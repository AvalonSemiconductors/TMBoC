magic
tech sky130B
magscale 1 2
timestamp 1682099404
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 397454 700884 397460 700936
rect 397512 700924 397518 700936
rect 446490 700924 446496 700936
rect 397512 700896 446496 700924
rect 397512 700884 397518 700896
rect 446490 700884 446496 700896
rect 446548 700884 446554 700936
rect 364978 700816 364984 700868
rect 365036 700856 365042 700868
rect 445018 700856 445024 700868
rect 365036 700828 445024 700856
rect 365036 700816 365042 700828
rect 445018 700816 445024 700828
rect 445076 700816 445082 700868
rect 283834 700748 283840 700800
rect 283892 700788 283898 700800
rect 446582 700788 446588 700800
rect 283892 700760 446588 700788
rect 283892 700748 283898 700760
rect 446582 700748 446588 700760
rect 446640 700748 446646 700800
rect 235166 700680 235172 700732
rect 235224 700720 235230 700732
rect 445110 700720 445116 700732
rect 235224 700692 445116 700720
rect 235224 700680 235230 700692
rect 445110 700680 445116 700692
rect 445168 700680 445174 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 416038 700652 416044 700664
rect 154172 700624 416044 700652
rect 154172 700612 154178 700624
rect 416038 700612 416044 700624
rect 416096 700612 416102 700664
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 450538 700584 450544 700596
rect 137888 700556 450544 700584
rect 137888 700544 137894 700556
rect 450538 700544 450544 700556
rect 450596 700544 450602 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 444282 700516 444288 700528
rect 105504 700488 444288 700516
rect 105504 700476 105510 700488
rect 444282 700476 444288 700488
rect 444340 700476 444346 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 444098 700448 444104 700460
rect 73028 700420 444104 700448
rect 73028 700408 73034 700420
rect 444098 700408 444104 700420
rect 444156 700408 444162 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 450630 700380 450636 700392
rect 40552 700352 450636 700380
rect 40552 700340 40558 700352
rect 450630 700340 450636 700352
rect 450688 700340 450694 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 418798 700312 418804 700324
rect 8168 700284 418804 700312
rect 8168 700272 8174 700284
rect 418798 700272 418804 700284
rect 418856 700272 418862 700324
rect 429838 700272 429844 700324
rect 429896 700312 429902 700324
rect 446398 700312 446404 700324
rect 429896 700284 446404 700312
rect 429896 700272 429902 700284
rect 446398 700272 446404 700284
rect 446456 700272 446462 700324
rect 447778 700272 447784 700324
rect 447836 700312 447842 700324
rect 478506 700312 478512 700324
rect 447836 700284 478512 700312
rect 447836 700272 447842 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 573358 696940 573364 696992
rect 573416 696980 573422 696992
rect 580166 696980 580172 696992
rect 573416 696952 580172 696980
rect 573416 696940 573422 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 218054 686536 218060 686588
rect 218112 686576 218118 686588
rect 445202 686576 445208 686588
rect 218112 686548 445208 686576
rect 218112 686536 218118 686548
rect 445202 686536 445208 686548
rect 445260 686536 445266 686588
rect 201494 686468 201500 686520
rect 201552 686508 201558 686520
rect 445294 686508 445300 686520
rect 201552 686480 445300 686508
rect 201552 686468 201558 686480
rect 445294 686468 445300 686480
rect 445352 686468 445358 686520
rect 347774 685176 347780 685228
rect 347832 685216 347838 685228
rect 446674 685216 446680 685228
rect 347832 685188 446680 685216
rect 347832 685176 347838 685188
rect 446674 685176 446680 685188
rect 446732 685176 446738 685228
rect 266354 685108 266360 685160
rect 266412 685148 266418 685160
rect 418982 685148 418988 685160
rect 266412 685120 418988 685148
rect 266412 685108 266418 685120
rect 418982 685108 418988 685120
rect 419040 685108 419046 685160
rect 19978 684768 19984 684820
rect 20036 684808 20042 684820
rect 418890 684808 418896 684820
rect 20036 684780 418896 684808
rect 20036 684768 20042 684780
rect 418890 684768 418896 684780
rect 418948 684768 418954 684820
rect 3602 684700 3608 684752
rect 3660 684740 3666 684752
rect 420178 684740 420184 684752
rect 3660 684712 420184 684740
rect 3660 684700 3666 684712
rect 420178 684700 420184 684712
rect 420236 684700 420242 684752
rect 3326 684632 3332 684684
rect 3384 684672 3390 684684
rect 420270 684672 420276 684684
rect 3384 684644 420276 684672
rect 3384 684632 3390 684644
rect 420270 684632 420276 684644
rect 420328 684632 420334 684684
rect 3142 684564 3148 684616
rect 3200 684604 3206 684616
rect 420362 684604 420368 684616
rect 3200 684576 420368 684604
rect 3200 684564 3206 684576
rect 420362 684564 420368 684576
rect 420420 684564 420426 684616
rect 3878 684496 3884 684548
rect 3936 684536 3942 684548
rect 445386 684536 445392 684548
rect 3936 684508 445392 684536
rect 3936 684496 3942 684508
rect 445386 684496 445392 684508
rect 445444 684496 445450 684548
rect 17954 683544 17960 683596
rect 18012 683584 18018 683596
rect 359458 683584 359464 683596
rect 18012 683556 359464 683584
rect 18012 683544 18018 683556
rect 359458 683544 359464 683556
rect 359516 683544 359522 683596
rect 21358 683476 21364 683528
rect 21416 683516 21422 683528
rect 420546 683516 420552 683528
rect 21416 683488 420552 683516
rect 21416 683476 21422 683488
rect 420546 683476 420552 683488
rect 420604 683476 420610 683528
rect 4062 683408 4068 683460
rect 4120 683448 4126 683460
rect 420638 683448 420644 683460
rect 4120 683420 420644 683448
rect 4120 683408 4126 683420
rect 420638 683408 420644 683420
rect 420696 683408 420702 683460
rect 3510 683340 3516 683392
rect 3568 683380 3574 683392
rect 420730 683380 420736 683392
rect 3568 683352 420736 683380
rect 3568 683340 3574 683352
rect 420730 683340 420736 683352
rect 420788 683340 420794 683392
rect 3694 683272 3700 683324
rect 3752 683312 3758 683324
rect 445478 683312 445484 683324
rect 3752 683284 445484 683312
rect 3752 683272 3758 683284
rect 445478 683272 445484 683284
rect 445536 683272 445542 683324
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 445570 683244 445576 683256
rect 3476 683216 445576 683244
rect 3476 683204 3482 683216
rect 445570 683204 445576 683216
rect 445628 683204 445634 683256
rect 3970 683136 3976 683188
rect 4028 683176 4034 683188
rect 446766 683176 446772 683188
rect 4028 683148 446772 683176
rect 4028 683136 4034 683148
rect 446766 683136 446772 683148
rect 446824 683136 446830 683188
rect 2958 682728 2964 682780
rect 3016 682768 3022 682780
rect 420086 682768 420092 682780
rect 3016 682740 420092 682768
rect 3016 682728 3022 682740
rect 420086 682728 420092 682740
rect 420144 682728 420150 682780
rect 2866 682660 2872 682712
rect 2924 682700 2930 682712
rect 450446 682700 450452 682712
rect 2924 682672 450452 682700
rect 2924 682660 2930 682672
rect 450446 682660 450452 682672
rect 450504 682660 450510 682712
rect 17862 680388 17868 680400
rect 16546 680360 17868 680388
rect 12894 680280 12900 680332
rect 12952 680320 12958 680332
rect 16546 680320 16574 680360
rect 17862 680348 17868 680360
rect 17920 680348 17926 680400
rect 12952 680292 16574 680320
rect 12952 680280 12958 680292
rect 361758 678988 361764 679040
rect 361816 679028 361822 679040
rect 364978 679028 364984 679040
rect 361816 679000 364984 679028
rect 361816 678988 361822 679000
rect 364978 678988 364984 679000
rect 365036 678988 365042 679040
rect 3510 678512 3516 678564
rect 3568 678512 3574 678564
rect 3602 678512 3608 678564
rect 3660 678552 3666 678564
rect 3660 678524 3924 678552
rect 3660 678512 3666 678524
rect 3528 678360 3556 678512
rect 3510 678308 3516 678360
rect 3568 678308 3574 678360
rect 3896 678224 3924 678524
rect 3878 678172 3884 678224
rect 3936 678172 3942 678224
rect 12894 676240 12900 676252
rect 11072 676212 12900 676240
rect 10410 676132 10416 676184
rect 10468 676172 10474 676184
rect 11072 676172 11100 676212
rect 12894 676200 12900 676212
rect 12952 676200 12958 676252
rect 10468 676144 11100 676172
rect 10468 676132 10474 676144
rect 569218 670692 569224 670744
rect 569276 670732 569282 670744
rect 580166 670732 580172 670744
rect 569276 670704 580172 670732
rect 569276 670692 569282 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 8018 667904 8024 667956
rect 8076 667944 8082 667956
rect 10410 667944 10416 667956
rect 8076 667916 10416 667944
rect 8076 667904 8082 667916
rect 10410 667904 10416 667916
rect 10468 667904 10474 667956
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 381538 667944 381544 667956
rect 361816 667916 381544 667944
rect 361816 667904 361822 667916
rect 381538 667904 381544 667916
rect 381596 667904 381602 667956
rect 4798 665184 4804 665236
rect 4856 665224 4862 665236
rect 8018 665224 8024 665236
rect 4856 665196 8024 665224
rect 4856 665184 4862 665196
rect 8018 665184 8024 665196
rect 8076 665184 8082 665236
rect 3142 658180 3148 658232
rect 3200 658220 3206 658232
rect 19978 658220 19984 658232
rect 3200 658192 19984 658220
rect 3200 658180 3206 658192
rect 19978 658180 19984 658192
rect 20036 658180 20042 658232
rect 361666 656140 361672 656192
rect 361724 656180 361730 656192
rect 406378 656180 406384 656192
rect 361724 656152 406384 656180
rect 361724 656140 361730 656152
rect 406378 656140 406384 656152
rect 406436 656140 406442 656192
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 378778 645912 378784 645924
rect 361816 645884 378784 645912
rect 361816 645872 361822 645884
rect 378778 645872 378784 645884
rect 378836 645872 378842 645924
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 407758 634828 407764 634840
rect 361632 634800 407764 634828
rect 361632 634788 361638 634800
rect 407758 634788 407764 634800
rect 407816 634788 407822 634840
rect 3694 631320 3700 631372
rect 3752 631360 3758 631372
rect 20898 631360 20904 631372
rect 3752 631332 20904 631360
rect 3752 631320 3758 631332
rect 20898 631320 20904 631332
rect 20956 631320 20962 631372
rect 576118 630640 576124 630692
rect 576176 630680 576182 630692
rect 579982 630680 579988 630692
rect 576176 630652 579988 630680
rect 576176 630640 576182 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 376018 623812 376024 623824
rect 361632 623784 376024 623812
rect 361632 623772 361638 623784
rect 376018 623772 376024 623784
rect 376076 623772 376082 623824
rect 361574 612756 361580 612808
rect 361632 612796 361638 612808
rect 410518 612796 410524 612808
rect 361632 612768 410524 612796
rect 361632 612756 361638 612768
rect 410518 612756 410524 612768
rect 410576 612756 410582 612808
rect 359458 601672 359464 601724
rect 359516 601712 359522 601724
rect 359516 601684 360240 601712
rect 359516 601672 359522 601684
rect 360212 601644 360240 601684
rect 361758 601672 361764 601724
rect 361816 601712 361822 601724
rect 374730 601712 374736 601724
rect 361816 601684 374736 601712
rect 361816 601672 361822 601684
rect 374730 601672 374736 601684
rect 374788 601672 374794 601724
rect 366358 601644 366364 601656
rect 360212 601616 366364 601644
rect 366358 601604 366364 601616
rect 366416 601604 366422 601656
rect 457530 600584 457536 600636
rect 457588 600624 457594 600636
rect 461578 600624 461584 600636
rect 457588 600596 461584 600624
rect 457588 600584 457594 600596
rect 461578 600584 461584 600596
rect 461636 600584 461642 600636
rect 457346 599972 457352 600024
rect 457404 600012 457410 600024
rect 462958 600012 462964 600024
rect 457404 599984 462964 600012
rect 457404 599972 457410 599984
rect 462958 599972 462964 599984
rect 463016 599972 463022 600024
rect 460198 599768 460204 599820
rect 460256 599808 460262 599820
rect 463694 599808 463700 599820
rect 460256 599780 463700 599808
rect 460256 599768 460262 599780
rect 463694 599768 463700 599780
rect 463752 599768 463758 599820
rect 458818 599632 458824 599684
rect 458876 599672 458882 599684
rect 466454 599672 466460 599684
rect 458876 599644 466460 599672
rect 458876 599632 458882 599644
rect 466454 599632 466460 599644
rect 466512 599632 466518 599684
rect 457898 599564 457904 599616
rect 457956 599604 457962 599616
rect 469858 599604 469864 599616
rect 457956 599576 469864 599604
rect 457956 599564 457962 599576
rect 469858 599564 469864 599576
rect 469916 599564 469922 599616
rect 459922 598340 459928 598392
rect 459980 598380 459986 598392
rect 463786 598380 463792 598392
rect 459980 598352 463792 598380
rect 459980 598340 459986 598352
rect 463786 598340 463792 598352
rect 463844 598340 463850 598392
rect 457714 598272 457720 598324
rect 457772 598312 457778 598324
rect 464338 598312 464344 598324
rect 457772 598284 464344 598312
rect 457772 598272 457778 598284
rect 464338 598272 464344 598284
rect 464396 598272 464402 598324
rect 488626 598272 488632 598324
rect 488684 598312 488690 598324
rect 494238 598312 494244 598324
rect 488684 598284 494244 598312
rect 488684 598272 488690 598284
rect 494238 598272 494244 598284
rect 494296 598272 494302 598324
rect 457622 598204 457628 598256
rect 457680 598244 457686 598256
rect 468478 598244 468484 598256
rect 457680 598216 468484 598244
rect 457680 598204 457686 598216
rect 468478 598204 468484 598216
rect 468536 598204 468542 598256
rect 482278 598204 482284 598256
rect 482336 598244 482342 598256
rect 494054 598244 494060 598256
rect 482336 598216 494060 598244
rect 482336 598204 482342 598216
rect 494054 598204 494060 598216
rect 494112 598204 494118 598256
rect 493318 597864 493324 597916
rect 493376 597904 493382 597916
rect 494974 597904 494980 597916
rect 493376 597876 494980 597904
rect 493376 597864 493382 597876
rect 494974 597864 494980 597876
rect 495032 597864 495038 597916
rect 458726 596912 458732 596964
rect 458784 596952 458790 596964
rect 465074 596952 465080 596964
rect 458784 596924 465080 596952
rect 458784 596912 458790 596924
rect 465074 596912 465080 596924
rect 465132 596912 465138 596964
rect 459830 596844 459836 596896
rect 459888 596884 459894 596896
rect 466546 596884 466552 596896
rect 459888 596856 466552 596884
rect 459888 596844 459894 596856
rect 466546 596844 466552 596856
rect 466604 596844 466610 596896
rect 459738 596776 459744 596828
rect 459796 596816 459802 596828
rect 470870 596816 470876 596828
rect 459796 596788 470876 596816
rect 459796 596776 459802 596788
rect 470870 596776 470876 596788
rect 470928 596776 470934 596828
rect 457438 596164 457444 596216
rect 457496 596204 457502 596216
rect 461670 596204 461676 596216
rect 457496 596176 461676 596204
rect 457496 596164 457502 596176
rect 461670 596164 461676 596176
rect 461728 596164 461734 596216
rect 361758 590656 361764 590708
rect 361816 590696 361822 590708
rect 371878 590696 371884 590708
rect 361816 590668 371884 590696
rect 361816 590656 361822 590668
rect 371878 590656 371884 590668
rect 371936 590656 371942 590708
rect 571978 590656 571984 590708
rect 572036 590696 572042 590708
rect 579614 590696 579620 590708
rect 572036 590668 579620 590696
rect 572036 590656 572042 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 366358 590588 366364 590640
rect 366416 590628 366422 590640
rect 367554 590628 367560 590640
rect 366416 590600 367560 590628
rect 366416 590588 366422 590600
rect 367554 590588 367560 590600
rect 367612 590588 367618 590640
rect 367554 586508 367560 586560
rect 367612 586548 367618 586560
rect 367612 586520 369900 586548
rect 367612 586508 367618 586520
rect 369872 586480 369900 586520
rect 372522 586480 372528 586492
rect 369872 586452 372528 586480
rect 372522 586440 372528 586452
rect 372580 586440 372586 586492
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 370498 579680 370504 579692
rect 361816 579652 370504 579680
rect 361816 579640 361822 579652
rect 370498 579640 370504 579652
rect 370556 579640 370562 579692
rect 372614 577396 372620 577448
rect 372672 577436 372678 577448
rect 374822 577436 374828 577448
rect 372672 577408 374828 577436
rect 372672 577396 372678 577408
rect 374822 577396 374828 577408
rect 374880 577396 374886 577448
rect 511258 576852 511264 576904
rect 511316 576892 511322 576904
rect 579614 576892 579620 576904
rect 511316 576864 579620 576892
rect 511316 576852 511322 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 374822 571956 374828 572008
rect 374880 571996 374886 572008
rect 376202 571996 376208 572008
rect 374880 571968 376208 571996
rect 374880 571956 374886 571968
rect 376202 571956 376208 571968
rect 376260 571956 376266 572008
rect 361758 568556 361764 568608
rect 361816 568596 361822 568608
rect 367738 568596 367744 568608
rect 361816 568568 367744 568596
rect 361816 568556 361822 568568
rect 367738 568556 367744 568568
rect 367796 568556 367802 568608
rect 376202 568488 376208 568540
rect 376260 568528 376266 568540
rect 377398 568528 377404 568540
rect 376260 568500 377404 568528
rect 376260 568488 376266 568500
rect 377398 568488 377404 568500
rect 377456 568488 377462 568540
rect 377398 564068 377404 564120
rect 377456 564108 377462 564120
rect 380342 564108 380348 564120
rect 377456 564080 380348 564108
rect 377456 564068 377462 564080
rect 380342 564068 380348 564080
rect 380400 564068 380406 564120
rect 380342 559172 380348 559224
rect 380400 559212 380406 559224
rect 384942 559212 384948 559224
rect 380400 559184 384948 559212
rect 380400 559172 380406 559184
rect 384942 559172 384948 559184
rect 385000 559172 385006 559224
rect 361574 557744 361580 557796
rect 361632 557784 361638 557796
rect 363598 557784 363604 557796
rect 361632 557756 363604 557784
rect 361632 557744 361638 557756
rect 363598 557744 363604 557756
rect 363656 557744 363662 557796
rect 385034 551964 385040 552016
rect 385092 552004 385098 552016
rect 387058 552004 387064 552016
rect 385092 551976 387064 552004
rect 385092 551964 385098 551976
rect 387058 551964 387064 551976
rect 387116 551964 387122 552016
rect 361574 546592 361580 546644
rect 361632 546632 361638 546644
rect 363690 546632 363696 546644
rect 361632 546604 363696 546632
rect 361632 546592 361638 546604
rect 363690 546592 363696 546604
rect 363748 546592 363754 546644
rect 457806 542988 457812 543040
rect 457864 543028 457870 543040
rect 468570 543028 468576 543040
rect 457864 543000 468576 543028
rect 457864 542988 457870 543000
rect 468570 542988 468576 543000
rect 468628 542988 468634 543040
rect 459554 541628 459560 541680
rect 459612 541668 459618 541680
rect 470686 541668 470692 541680
rect 459612 541640 470692 541668
rect 459612 541628 459618 541640
rect 470686 541628 470692 541640
rect 470744 541628 470750 541680
rect 387058 540880 387064 540932
rect 387116 540920 387122 540932
rect 388438 540920 388444 540932
rect 387116 540892 388444 540920
rect 387116 540880 387122 540892
rect 388438 540880 388444 540892
rect 388496 540880 388502 540932
rect 519538 536800 519544 536852
rect 519596 536840 519602 536852
rect 580166 536840 580172 536852
rect 519596 536812 580172 536840
rect 519596 536800 519602 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 361574 535712 361580 535764
rect 361632 535752 361638 535764
rect 363782 535752 363788 535764
rect 361632 535724 363788 535752
rect 361632 535712 361638 535724
rect 363782 535712 363788 535724
rect 363840 535712 363846 535764
rect 448054 526396 448060 526448
rect 448112 526436 448118 526448
rect 500954 526436 500960 526448
rect 448112 526408 500960 526436
rect 448112 526396 448118 526408
rect 500954 526396 500960 526408
rect 501012 526396 501018 526448
rect 457254 525036 457260 525088
rect 457312 525076 457318 525088
rect 465166 525076 465172 525088
rect 457312 525048 465172 525076
rect 457312 525036 457318 525048
rect 465166 525036 465172 525048
rect 465224 525036 465230 525088
rect 361758 524424 361764 524476
rect 361816 524464 361822 524476
rect 411898 524464 411904 524476
rect 361816 524436 411904 524464
rect 361816 524424 361822 524436
rect 411898 524424 411904 524436
rect 411956 524424 411962 524476
rect 511350 524424 511356 524476
rect 511408 524464 511414 524476
rect 580166 524464 580172 524476
rect 511408 524436 580172 524464
rect 511408 524424 511414 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 448422 523676 448428 523728
rect 448480 523716 448486 523728
rect 506474 523716 506480 523728
rect 448480 523688 506480 523716
rect 448480 523676 448486 523688
rect 506474 523676 506480 523688
rect 506532 523676 506538 523728
rect 448330 522248 448336 522300
rect 448388 522288 448394 522300
rect 493318 522288 493324 522300
rect 448388 522260 493324 522288
rect 448388 522248 448394 522260
rect 493318 522248 493324 522260
rect 493376 522248 493382 522300
rect 474734 521636 474740 521688
rect 474792 521676 474798 521688
rect 475194 521676 475200 521688
rect 474792 521648 475200 521676
rect 474792 521636 474798 521648
rect 475194 521636 475200 521648
rect 475252 521676 475258 521688
rect 494330 521676 494336 521688
rect 475252 521648 494336 521676
rect 475252 521636 475258 521648
rect 494330 521636 494336 521648
rect 494388 521636 494394 521688
rect 458082 520956 458088 521008
rect 458140 520996 458146 521008
rect 465718 520996 465724 521008
rect 458140 520968 465724 520996
rect 458140 520956 458146 520968
rect 465718 520956 465724 520968
rect 465776 520956 465782 521008
rect 449710 520888 449716 520940
rect 449768 520928 449774 520940
rect 475194 520928 475200 520940
rect 449768 520900 475200 520928
rect 449768 520888 449774 520900
rect 475194 520888 475200 520900
rect 475252 520888 475258 520940
rect 482646 520888 482652 520940
rect 482704 520928 482710 520940
rect 520274 520928 520280 520940
rect 482704 520900 520280 520928
rect 482704 520888 482710 520900
rect 520274 520888 520280 520900
rect 520332 520888 520338 520940
rect 461762 520412 461768 520464
rect 461820 520452 461826 520464
rect 488626 520452 488632 520464
rect 461820 520424 488632 520452
rect 461820 520412 461826 520424
rect 488626 520412 488632 520424
rect 488684 520412 488690 520464
rect 467834 520344 467840 520396
rect 467892 520384 467898 520396
rect 469122 520384 469128 520396
rect 467892 520356 469128 520384
rect 467892 520344 467898 520356
rect 469122 520344 469128 520356
rect 469180 520384 469186 520396
rect 494238 520384 494244 520396
rect 469180 520356 494244 520384
rect 469180 520344 469186 520356
rect 494238 520344 494244 520356
rect 494296 520344 494302 520396
rect 477402 520276 477408 520328
rect 477460 520316 477466 520328
rect 482646 520316 482652 520328
rect 477460 520288 482652 520316
rect 477460 520276 477466 520288
rect 482646 520276 482652 520288
rect 482704 520276 482710 520328
rect 457990 519596 457996 519648
rect 458048 519636 458054 519648
rect 468754 519636 468760 519648
rect 458048 519608 468760 519636
rect 458048 519596 458054 519608
rect 468754 519596 468760 519608
rect 468812 519596 468818 519648
rect 447962 519528 447968 519580
rect 448020 519568 448026 519580
rect 467834 519568 467840 519580
rect 448020 519540 467840 519568
rect 448020 519528 448026 519540
rect 467834 519528 467840 519540
rect 467892 519528 467898 519580
rect 449802 518168 449808 518220
rect 449860 518208 449866 518220
rect 462406 518208 462412 518220
rect 449860 518180 462412 518208
rect 449860 518168 449866 518180
rect 462406 518168 462412 518180
rect 462464 518168 462470 518220
rect 388438 517488 388444 517540
rect 388496 517528 388502 517540
rect 389450 517528 389456 517540
rect 388496 517500 389456 517528
rect 388496 517488 388502 517500
rect 389450 517488 389456 517500
rect 389508 517488 389514 517540
rect 459646 517488 459652 517540
rect 459704 517528 459710 517540
rect 462498 517528 462504 517540
rect 459704 517500 462504 517528
rect 459704 517488 459710 517500
rect 462498 517488 462504 517500
rect 462556 517488 462562 517540
rect 491846 516168 491852 516180
rect 448440 516140 491852 516168
rect 448440 516112 448468 516140
rect 491846 516128 491852 516140
rect 491904 516128 491910 516180
rect 448422 516060 448428 516112
rect 448480 516060 448486 516112
rect 494054 515380 494060 515432
rect 494112 515420 494118 515432
rect 538214 515420 538220 515432
rect 494112 515392 538220 515420
rect 494112 515380 494118 515392
rect 538214 515380 538220 515392
rect 538272 515380 538278 515432
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 414658 513380 414664 513392
rect 361816 513352 414664 513380
rect 361816 513340 361822 513352
rect 414658 513340 414664 513352
rect 414716 513340 414722 513392
rect 494054 512592 494060 512644
rect 494112 512632 494118 512644
rect 494422 512632 494428 512644
rect 494112 512604 494428 512632
rect 494112 512592 494118 512604
rect 494422 512592 494428 512604
rect 494480 512632 494486 512644
rect 535454 512632 535460 512644
rect 494480 512604 535460 512632
rect 494480 512592 494486 512604
rect 535454 512592 535460 512604
rect 535512 512592 535518 512644
rect 389450 511980 389456 512032
rect 389508 512020 389514 512032
rect 389508 511992 390876 512020
rect 389508 511980 389514 511992
rect 390848 511952 390876 511992
rect 393222 511952 393228 511964
rect 390848 511924 393228 511952
rect 393222 511912 393228 511924
rect 393280 511912 393286 511964
rect 567838 510620 567844 510672
rect 567896 510660 567902 510672
rect 580166 510660 580172 510672
rect 567896 510632 580172 510660
rect 567896 510620 567902 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 494330 508512 494336 508564
rect 494388 508552 494394 508564
rect 532694 508552 532700 508564
rect 494388 508524 532700 508552
rect 494388 508512 494394 508524
rect 532694 508512 532700 508524
rect 532752 508512 532758 508564
rect 393314 506744 393320 506796
rect 393372 506784 393378 506796
rect 396718 506784 396724 506796
rect 393372 506756 396724 506784
rect 393372 506744 393378 506756
rect 396718 506744 396724 506756
rect 396776 506744 396782 506796
rect 495066 505724 495072 505776
rect 495124 505764 495130 505776
rect 529934 505764 529940 505776
rect 495124 505736 529940 505764
rect 495124 505724 495130 505736
rect 529934 505724 529940 505736
rect 529992 505724 529998 505776
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 416130 502364 416136 502376
rect 361816 502336 416136 502364
rect 361816 502324 361822 502336
rect 416130 502324 416136 502336
rect 416188 502324 416194 502376
rect 448514 500216 448520 500268
rect 448572 500256 448578 500268
rect 545114 500256 545120 500268
rect 448572 500228 545120 500256
rect 448572 500216 448578 500228
rect 545114 500216 545120 500228
rect 545172 500216 545178 500268
rect 448514 498788 448520 498840
rect 448572 498828 448578 498840
rect 542446 498828 542452 498840
rect 448572 498800 542452 498828
rect 448572 498788 448578 498800
rect 542446 498788 542452 498800
rect 542504 498788 542510 498840
rect 453298 497428 453304 497480
rect 453356 497468 453362 497480
rect 480254 497468 480260 497480
rect 453356 497440 480260 497468
rect 453356 497428 453362 497440
rect 480254 497428 480260 497440
rect 480312 497428 480318 497480
rect 454034 497020 454040 497072
rect 454092 497060 454098 497072
rect 459554 497060 459560 497072
rect 454092 497032 459560 497060
rect 454092 497020 454098 497032
rect 459554 497020 459560 497032
rect 459612 497020 459618 497072
rect 454126 496952 454132 497004
rect 454184 496992 454190 497004
rect 458082 496992 458088 497004
rect 454184 496964 458088 496992
rect 454184 496952 454190 496964
rect 458082 496952 458088 496964
rect 458140 496952 458146 497004
rect 452838 496884 452844 496936
rect 452896 496924 452902 496936
rect 455138 496924 455144 496936
rect 452896 496896 455144 496924
rect 452896 496884 452902 496896
rect 455138 496884 455144 496896
rect 455196 496884 455202 496936
rect 455414 496884 455420 496936
rect 455472 496924 455478 496936
rect 461026 496924 461032 496936
rect 455472 496896 461032 496924
rect 455472 496884 455478 496896
rect 461026 496884 461032 496896
rect 461084 496884 461090 496936
rect 451366 496816 451372 496868
rect 451424 496856 451430 496868
rect 453666 496856 453672 496868
rect 451424 496828 453672 496856
rect 451424 496816 451430 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 454678 496816 454684 496868
rect 454736 496856 454742 496868
rect 456610 496856 456616 496868
rect 454736 496828 456616 496856
rect 454736 496816 454742 496828
rect 456610 496816 456616 496828
rect 456668 496816 456674 496868
rect 448422 496068 448428 496120
rect 448480 496108 448486 496120
rect 547874 496108 547880 496120
rect 448480 496080 547880 496108
rect 448480 496068 448486 496080
rect 547874 496068 547880 496080
rect 547932 496068 547938 496120
rect 449986 494708 449992 494760
rect 450044 494748 450050 494760
rect 450722 494748 450728 494760
rect 450044 494720 450728 494748
rect 450044 494708 450050 494720
rect 450722 494708 450728 494720
rect 450780 494708 450786 494760
rect 361758 491308 361764 491360
rect 361816 491348 361822 491360
rect 417418 491348 417424 491360
rect 361816 491320 417424 491348
rect 361816 491308 361822 491320
rect 417418 491308 417424 491320
rect 417476 491308 417482 491360
rect 518158 484372 518164 484424
rect 518216 484412 518222 484424
rect 580166 484412 580172 484424
rect 518216 484384 580172 484412
rect 518216 484372 518222 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 419074 480264 419080 480276
rect 361816 480236 419080 480264
rect 361816 480224 361822 480236
rect 419074 480224 419080 480236
rect 419132 480224 419138 480276
rect 396718 476076 396724 476128
rect 396776 476116 396782 476128
rect 396776 476088 397500 476116
rect 396776 476076 396782 476088
rect 397472 476048 397500 476088
rect 400858 476048 400864 476060
rect 397472 476020 400864 476048
rect 400858 476008 400864 476020
rect 400916 476008 400922 476060
rect 516778 470568 516784 470620
rect 516836 470608 516842 470620
rect 579614 470608 579620 470620
rect 516836 470580 579620 470608
rect 516836 470568 516842 470580
rect 579614 470568 579620 470580
rect 579672 470568 579678 470620
rect 400858 468188 400864 468240
rect 400916 468228 400922 468240
rect 401962 468228 401968 468240
rect 400916 468200 401968 468228
rect 400916 468188 400922 468200
rect 401962 468188 401968 468200
rect 402020 468188 402026 468240
rect 401962 464992 401968 465044
rect 402020 465032 402026 465044
rect 403618 465032 403624 465044
rect 402020 465004 403624 465032
rect 402020 464992 402026 465004
rect 403618 464992 403624 465004
rect 403676 464992 403682 465044
rect 515398 464380 515404 464432
rect 515456 464420 515462 464432
rect 542354 464420 542360 464432
rect 515456 464392 542360 464420
rect 515456 464380 515462 464392
rect 542354 464380 542360 464392
rect 542412 464380 542418 464432
rect 449802 464312 449808 464364
rect 449860 464352 449866 464364
rect 525794 464352 525800 464364
rect 449860 464324 525800 464352
rect 449860 464312 449866 464324
rect 525794 464312 525800 464324
rect 525852 464312 525858 464364
rect 488258 462952 488264 463004
rect 488316 462992 488322 463004
rect 494054 462992 494060 463004
rect 488316 462964 494060 462992
rect 488316 462952 488322 462964
rect 494054 462952 494060 462964
rect 494112 462992 494118 463004
rect 527634 462992 527640 463004
rect 494112 462964 527640 462992
rect 494112 462952 494118 462964
rect 527634 462952 527640 462964
rect 527692 462952 527698 463004
rect 436094 462408 436100 462460
rect 436152 462448 436158 462460
rect 554130 462448 554136 462460
rect 436152 462420 554136 462448
rect 436152 462408 436158 462420
rect 554130 462408 554136 462420
rect 554188 462408 554194 462460
rect 431954 462340 431960 462392
rect 432012 462380 432018 462392
rect 551186 462380 551192 462392
rect 432012 462352 551192 462380
rect 432012 462340 432018 462352
rect 551186 462340 551192 462352
rect 551244 462340 551250 462392
rect 477402 461592 477408 461644
rect 477460 461632 477466 461644
rect 521746 461632 521752 461644
rect 477460 461604 521752 461632
rect 477460 461592 477466 461604
rect 521746 461592 521752 461604
rect 521804 461592 521810 461644
rect 476022 461456 476028 461508
rect 476080 461496 476086 461508
rect 477402 461496 477408 461508
rect 476080 461468 477408 461496
rect 476080 461456 476086 461468
rect 477402 461456 477408 461468
rect 477460 461456 477466 461508
rect 449894 460912 449900 460964
rect 449952 460952 449958 460964
rect 524414 460952 524420 460964
rect 449952 460924 524420 460952
rect 449952 460912 449958 460924
rect 524414 460912 524420 460924
rect 524472 460912 524478 460964
rect 449710 460164 449716 460216
rect 449768 460204 449774 460216
rect 485774 460204 485780 460216
rect 449768 460176 485780 460204
rect 449768 460164 449774 460176
rect 485774 460164 485780 460176
rect 485832 460164 485838 460216
rect 449618 458804 449624 458856
rect 449676 458844 449682 458856
rect 488534 458844 488540 458856
rect 449676 458816 488540 458844
rect 449676 458804 449682 458816
rect 488534 458804 488540 458816
rect 488592 458804 488598 458856
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 383010 458232 383016 458244
rect 361816 458204 383016 458232
rect 361816 458192 361822 458204
rect 383010 458192 383016 458204
rect 383068 458192 383074 458244
rect 449434 457444 449440 457496
rect 449492 457484 449498 457496
rect 487154 457484 487160 457496
rect 449492 457456 487160 457484
rect 449492 457444 449498 457456
rect 487154 457444 487160 457456
rect 487212 457444 487218 457496
rect 403618 456764 403624 456816
rect 403676 456804 403682 456816
rect 403676 456776 405780 456804
rect 403676 456764 403682 456776
rect 405752 456736 405780 456776
rect 408402 456736 408408 456748
rect 405752 456708 408408 456736
rect 408402 456696 408408 456708
rect 408460 456696 408466 456748
rect 473722 456492 473728 456544
rect 473780 456532 473786 456544
rect 476022 456532 476028 456544
rect 473780 456504 476028 456532
rect 473780 456492 473786 456504
rect 476022 456492 476028 456504
rect 476080 456492 476086 456544
rect 451918 455472 451924 455524
rect 451976 455512 451982 455524
rect 480990 455512 480996 455524
rect 451976 455484 480996 455512
rect 451976 455472 451982 455484
rect 480990 455472 480996 455484
rect 481048 455472 481054 455524
rect 423582 455404 423588 455456
rect 423640 455444 423646 455456
rect 473722 455444 473728 455456
rect 423640 455416 473728 455444
rect 423640 455404 423646 455416
rect 473722 455404 473728 455416
rect 473780 455404 473786 455456
rect 449526 454724 449532 454776
rect 449584 454764 449590 454776
rect 481634 454764 481640 454776
rect 449584 454736 481640 454764
rect 449584 454724 449590 454736
rect 481634 454724 481640 454736
rect 481692 454724 481698 454776
rect 449342 454656 449348 454708
rect 449400 454696 449406 454708
rect 484394 454696 484400 454708
rect 449400 454668 484400 454696
rect 449400 454656 449406 454668
rect 484394 454656 484400 454668
rect 484452 454656 484458 454708
rect 408494 452548 408500 452600
rect 408552 452588 408558 452600
rect 410334 452588 410340 452600
rect 408552 452560 410340 452588
rect 408552 452548 408558 452560
rect 410334 452548 410340 452560
rect 410392 452548 410398 452600
rect 422478 447516 422484 447568
rect 422536 447556 422542 447568
rect 423582 447556 423588 447568
rect 422536 447528 423588 447556
rect 422536 447516 422542 447528
rect 423582 447516 423588 447528
rect 423640 447516 423646 447568
rect 427446 447176 427452 447228
rect 427504 447216 427510 447228
rect 446858 447216 446864 447228
rect 427504 447188 446864 447216
rect 427504 447176 427510 447188
rect 446858 447176 446864 447188
rect 446916 447176 446922 447228
rect 423582 447108 423588 447160
rect 423640 447148 423646 447160
rect 443362 447148 443368 447160
rect 423640 447120 443368 447148
rect 423640 447108 423646 447120
rect 443362 447108 443368 447120
rect 443420 447108 443426 447160
rect 410334 447040 410340 447092
rect 410392 447080 410398 447092
rect 413278 447080 413284 447092
rect 410392 447052 413284 447080
rect 410392 447040 410398 447052
rect 413278 447040 413284 447052
rect 413336 447040 413342 447092
rect 436094 445680 436100 445732
rect 436152 445720 436158 445732
rect 437382 445720 437388 445732
rect 436152 445692 437388 445720
rect 436152 445680 436158 445692
rect 437382 445680 437388 445692
rect 437440 445680 437446 445732
rect 432690 444524 432696 444576
rect 432748 444564 432754 444576
rect 445754 444564 445760 444576
rect 432748 444536 445760 444564
rect 432748 444524 432754 444536
rect 445754 444524 445760 444536
rect 445812 444524 445818 444576
rect 437290 444456 437296 444508
rect 437348 444496 437354 444508
rect 445846 444496 445852 444508
rect 437348 444468 445852 444496
rect 437348 444456 437354 444468
rect 445846 444456 445852 444468
rect 445904 444456 445910 444508
rect 442626 444388 442632 444440
rect 442684 444428 442690 444440
rect 445938 444428 445944 444440
rect 442684 444400 445944 444428
rect 442684 444388 442690 444400
rect 445938 444388 445944 444400
rect 445996 444388 446002 444440
rect 443362 444320 443368 444372
rect 443420 444360 443426 444372
rect 447870 444360 447876 444372
rect 443420 444332 447876 444360
rect 443420 444320 443426 444332
rect 447870 444320 447876 444332
rect 447928 444320 447934 444372
rect 413278 438268 413284 438320
rect 413336 438308 413342 438320
rect 414750 438308 414756 438320
rect 413336 438280 414756 438308
rect 413336 438268 413342 438280
rect 414750 438268 414756 438280
rect 414808 438268 414814 438320
rect 361758 436092 361764 436144
rect 361816 436132 361822 436144
rect 419166 436132 419172 436144
rect 361816 436104 419172 436132
rect 361816 436092 361822 436104
rect 419166 436092 419172 436104
rect 419224 436092 419230 436144
rect 574738 430584 574744 430636
rect 574796 430624 574802 430636
rect 579614 430624 579620 430636
rect 574796 430596 579620 430624
rect 574796 430584 574802 430596
rect 579614 430584 579620 430596
rect 579672 430584 579678 430636
rect 456886 429972 456892 430024
rect 456944 430012 456950 430024
rect 474274 430012 474280 430024
rect 456944 429984 474280 430012
rect 456944 429972 456950 429984
rect 474274 429972 474280 429984
rect 474332 429972 474338 430024
rect 458174 429904 458180 429956
rect 458232 429944 458238 429956
rect 476942 429944 476948 429956
rect 458232 429916 476948 429944
rect 458232 429904 458238 429916
rect 476942 429904 476948 429916
rect 477000 429904 477006 429956
rect 458358 429836 458364 429888
rect 458416 429876 458422 429888
rect 479334 429876 479340 429888
rect 458416 429848 479340 429876
rect 458416 429836 458422 429848
rect 479334 429836 479340 429848
rect 479392 429836 479398 429888
rect 479518 429836 479524 429888
rect 479576 429876 479582 429888
rect 484946 429876 484952 429888
rect 479576 429848 484952 429876
rect 479576 429836 479582 429848
rect 484946 429836 484952 429848
rect 485004 429836 485010 429888
rect 486418 429156 486424 429208
rect 486476 429196 486482 429208
rect 487614 429196 487620 429208
rect 486476 429168 487620 429196
rect 486476 429156 486482 429168
rect 487614 429156 487620 429168
rect 487672 429156 487678 429208
rect 457438 428408 457444 428460
rect 457496 428448 457502 428460
rect 471606 428448 471612 428460
rect 457496 428420 471612 428448
rect 457496 428408 457502 428420
rect 471606 428408 471612 428420
rect 471664 428408 471670 428460
rect 414750 426368 414756 426420
rect 414808 426408 414814 426420
rect 417510 426408 417516 426420
rect 414808 426380 417516 426408
rect 414808 426368 414814 426380
rect 417510 426368 417516 426380
rect 417568 426368 417574 426420
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 502978 423512 502984 423564
rect 503036 423552 503042 423564
rect 523770 423552 523776 423564
rect 503036 423524 523776 423552
rect 503036 423512 503042 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 444190 423376 444196 423428
rect 444248 423416 444254 423428
rect 447778 423416 447784 423428
rect 444248 423388 447784 423416
rect 444248 423376 444254 423388
rect 447778 423376 447784 423388
rect 447836 423376 447842 423428
rect 483014 423376 483020 423428
rect 483072 423416 483078 423428
rect 522482 423416 522488 423428
rect 483072 423388 522488 423416
rect 483072 423376 483078 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 485774 423308 485780 423360
rect 485832 423348 485838 423360
rect 526346 423348 526352 423360
rect 485832 423320 526352 423348
rect 485832 423308 485838 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 487154 423240 487160 423292
rect 487212 423280 487218 423292
rect 528922 423280 528928 423292
rect 487212 423252 528928 423280
rect 487212 423240 487218 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 488534 423172 488540 423224
rect 488592 423212 488598 423224
rect 531498 423212 531504 423224
rect 488592 423184 531504 423212
rect 488592 423172 488598 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 496814 423104 496820 423156
rect 496872 423144 496878 423156
rect 545666 423144 545672 423156
rect 496872 423116 545672 423144
rect 496872 423104 496878 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 498194 423036 498200 423088
rect 498252 423076 498258 423088
rect 548242 423076 548248 423088
rect 498252 423048 548248 423076
rect 498252 423036 498258 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 499574 422968 499580 423020
rect 499632 423008 499638 423020
rect 550818 423008 550824 423020
rect 499632 422980 550824 423008
rect 499632 422968 499638 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 501046 422900 501052 422952
rect 501104 422940 501110 422952
rect 553394 422940 553400 422952
rect 501104 422912 553400 422940
rect 501104 422900 501110 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 483106 421540 483112 421592
rect 483164 421580 483170 421592
rect 521194 421580 521200 421592
rect 483164 421552 521200 421580
rect 483164 421540 483170 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 417510 420452 417516 420504
rect 417568 420492 417574 420504
rect 424318 420492 424324 420504
rect 417568 420464 424324 420492
rect 417568 420452 417574 420464
rect 424318 420452 424324 420464
rect 424376 420452 424382 420504
rect 494054 420180 494060 420232
rect 494112 420220 494118 420232
rect 541802 420220 541808 420232
rect 494112 420192 541808 420220
rect 494112 420180 494118 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 362402 418752 362408 418804
rect 362460 418792 362466 418804
rect 443638 418792 443644 418804
rect 362460 418764 443644 418792
rect 362460 418752 362466 418764
rect 443638 418752 443644 418764
rect 443696 418752 443702 418804
rect 509878 418140 509884 418192
rect 509936 418180 509942 418192
rect 579706 418180 579712 418192
rect 509936 418152 579712 418180
rect 509936 418140 509942 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 421466 417732 421472 417784
rect 421524 417772 421530 417784
rect 503714 417772 503720 417784
rect 421524 417744 503720 417772
rect 421524 417732 421530 417744
rect 503714 417732 503720 417744
rect 503772 417732 503778 417784
rect 425974 417664 425980 417716
rect 426032 417704 426038 417716
rect 507854 417704 507860 417716
rect 426032 417676 507860 417704
rect 426032 417664 426038 417676
rect 507854 417664 507860 417676
rect 507912 417664 507918 417716
rect 425330 417596 425336 417648
rect 425388 417636 425394 417648
rect 507946 417636 507952 417648
rect 425388 417608 507952 417636
rect 425388 417596 425394 417608
rect 507946 417596 507952 417608
rect 508004 417596 508010 417648
rect 424042 417528 424048 417580
rect 424100 417568 424106 417580
rect 506474 417568 506480 417580
rect 424100 417540 506480 417568
rect 424100 417528 424106 417540
rect 506474 417528 506480 417540
rect 506532 417528 506538 417580
rect 424686 417460 424692 417512
rect 424744 417500 424750 417512
rect 506566 417500 506572 417512
rect 424744 417472 506572 417500
rect 424744 417460 424750 417472
rect 506566 417460 506572 417472
rect 506624 417460 506630 417512
rect 422110 417392 422116 417444
rect 422168 417432 422174 417444
rect 503990 417432 503996 417444
rect 422168 417404 503996 417432
rect 422168 417392 422174 417404
rect 503990 417392 503996 417404
rect 504048 417392 504054 417444
rect 362310 416032 362316 416084
rect 362368 416072 362374 416084
rect 440878 416072 440884 416084
rect 362368 416044 440884 416072
rect 362368 416032 362374 416044
rect 440878 416032 440884 416044
rect 440936 416032 440942 416084
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 442258 414032 442264 414044
rect 361632 414004 442264 414032
rect 361632 413992 361638 414004
rect 442258 413992 442264 414004
rect 442316 413992 442322 414044
rect 362218 413244 362224 413296
rect 362276 413284 362282 413296
rect 436738 413284 436744 413296
rect 362276 413256 436744 413284
rect 362276 413244 362282 413256
rect 436738 413244 436744 413256
rect 436796 413244 436802 413296
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 439498 403016 439504 403028
rect 361632 402988 439504 403016
rect 361632 402976 361638 402988
rect 439498 402976 439504 402988
rect 439556 402976 439562 403028
rect 502610 402228 502616 402280
rect 502668 402268 502674 402280
rect 557534 402268 557540 402280
rect 502668 402240 557540 402268
rect 502668 402228 502674 402240
rect 557534 402228 557540 402240
rect 557592 402228 557598 402280
rect 497458 400868 497464 400920
rect 497516 400908 497522 400920
rect 546494 400908 546500 400920
rect 497516 400880 546500 400908
rect 497516 400868 497522 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 494146 399440 494152 399492
rect 494204 399480 494210 399492
rect 539594 399480 539600 399492
rect 494204 399452 539600 399480
rect 494204 399440 494210 399452
rect 539594 399440 539600 399452
rect 539652 399440 539658 399492
rect 492674 398080 492680 398132
rect 492732 398120 492738 398132
rect 538214 398120 538220 398132
rect 492732 398092 538220 398120
rect 492732 398080 492738 398092
rect 538214 398080 538220 398092
rect 538272 398080 538278 398132
rect 492766 396720 492772 396772
rect 492824 396760 492830 396772
rect 536834 396760 536840 396772
rect 492824 396732 536840 396760
rect 492824 396720 492830 396732
rect 536834 396720 536840 396732
rect 536892 396720 536898 396772
rect 460934 395292 460940 395344
rect 460992 395332 460998 395344
rect 490006 395332 490012 395344
rect 460992 395304 490012 395332
rect 460992 395292 460998 395304
rect 490006 395292 490012 395304
rect 490064 395292 490070 395344
rect 491570 395292 491576 395344
rect 491628 395332 491634 395344
rect 535454 395332 535460 395344
rect 491628 395304 535460 395332
rect 491628 395292 491634 395304
rect 535454 395292 535460 395304
rect 535512 395292 535518 395344
rect 461026 393932 461032 393984
rect 461084 393972 461090 393984
rect 486418 393972 486424 393984
rect 461084 393944 486424 393972
rect 461084 393932 461090 393944
rect 486418 393932 486424 393944
rect 486476 393932 486482 393984
rect 491386 393932 491392 393984
rect 491444 393972 491450 393984
rect 534166 393972 534172 393984
rect 491444 393944 534172 393972
rect 491444 393932 491450 393944
rect 534166 393932 534172 393944
rect 534224 393932 534230 393984
rect 463602 392572 463608 392624
rect 463660 392612 463666 392624
rect 481634 392612 481640 392624
rect 463660 392584 481640 392612
rect 463660 392572 463666 392584
rect 481634 392572 481640 392584
rect 481692 392572 481698 392624
rect 490558 392572 490564 392624
rect 490616 392612 490622 392624
rect 534074 392612 534080 392624
rect 490616 392584 534080 392612
rect 490616 392572 490622 392584
rect 534074 392572 534080 392584
rect 534132 392572 534138 392624
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 440970 392000 440976 392012
rect 361632 391972 440976 392000
rect 361632 391960 361638 391972
rect 440970 391960 440976 391972
rect 441028 391960 441034 392012
rect 450078 391280 450084 391332
rect 450136 391320 450142 391332
rect 491110 391320 491116 391332
rect 450136 391292 491116 391320
rect 450136 391280 450142 391292
rect 491110 391280 491116 391292
rect 491168 391280 491174 391332
rect 496446 391280 496452 391332
rect 496504 391320 496510 391332
rect 543734 391320 543740 391332
rect 496504 391292 543740 391320
rect 496504 391280 496510 391292
rect 543734 391280 543740 391292
rect 543792 391280 543798 391332
rect 422386 391212 422392 391264
rect 422444 391252 422450 391264
rect 506014 391252 506020 391264
rect 422444 391224 506020 391252
rect 422444 391212 422450 391224
rect 506014 391212 506020 391224
rect 506072 391212 506078 391264
rect 460382 389852 460388 389904
rect 460440 389892 460446 389904
rect 479518 389892 479524 389904
rect 460440 389864 479524 389892
rect 460440 389852 460446 389864
rect 479518 389852 479524 389864
rect 479576 389852 479582 389904
rect 495710 389852 495716 389904
rect 495768 389892 495774 389904
rect 542354 389892 542360 389904
rect 495768 389864 542360 389892
rect 495768 389852 495774 389864
rect 542354 389852 542360 389864
rect 542412 389852 542418 389904
rect 422294 389784 422300 389836
rect 422352 389824 422358 389836
rect 505278 389824 505284 389836
rect 422352 389796 505284 389824
rect 422352 389784 422358 389796
rect 505278 389784 505284 389796
rect 505336 389784 505342 389836
rect 449986 389240 449992 389292
rect 450044 389280 450050 389292
rect 450722 389280 450728 389292
rect 450044 389252 450728 389280
rect 450044 389240 450050 389252
rect 450722 389240 450728 389252
rect 450780 389240 450786 389292
rect 454034 389240 454040 389292
rect 454092 389280 454098 389292
rect 454862 389280 454868 389292
rect 454092 389252 454868 389280
rect 454092 389240 454098 389252
rect 454862 389240 454868 389252
rect 454920 389240 454926 389292
rect 460934 389240 460940 389292
rect 460992 389280 460998 389292
rect 461486 389280 461492 389292
rect 460992 389252 461492 389280
rect 460992 389240 460998 389252
rect 461486 389240 461492 389252
rect 461544 389240 461550 389292
rect 483014 389240 483020 389292
rect 483072 389280 483078 389292
rect 483566 389280 483572 389292
rect 483072 389252 483572 389280
rect 483072 389240 483078 389252
rect 483566 389240 483572 389252
rect 483624 389240 483630 389292
rect 492674 389240 492680 389292
rect 492732 389280 492738 389292
rect 493134 389280 493140 389292
rect 492732 389252 493140 389280
rect 492732 389240 492738 389252
rect 493134 389240 493140 389252
rect 493192 389240 493198 389292
rect 494054 389240 494060 389292
rect 494112 389280 494118 389292
rect 494606 389280 494612 389292
rect 494112 389252 494612 389280
rect 494112 389240 494118 389252
rect 494606 389240 494612 389252
rect 494664 389240 494670 389292
rect 507854 389240 507860 389292
rect 507912 389280 507918 389292
rect 508590 389280 508596 389292
rect 507912 389252 508596 389280
rect 507912 389240 507918 389252
rect 508590 389240 508596 389252
rect 508648 389240 508654 389292
rect 453758 389104 453764 389156
rect 453816 389144 453822 389156
rect 454678 389144 454684 389156
rect 453816 389116 454684 389144
rect 453816 389104 453822 389116
rect 454678 389104 454684 389116
rect 454736 389104 454742 389156
rect 456702 389104 456708 389156
rect 456760 389144 456766 389156
rect 457438 389144 457444 389156
rect 456760 389116 457444 389144
rect 456760 389104 456766 389116
rect 457438 389104 457444 389116
rect 457496 389104 457502 389156
rect 468570 389104 468576 389156
rect 468628 389144 468634 389156
rect 469214 389144 469220 389156
rect 468628 389116 469220 389144
rect 468628 389104 468634 389116
rect 469214 389104 469220 389116
rect 469272 389104 469278 389156
rect 469858 388900 469864 388952
rect 469916 388940 469922 388952
rect 478046 388940 478052 388952
rect 469916 388912 478052 388940
rect 469916 388900 469922 388912
rect 478046 388900 478052 388912
rect 478104 388900 478110 388952
rect 484670 388900 484676 388952
rect 484728 388940 484734 388952
rect 502978 388940 502984 388952
rect 484728 388912 502984 388940
rect 484728 388900 484734 388912
rect 502978 388900 502984 388912
rect 503036 388900 503042 388952
rect 499390 388832 499396 388884
rect 499448 388872 499454 388884
rect 522298 388872 522304 388884
rect 499448 388844 522304 388872
rect 499448 388832 499454 388844
rect 522298 388832 522304 388844
rect 522356 388832 522362 388884
rect 468478 388764 468484 388816
rect 468536 388804 468542 388816
rect 478782 388804 478788 388816
rect 468536 388776 478788 388804
rect 468536 388764 468542 388776
rect 478782 388764 478788 388776
rect 478840 388764 478846 388816
rect 500862 388764 500868 388816
rect 500920 388804 500926 388816
rect 523678 388804 523684 388816
rect 500920 388776 523684 388804
rect 500920 388764 500926 388776
rect 523678 388764 523684 388776
rect 523736 388764 523742 388816
rect 459646 388696 459652 388748
rect 459704 388736 459710 388748
rect 463602 388736 463608 388748
rect 459704 388708 463608 388736
rect 459704 388696 459710 388708
rect 463602 388696 463608 388708
rect 463660 388696 463666 388748
rect 468754 388696 468760 388748
rect 468812 388736 468818 388748
rect 480254 388736 480260 388748
rect 468812 388708 480260 388736
rect 468812 388696 468818 388708
rect 480254 388696 480260 388708
rect 480312 388696 480318 388748
rect 502334 388696 502340 388748
rect 502392 388736 502398 388748
rect 526438 388736 526444 388748
rect 502392 388708 526444 388736
rect 502392 388696 502398 388708
rect 526438 388696 526444 388708
rect 526496 388696 526502 388748
rect 461670 388628 461676 388680
rect 461728 388668 461734 388680
rect 468478 388668 468484 388680
rect 461728 388640 468484 388668
rect 461728 388628 461734 388640
rect 468478 388628 468484 388640
rect 468536 388628 468542 388680
rect 468662 388628 468668 388680
rect 468720 388668 468726 388680
rect 482462 388668 482468 388680
rect 468720 388640 482468 388668
rect 468720 388628 468726 388640
rect 482462 388628 482468 388640
rect 482520 388628 482526 388680
rect 485406 388628 485412 388680
rect 485464 388668 485470 388680
rect 524414 388668 524420 388680
rect 485464 388640 524420 388668
rect 485464 388628 485470 388640
rect 524414 388628 524420 388640
rect 524472 388628 524478 388680
rect 461578 388560 461584 388612
rect 461636 388600 461642 388612
rect 476574 388600 476580 388612
rect 461636 388572 476580 388600
rect 461636 388560 461642 388572
rect 476574 388560 476580 388572
rect 476632 388560 476638 388612
rect 486878 388560 486884 388612
rect 486936 388600 486942 388612
rect 527174 388600 527180 388612
rect 486936 388572 527180 388600
rect 486936 388560 486942 388572
rect 527174 388560 527180 388572
rect 527232 388560 527238 388612
rect 465718 388492 465724 388544
rect 465776 388532 465782 388544
rect 481726 388532 481732 388544
rect 465776 388504 481732 388532
rect 465776 388492 465782 388504
rect 481726 388492 481732 388504
rect 481784 388492 481790 388544
rect 489822 388492 489828 388544
rect 489880 388532 489886 388544
rect 530578 388532 530584 388544
rect 489880 388504 530584 388532
rect 489880 388492 489886 388504
rect 530578 388492 530584 388504
rect 530636 388492 530642 388544
rect 448422 388424 448428 388476
rect 448480 388464 448486 388476
rect 461762 388464 461768 388476
rect 448480 388436 461768 388464
rect 448480 388424 448486 388436
rect 461762 388424 461768 388436
rect 461820 388424 461826 388476
rect 464338 388424 464344 388476
rect 464396 388464 464402 388476
rect 480990 388464 480996 388476
rect 464396 388436 480996 388464
rect 464396 388424 464402 388436
rect 480990 388424 480996 388436
rect 481048 388424 481054 388476
rect 488350 388424 488356 388476
rect 488408 388464 488414 388476
rect 529198 388464 529204 388476
rect 488408 388436 529204 388464
rect 488408 388424 488414 388436
rect 529198 388424 529204 388436
rect 529256 388424 529262 388476
rect 462958 388152 462964 388204
rect 463016 388192 463022 388204
rect 469950 388192 469956 388204
rect 463016 388164 469956 388192
rect 463016 388152 463022 388164
rect 469950 388152 469956 388164
rect 470008 388152 470014 388204
rect 466454 387744 466460 387796
rect 466512 387784 466518 387796
rect 467374 387784 467380 387796
rect 466512 387756 467380 387784
rect 466512 387744 466518 387756
rect 467374 387744 467380 387756
rect 467432 387744 467438 387796
rect 450262 387132 450268 387184
rect 450320 387172 450326 387184
rect 491294 387172 491300 387184
rect 450320 387144 491300 387172
rect 450320 387132 450326 387144
rect 491294 387132 491300 387144
rect 491352 387132 491358 387184
rect 449158 387064 449164 387116
rect 449216 387104 449222 387116
rect 513374 387104 513380 387116
rect 449216 387076 513380 387104
rect 449216 387064 449222 387076
rect 513374 387064 513380 387076
rect 513432 387064 513438 387116
rect 447870 386588 447876 386640
rect 447928 386628 447934 386640
rect 553946 386628 553952 386640
rect 447928 386600 553952 386628
rect 447928 386588 447934 386600
rect 553946 386588 553952 386600
rect 554004 386588 554010 386640
rect 382918 386520 382924 386572
rect 382976 386560 382982 386572
rect 512178 386560 512184 386572
rect 382976 386532 512184 386560
rect 382976 386520 382982 386532
rect 512178 386520 512184 386532
rect 512236 386520 512242 386572
rect 380250 386452 380256 386504
rect 380308 386492 380314 386504
rect 512270 386492 512276 386504
rect 380308 386464 512276 386492
rect 380308 386452 380314 386464
rect 512270 386452 512276 386464
rect 512328 386452 512334 386504
rect 380158 386384 380164 386436
rect 380216 386424 380222 386436
rect 511994 386424 512000 386436
rect 380216 386396 512000 386424
rect 380216 386384 380222 386396
rect 511994 386384 512000 386396
rect 512052 386384 512058 386436
rect 447778 385976 447784 386028
rect 447836 386016 447842 386028
rect 451918 386016 451924 386028
rect 447836 385988 451924 386016
rect 447836 385976 447842 385988
rect 451918 385976 451924 385988
rect 451976 385976 451982 386028
rect 447594 385364 447600 385416
rect 447652 385404 447658 385416
rect 453298 385404 453304 385416
rect 447652 385376 453304 385404
rect 447652 385364 447658 385376
rect 453298 385364 453304 385376
rect 453356 385364 453362 385416
rect 447686 385092 447692 385144
rect 447744 385132 447750 385144
rect 563422 385132 563428 385144
rect 447744 385104 563428 385132
rect 447744 385092 447750 385104
rect 563422 385092 563428 385104
rect 563480 385092 563486 385144
rect 374638 385024 374644 385076
rect 374696 385064 374702 385076
rect 512086 385064 512092 385076
rect 374696 385036 512092 385064
rect 374696 385024 374702 385036
rect 512086 385024 512092 385036
rect 512144 385024 512150 385076
rect 364978 384956 364984 385008
rect 365036 384996 365042 385008
rect 447134 384996 447140 385008
rect 365036 384968 447140 384996
rect 365036 384956 365042 384968
rect 447134 384956 447140 384968
rect 447192 384956 447198 385008
rect 512730 383732 512736 383784
rect 512788 383772 512794 383784
rect 534718 383772 534724 383784
rect 512788 383744 534724 383772
rect 512788 383732 512794 383744
rect 534718 383732 534724 383744
rect 534776 383732 534782 383784
rect 513282 383664 513288 383716
rect 513340 383704 513346 383716
rect 548518 383704 548524 383716
rect 513340 383676 548524 383704
rect 513340 383664 513346 383676
rect 548518 383664 548524 383676
rect 548576 383664 548582 383716
rect 381538 383596 381544 383648
rect 381596 383636 381602 383648
rect 447134 383636 447140 383648
rect 381596 383608 447140 383636
rect 381596 383596 381602 383608
rect 447134 383596 447140 383608
rect 447192 383596 447198 383648
rect 406378 383528 406384 383580
rect 406436 383568 406442 383580
rect 447226 383568 447232 383580
rect 406436 383540 447232 383568
rect 406436 383528 406442 383540
rect 447226 383528 447232 383540
rect 447284 383528 447290 383580
rect 513190 382440 513196 382492
rect 513248 382480 513254 382492
rect 518342 382480 518348 382492
rect 513248 382452 518348 382480
rect 513248 382440 513254 382452
rect 518342 382440 518348 382452
rect 518400 382440 518406 382492
rect 513282 382372 513288 382424
rect 513340 382412 513346 382424
rect 519630 382412 519636 382424
rect 513340 382384 519636 382412
rect 513340 382372 513346 382384
rect 519630 382372 519636 382384
rect 519688 382372 519694 382424
rect 512914 382236 512920 382288
rect 512972 382276 512978 382288
rect 522298 382276 522304 382288
rect 512972 382248 522304 382276
rect 512972 382236 512978 382248
rect 522298 382236 522304 382248
rect 522356 382236 522362 382288
rect 378778 382168 378784 382220
rect 378836 382208 378842 382220
rect 447134 382208 447140 382220
rect 378836 382180 447140 382208
rect 378836 382168 378842 382180
rect 447134 382168 447140 382180
rect 447192 382168 447198 382220
rect 407758 382100 407764 382152
rect 407816 382140 407822 382152
rect 447226 382140 447232 382152
rect 407816 382112 447232 382140
rect 407816 382100 407822 382112
rect 447226 382100 447232 382112
rect 447284 382100 447290 382152
rect 512362 381080 512368 381132
rect 512420 381120 512426 381132
rect 515490 381120 515496 381132
rect 512420 381092 515496 381120
rect 512420 381080 512426 381092
rect 515490 381080 515496 381092
rect 515548 381080 515554 381132
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 442350 380916 442356 380928
rect 361632 380888 442356 380916
rect 361632 380876 361638 380888
rect 442350 380876 442356 380888
rect 442408 380876 442414 380928
rect 513282 380876 513288 380928
rect 513340 380916 513346 380928
rect 548610 380916 548616 380928
rect 513340 380888 548616 380916
rect 513340 380876 513346 380888
rect 548610 380876 548616 380888
rect 548668 380876 548674 380928
rect 376018 380808 376024 380860
rect 376076 380848 376082 380860
rect 447134 380848 447140 380860
rect 376076 380820 447140 380848
rect 376076 380808 376082 380820
rect 447134 380808 447140 380820
rect 447192 380808 447198 380860
rect 410518 380740 410524 380792
rect 410576 380780 410582 380792
rect 447226 380780 447232 380792
rect 410576 380752 447232 380780
rect 410576 380740 410582 380752
rect 447226 380740 447232 380752
rect 447284 380740 447290 380792
rect 512086 380400 512092 380452
rect 512144 380440 512150 380452
rect 512454 380440 512460 380452
rect 512144 380412 512460 380440
rect 512144 380400 512150 380412
rect 512454 380400 512460 380412
rect 512512 380400 512518 380452
rect 512086 380128 512092 380180
rect 512144 380168 512150 380180
rect 514110 380168 514116 380180
rect 512144 380140 514116 380168
rect 512144 380128 512150 380140
rect 514110 380128 514116 380140
rect 514168 380128 514174 380180
rect 512822 379516 512828 379568
rect 512880 379556 512886 379568
rect 544378 379556 544384 379568
rect 512880 379528 544384 379556
rect 512880 379516 512886 379528
rect 544378 379516 544384 379528
rect 544436 379516 544442 379568
rect 371878 379448 371884 379500
rect 371936 379488 371942 379500
rect 447226 379488 447232 379500
rect 371936 379460 447232 379488
rect 371936 379448 371942 379460
rect 447226 379448 447232 379460
rect 447284 379448 447290 379500
rect 374730 379380 374736 379432
rect 374788 379420 374794 379432
rect 447134 379420 447140 379432
rect 374788 379392 447140 379420
rect 374788 379380 374794 379392
rect 447134 379380 447140 379392
rect 447192 379380 447198 379432
rect 512178 378292 512184 378344
rect 512236 378332 512242 378344
rect 523678 378332 523684 378344
rect 512236 378304 523684 378332
rect 512236 378292 512242 378304
rect 523678 378292 523684 378304
rect 523736 378292 523742 378344
rect 513282 378224 513288 378276
rect 513340 378264 513346 378276
rect 547138 378264 547144 378276
rect 513340 378236 547144 378264
rect 513340 378224 513346 378236
rect 547138 378224 547144 378236
rect 547196 378224 547202 378276
rect 514018 378156 514024 378208
rect 514076 378196 514082 378208
rect 579614 378196 579620 378208
rect 514076 378168 579620 378196
rect 514076 378156 514082 378168
rect 579614 378156 579620 378168
rect 579672 378156 579678 378208
rect 367738 378088 367744 378140
rect 367796 378128 367802 378140
rect 447226 378128 447232 378140
rect 367796 378100 447232 378128
rect 367796 378088 367802 378100
rect 447226 378088 447232 378100
rect 447284 378088 447290 378140
rect 370498 378020 370504 378072
rect 370556 378060 370562 378072
rect 447134 378060 447140 378072
rect 370556 378032 447140 378060
rect 370556 378020 370562 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 513190 376864 513196 376916
rect 513248 376904 513254 376916
rect 517514 376904 517520 376916
rect 513248 376876 517520 376904
rect 513248 376864 513254 376876
rect 517514 376864 517520 376876
rect 517572 376864 517578 376916
rect 363690 376660 363696 376712
rect 363748 376700 363754 376712
rect 447226 376700 447232 376712
rect 363748 376672 447232 376700
rect 363748 376660 363754 376672
rect 447226 376660 447232 376672
rect 447284 376660 447290 376712
rect 363598 376592 363604 376644
rect 363656 376632 363662 376644
rect 447134 376632 447140 376644
rect 363656 376604 447140 376632
rect 363656 376592 363662 376604
rect 447134 376592 447140 376604
rect 447192 376592 447198 376644
rect 512362 375980 512368 376032
rect 512420 376020 512426 376032
rect 549898 376020 549904 376032
rect 512420 375992 549904 376020
rect 512420 375980 512426 375992
rect 549898 375980 549904 375992
rect 549956 375980 549962 376032
rect 363782 375300 363788 375352
rect 363840 375340 363846 375352
rect 447134 375340 447140 375352
rect 363840 375312 447140 375340
rect 363840 375300 363846 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 411898 375232 411904 375284
rect 411956 375272 411962 375284
rect 447226 375272 447232 375284
rect 411956 375244 447232 375272
rect 411956 375232 411962 375244
rect 447226 375232 447232 375244
rect 447284 375232 447290 375284
rect 512730 374144 512736 374196
rect 512788 374184 512794 374196
rect 516134 374184 516140 374196
rect 512788 374156 516140 374184
rect 512788 374144 512794 374156
rect 516134 374144 516140 374156
rect 516192 374144 516198 374196
rect 414658 373940 414664 373992
rect 414716 373980 414722 373992
rect 447134 373980 447140 373992
rect 414716 373952 447140 373980
rect 414716 373940 414722 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 416130 373872 416136 373924
rect 416188 373912 416194 373924
rect 447226 373912 447232 373924
rect 416188 373884 447232 373912
rect 416188 373872 416194 373884
rect 447226 373872 447232 373884
rect 447284 373872 447290 373924
rect 512822 372648 512828 372700
rect 512880 372688 512886 372700
rect 517606 372688 517612 372700
rect 512880 372660 517612 372688
rect 512880 372648 512886 372660
rect 517606 372648 517612 372660
rect 517664 372648 517670 372700
rect 513282 372580 513288 372632
rect 513340 372620 513346 372632
rect 521654 372620 521660 372632
rect 513340 372592 521660 372620
rect 513340 372580 513346 372592
rect 521654 372580 521660 372592
rect 521712 372580 521718 372632
rect 417418 372512 417424 372564
rect 417476 372552 417482 372564
rect 447134 372552 447140 372564
rect 417476 372524 447140 372552
rect 417476 372512 417482 372524
rect 447134 372512 447140 372524
rect 447192 372512 447198 372564
rect 419074 372444 419080 372496
rect 419132 372484 419138 372496
rect 447226 372484 447232 372496
rect 419132 372456 447232 372484
rect 419132 372444 419138 372456
rect 447226 372444 447232 372456
rect 447284 372444 447290 372496
rect 512546 371220 512552 371272
rect 512604 371260 512610 371272
rect 517698 371260 517704 371272
rect 512604 371232 517704 371260
rect 512604 371220 512610 371232
rect 517698 371220 517704 371232
rect 517756 371220 517762 371272
rect 383010 371152 383016 371204
rect 383068 371192 383074 371204
rect 447226 371192 447232 371204
rect 383068 371164 447232 371192
rect 383068 371152 383074 371164
rect 447226 371152 447232 371164
rect 447284 371152 447290 371204
rect 436738 371084 436744 371136
rect 436796 371124 436802 371136
rect 447134 371124 447140 371136
rect 436796 371096 447140 371124
rect 436796 371084 436802 371096
rect 447134 371084 447140 371096
rect 447192 371084 447198 371136
rect 511994 370064 512000 370116
rect 512052 370104 512058 370116
rect 514202 370104 514208 370116
rect 512052 370076 514208 370104
rect 512052 370064 512058 370076
rect 514202 370064 514208 370076
rect 514260 370064 514266 370116
rect 513282 369996 513288 370048
rect 513340 370036 513346 370048
rect 521746 370036 521752 370048
rect 513340 370008 521752 370036
rect 513340 369996 513346 370008
rect 521746 369996 521752 370008
rect 521804 369996 521810 370048
rect 512086 369928 512092 369980
rect 512144 369968 512150 369980
rect 514938 369968 514944 369980
rect 512144 369940 514944 369968
rect 512144 369928 512150 369940
rect 514938 369928 514944 369940
rect 514996 369928 515002 369980
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 444006 369900 444012 369912
rect 361632 369872 444012 369900
rect 361632 369860 361638 369872
rect 444006 369860 444012 369872
rect 444064 369860 444070 369912
rect 419166 369792 419172 369844
rect 419224 369832 419230 369844
rect 447226 369832 447232 369844
rect 419224 369804 447232 369832
rect 419224 369792 419230 369804
rect 447226 369792 447232 369804
rect 447284 369792 447290 369844
rect 440878 369724 440884 369776
rect 440936 369764 440942 369776
rect 447134 369764 447140 369776
rect 440936 369736 447140 369764
rect 440936 369724 440942 369736
rect 447134 369724 447140 369736
rect 447192 369724 447198 369776
rect 513006 368568 513012 368620
rect 513064 368608 513070 368620
rect 518894 368608 518900 368620
rect 513064 368580 518900 368608
rect 513064 368568 513070 368580
rect 518894 368568 518900 368580
rect 518952 368568 518958 368620
rect 443638 368432 443644 368484
rect 443696 368472 443702 368484
rect 447134 368472 447140 368484
rect 443696 368444 447140 368472
rect 443696 368432 443702 368444
rect 447134 368432 447140 368444
rect 447192 368432 447198 368484
rect 442258 368364 442264 368416
rect 442316 368404 442322 368416
rect 447226 368404 447232 368416
rect 442316 368376 447232 368404
rect 442316 368364 442322 368376
rect 447226 368364 447232 368376
rect 447284 368364 447290 368416
rect 512638 367208 512644 367260
rect 512696 367248 512702 367260
rect 520274 367248 520280 367260
rect 512696 367220 520280 367248
rect 512696 367208 512702 367220
rect 520274 367208 520280 367220
rect 520332 367208 520338 367260
rect 439498 367004 439504 367056
rect 439556 367044 439562 367056
rect 447134 367044 447140 367056
rect 439556 367016 447140 367044
rect 439556 367004 439562 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 440970 366936 440976 366988
rect 441028 366976 441034 366988
rect 447226 366976 447232 366988
rect 441028 366948 447232 366976
rect 441028 366936 441034 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 512454 365848 512460 365900
rect 512512 365888 512518 365900
rect 515582 365888 515588 365900
rect 512512 365860 515588 365888
rect 512512 365848 512518 365860
rect 515582 365848 515588 365860
rect 515640 365848 515646 365900
rect 444006 365644 444012 365696
rect 444064 365684 444070 365696
rect 447134 365684 447140 365696
rect 444064 365656 447140 365684
rect 444064 365644 444070 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 442350 365576 442356 365628
rect 442408 365616 442414 365628
rect 447226 365616 447232 365628
rect 442408 365588 447232 365616
rect 442408 365576 442414 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 512086 364488 512092 364540
rect 512144 364528 512150 364540
rect 514846 364528 514852 364540
rect 512144 364500 514852 364528
rect 512144 364488 512150 364500
rect 514846 364488 514852 364500
rect 514904 364488 514910 364540
rect 570598 364352 570604 364404
rect 570656 364392 570662 364404
rect 580166 364392 580172 364404
rect 570656 364364 580172 364392
rect 570656 364352 570662 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 513282 363060 513288 363112
rect 513340 363100 513346 363112
rect 518250 363100 518256 363112
rect 513340 363072 518256 363100
rect 513340 363060 513346 363072
rect 518250 363060 518256 363072
rect 518308 363060 518314 363112
rect 442258 362992 442264 363044
rect 442316 363032 442322 363044
rect 447226 363032 447232 363044
rect 442316 363004 447232 363032
rect 442316 362992 442322 363004
rect 447226 362992 447232 363004
rect 447284 362992 447290 363044
rect 511994 362992 512000 363044
rect 512052 363032 512058 363044
rect 515030 363032 515036 363044
rect 512052 363004 515036 363032
rect 512052 362992 512058 363004
rect 515030 362992 515036 363004
rect 515088 362992 515094 363044
rect 432598 362924 432604 362976
rect 432656 362964 432662 362976
rect 447134 362964 447140 362976
rect 432656 362936 447140 362964
rect 432656 362924 432662 362936
rect 447134 362924 447140 362936
rect 447192 362924 447198 362976
rect 511994 362176 512000 362228
rect 512052 362216 512058 362228
rect 513742 362216 513748 362228
rect 512052 362188 513748 362216
rect 512052 362176 512058 362188
rect 513742 362176 513748 362188
rect 513800 362176 513806 362228
rect 513282 362040 513288 362092
rect 513340 362080 513346 362092
rect 518986 362080 518992 362092
rect 513340 362052 518992 362080
rect 513340 362040 513346 362052
rect 518986 362040 518992 362052
rect 519044 362040 519050 362092
rect 513098 361768 513104 361820
rect 513156 361808 513162 361820
rect 516870 361808 516876 361820
rect 513156 361780 516876 361808
rect 513156 361768 513162 361780
rect 516870 361768 516876 361780
rect 516928 361768 516934 361820
rect 443638 361632 443644 361684
rect 443696 361672 443702 361684
rect 447226 361672 447232 361684
rect 443696 361644 447232 361672
rect 443696 361632 443702 361644
rect 447226 361632 447232 361644
rect 447284 361632 447290 361684
rect 435450 361564 435456 361616
rect 435508 361604 435514 361616
rect 447134 361604 447140 361616
rect 435508 361576 447140 361604
rect 435508 361564 435514 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 442442 360272 442448 360324
rect 442500 360312 442506 360324
rect 447226 360312 447232 360324
rect 442500 360284 447232 360312
rect 442500 360272 442506 360284
rect 447226 360272 447232 360284
rect 447284 360272 447290 360324
rect 513282 360272 513288 360324
rect 513340 360312 513346 360324
rect 520366 360312 520372 360324
rect 513340 360284 520372 360312
rect 513340 360272 513346 360284
rect 520366 360272 520372 360284
rect 520424 360272 520430 360324
rect 439590 360204 439596 360256
rect 439648 360244 439654 360256
rect 447134 360244 447140 360256
rect 439648 360216 447140 360244
rect 439648 360204 439654 360216
rect 447134 360204 447140 360216
rect 447192 360204 447198 360256
rect 547138 359184 547144 359236
rect 547196 359224 547202 359236
rect 552290 359224 552296 359236
rect 547196 359196 552296 359224
rect 547196 359184 547202 359196
rect 552290 359184 552296 359196
rect 552348 359184 552354 359236
rect 548610 359116 548616 359168
rect 548668 359156 548674 359168
rect 558178 359156 558184 359168
rect 548668 359128 558184 359156
rect 548668 359116 548674 359128
rect 558178 359116 558184 359128
rect 558236 359116 558242 359168
rect 544378 359048 544384 359100
rect 544436 359088 544442 359100
rect 553762 359088 553768 359100
rect 544436 359060 553768 359088
rect 544436 359048 544442 359060
rect 553762 359048 553768 359060
rect 553820 359048 553826 359100
rect 548518 358980 548524 359032
rect 548576 359020 548582 359032
rect 565538 359020 565544 359032
rect 548576 358992 565544 359020
rect 548576 358980 548582 358992
rect 565538 358980 565544 358992
rect 565596 358980 565602 359032
rect 523678 358912 523684 358964
rect 523736 358952 523742 358964
rect 550818 358952 550824 358964
rect 523736 358924 550824 358952
rect 523736 358912 523742 358924
rect 550818 358912 550824 358924
rect 550876 358912 550882 358964
rect 441062 358844 441068 358896
rect 441120 358884 441126 358896
rect 447226 358884 447232 358896
rect 441120 358856 447232 358884
rect 441120 358844 441126 358856
rect 447226 358844 447232 358856
rect 447284 358844 447290 358896
rect 513282 358844 513288 358896
rect 513340 358884 513346 358896
rect 519170 358884 519176 358896
rect 513340 358856 519176 358884
rect 513340 358844 513346 358856
rect 519170 358844 519176 358856
rect 519228 358844 519234 358896
rect 534718 358844 534724 358896
rect 534776 358884 534782 358896
rect 567010 358884 567016 358896
rect 534776 358856 567016 358884
rect 534776 358844 534782 358856
rect 567010 358844 567016 358856
rect 567068 358844 567074 358896
rect 436830 358776 436836 358828
rect 436888 358816 436894 358828
rect 447134 358816 447140 358828
rect 436888 358788 447140 358816
rect 436888 358776 436894 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 514110 358776 514116 358828
rect 514168 358816 514174 358828
rect 555234 358816 555240 358828
rect 514168 358788 555240 358816
rect 514168 358776 514174 358788
rect 555234 358776 555240 358788
rect 555292 358776 555298 358828
rect 549898 358708 549904 358760
rect 549956 358748 549962 358760
rect 556706 358748 556712 358760
rect 549956 358720 556712 358748
rect 549956 358708 549962 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 519630 358640 519636 358692
rect 519688 358680 519694 358692
rect 562594 358680 562600 358692
rect 519688 358652 562600 358680
rect 519688 358640 519694 358652
rect 562594 358640 562600 358652
rect 562652 358640 562658 358692
rect 518342 358572 518348 358624
rect 518400 358612 518406 358624
rect 561122 358612 561128 358624
rect 518400 358584 561128 358612
rect 518400 358572 518406 358584
rect 561122 358572 561128 358584
rect 561180 358572 561186 358624
rect 522298 358504 522304 358556
rect 522356 358544 522362 358556
rect 564066 358544 564072 358556
rect 522356 358516 564072 358544
rect 522356 358504 522362 358516
rect 564066 358504 564072 358516
rect 564124 358504 564130 358556
rect 515490 358436 515496 358488
rect 515548 358476 515554 358488
rect 559650 358476 559656 358488
rect 515548 358448 559656 358476
rect 515548 358436 515554 358448
rect 559650 358436 559656 358448
rect 559708 358436 559714 358488
rect 512086 357620 512092 357672
rect 512144 357660 512150 357672
rect 519262 357660 519268 357672
rect 512144 357632 519268 357660
rect 512144 357620 512150 357632
rect 519262 357620 519268 357632
rect 519320 357620 519326 357672
rect 512086 357416 512092 357468
rect 512144 357456 512150 357468
rect 513834 357456 513840 357468
rect 512144 357428 513840 357456
rect 512144 357416 512150 357428
rect 513834 357416 513840 357428
rect 513892 357416 513898 357468
rect 512086 356328 512092 356380
rect 512144 356368 512150 356380
rect 513650 356368 513656 356380
rect 512144 356340 513656 356368
rect 512144 356328 512150 356340
rect 513650 356328 513656 356340
rect 513708 356328 513714 356380
rect 512730 356124 512736 356176
rect 512788 356164 512794 356176
rect 521838 356164 521844 356176
rect 512788 356136 521844 356164
rect 512788 356124 512794 356136
rect 521838 356124 521844 356136
rect 521896 356124 521902 356176
rect 513282 354764 513288 354816
rect 513340 354804 513346 354816
rect 519446 354804 519452 354816
rect 513340 354776 519452 354804
rect 513340 354764 513346 354776
rect 519446 354764 519452 354776
rect 519504 354764 519510 354816
rect 513190 354696 513196 354748
rect 513248 354736 513254 354748
rect 521930 354736 521936 354748
rect 513248 354708 521936 354736
rect 513248 354696 513254 354708
rect 521930 354696 521936 354708
rect 521988 354696 521994 354748
rect 512086 353744 512092 353796
rect 512144 353784 512150 353796
rect 515122 353784 515128 353796
rect 512144 353756 515128 353784
rect 512144 353744 512150 353756
rect 515122 353744 515128 353756
rect 515180 353744 515186 353796
rect 513282 353268 513288 353320
rect 513340 353308 513346 353320
rect 519078 353308 519084 353320
rect 513340 353280 519084 353308
rect 513340 353268 513346 353280
rect 519078 353268 519084 353280
rect 519136 353268 519142 353320
rect 512914 352112 512920 352164
rect 512972 352152 512978 352164
rect 516318 352152 516324 352164
rect 512972 352124 516324 352152
rect 512972 352112 512978 352124
rect 516318 352112 516324 352124
rect 516376 352112 516382 352164
rect 424318 352044 424324 352096
rect 424376 352084 424382 352096
rect 426894 352084 426900 352096
rect 424376 352056 426900 352084
rect 424376 352044 424382 352056
rect 426894 352044 426900 352056
rect 426952 352044 426958 352096
rect 394694 351908 394700 351960
rect 394752 351948 394758 351960
rect 447134 351948 447140 351960
rect 394752 351920 447140 351948
rect 394752 351908 394758 351920
rect 447134 351908 447140 351920
rect 447192 351908 447198 351960
rect 513282 351908 513288 351960
rect 513340 351948 513346 351960
rect 522022 351948 522028 351960
rect 513340 351920 522028 351948
rect 513340 351908 513346 351920
rect 522022 351908 522028 351920
rect 522080 351908 522086 351960
rect 512822 351432 512828 351484
rect 512880 351472 512886 351484
rect 517882 351472 517888 351484
rect 512880 351444 517888 351472
rect 512880 351432 512886 351444
rect 517882 351432 517888 351444
rect 517940 351432 517946 351484
rect 512086 350752 512092 350804
rect 512144 350792 512150 350804
rect 515214 350792 515220 350804
rect 512144 350764 515220 350792
rect 512144 350752 512150 350764
rect 515214 350752 515220 350764
rect 515272 350752 515278 350804
rect 405734 350548 405740 350600
rect 405792 350588 405798 350600
rect 447134 350588 447140 350600
rect 405792 350560 447140 350588
rect 405792 350548 405798 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 513006 349256 513012 349308
rect 513064 349296 513070 349308
rect 519354 349296 519360 349308
rect 513064 349268 519360 349296
rect 513064 349256 513070 349268
rect 519354 349256 519360 349268
rect 519412 349256 519418 349308
rect 512086 349188 512092 349240
rect 512144 349228 512150 349240
rect 513926 349228 513932 349240
rect 512144 349200 513932 349228
rect 512144 349188 512150 349200
rect 513926 349188 513932 349200
rect 513984 349188 513990 349240
rect 446858 349052 446864 349104
rect 446916 349092 446922 349104
rect 447594 349092 447600 349104
rect 446916 349064 447600 349092
rect 446916 349052 446922 349064
rect 447594 349052 447600 349064
rect 447652 349052 447658 349104
rect 432782 348372 432788 348424
rect 432840 348412 432846 348424
rect 442258 348412 442264 348424
rect 432840 348384 442264 348412
rect 432840 348372 432846 348384
rect 442258 348372 442264 348384
rect 442316 348372 442322 348424
rect 512822 347896 512828 347948
rect 512880 347936 512886 347948
rect 516226 347936 516232 347948
rect 512880 347908 516232 347936
rect 512880 347896 512886 347908
rect 516226 347896 516232 347908
rect 516284 347896 516290 347948
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 402238 347800 402244 347812
rect 361816 347772 402244 347800
rect 361816 347760 361822 347772
rect 402238 347760 402244 347772
rect 402296 347760 402302 347812
rect 512914 347760 512920 347812
rect 512972 347800 512978 347812
rect 516502 347800 516508 347812
rect 512972 347772 516508 347800
rect 512972 347760 512978 347772
rect 516502 347760 516508 347772
rect 516560 347760 516566 347812
rect 362218 347692 362224 347744
rect 362276 347732 362282 347744
rect 447134 347732 447140 347744
rect 362276 347704 447140 347732
rect 362276 347692 362282 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 426894 347624 426900 347676
rect 426952 347664 426958 347676
rect 430574 347664 430580 347676
rect 426952 347636 430580 347664
rect 426952 347624 426958 347636
rect 430574 347624 430580 347636
rect 430632 347624 430638 347676
rect 513282 346672 513288 346724
rect 513340 346712 513346 346724
rect 517790 346712 517796 346724
rect 513340 346684 517796 346712
rect 513340 346672 513346 346684
rect 517790 346672 517796 346684
rect 517848 346672 517854 346724
rect 512822 346536 512828 346588
rect 512880 346576 512886 346588
rect 517974 346576 517980 346588
rect 512880 346548 517980 346576
rect 512880 346536 512886 346548
rect 517974 346536 517980 346548
rect 518032 346536 518038 346588
rect 512638 346400 512644 346452
rect 512696 346440 512702 346452
rect 515306 346440 515312 346452
rect 512696 346412 515312 346440
rect 512696 346400 512702 346412
rect 515306 346400 515312 346412
rect 515364 346400 515370 346452
rect 512086 345924 512092 345976
rect 512144 345964 512150 345976
rect 514110 345964 514116 345976
rect 512144 345936 514116 345964
rect 512144 345924 512150 345936
rect 514110 345924 514116 345936
rect 514168 345924 514174 345976
rect 432782 344292 432788 344344
rect 432840 344332 432846 344344
rect 443638 344332 443644 344344
rect 432840 344304 443644 344332
rect 432840 344292 432846 344304
rect 443638 344292 443644 344304
rect 443696 344292 443702 344344
rect 512638 344224 512644 344276
rect 512696 344264 512702 344276
rect 515490 344264 515496 344276
rect 512696 344236 515496 344264
rect 512696 344224 512702 344236
rect 515490 344224 515496 344236
rect 515548 344224 515554 344276
rect 513282 343952 513288 344004
rect 513340 343992 513346 344004
rect 518066 343992 518072 344004
rect 513340 343964 518072 343992
rect 513340 343952 513346 343964
rect 518066 343952 518072 343964
rect 518124 343952 518130 344004
rect 512822 343816 512828 343868
rect 512880 343856 512886 343868
rect 516410 343856 516416 343868
rect 512880 343828 516416 343856
rect 512880 343816 512886 343828
rect 516410 343816 516416 343828
rect 516468 343816 516474 343868
rect 402238 342864 402244 342916
rect 402296 342904 402302 342916
rect 402974 342904 402980 342916
rect 402296 342876 402980 342904
rect 402296 342864 402302 342876
rect 402974 342864 402980 342876
rect 403032 342904 403038 342916
rect 447870 342904 447876 342916
rect 403032 342876 447876 342904
rect 403032 342864 403038 342876
rect 447870 342864 447876 342876
rect 447928 342864 447934 342916
rect 430574 342184 430580 342236
rect 430632 342224 430638 342236
rect 432690 342224 432696 342236
rect 430632 342196 432696 342224
rect 430632 342184 430638 342196
rect 432690 342184 432696 342196
rect 432748 342184 432754 342236
rect 513282 341232 513288 341284
rect 513340 341272 513346 341284
rect 519630 341272 519636 341284
rect 513340 341244 519636 341272
rect 513340 341232 513346 341244
rect 519630 341232 519636 341244
rect 519688 341232 519694 341284
rect 444098 340960 444104 341012
rect 444156 341000 444162 341012
rect 447226 341000 447232 341012
rect 444156 340972 447232 341000
rect 444156 340960 444162 340972
rect 447226 340960 447232 340972
rect 447284 340960 447290 341012
rect 513006 340960 513012 341012
rect 513064 341000 513070 341012
rect 516594 341000 516600 341012
rect 513064 340972 516600 341000
rect 513064 340960 513070 340972
rect 516594 340960 516600 340972
rect 516652 340960 516658 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447134 340932 447140 340944
rect 361816 340904 447140 340932
rect 361816 340892 361822 340904
rect 447134 340892 447140 340904
rect 447192 340892 447198 340944
rect 513282 339872 513288 339924
rect 513340 339912 513346 339924
rect 520550 339912 520556 339924
rect 513340 339884 520556 339912
rect 513340 339872 513346 339884
rect 520550 339872 520556 339884
rect 520608 339872 520614 339924
rect 442350 339532 442356 339584
rect 442408 339572 442414 339584
rect 447226 339572 447232 339584
rect 442408 339544 447232 339572
rect 442408 339532 442414 339544
rect 447226 339532 447232 339544
rect 447284 339532 447290 339584
rect 513006 339532 513012 339584
rect 513064 339572 513070 339584
rect 516686 339572 516692 339584
rect 513064 339544 516692 339572
rect 513064 339532 513070 339544
rect 516686 339532 516692 339544
rect 516744 339532 516750 339584
rect 399478 339464 399484 339516
rect 399536 339504 399542 339516
rect 447134 339504 447140 339516
rect 399536 339476 447140 339504
rect 399536 339464 399542 339476
rect 447134 339464 447140 339476
rect 447192 339464 447198 339516
rect 513190 339464 513196 339516
rect 513248 339504 513254 339516
rect 522114 339504 522120 339516
rect 513248 339476 522120 339504
rect 513248 339464 513254 339476
rect 522114 339464 522120 339476
rect 522172 339464 522178 339516
rect 401594 339396 401600 339448
rect 401652 339436 401658 339448
rect 402974 339436 402980 339448
rect 401652 339408 402980 339436
rect 401652 339396 401658 339408
rect 402974 339396 402980 339408
rect 403032 339396 403038 339448
rect 412634 338716 412640 338768
rect 412692 338756 412698 338768
rect 449158 338756 449164 338768
rect 412692 338728 449164 338756
rect 412692 338716 412698 338728
rect 449158 338716 449164 338728
rect 449216 338716 449222 338768
rect 513282 338240 513288 338292
rect 513340 338280 513346 338292
rect 519722 338280 519728 338292
rect 513340 338252 519728 338280
rect 513340 338240 513346 338252
rect 519722 338240 519728 338252
rect 519780 338240 519786 338292
rect 435358 338172 435364 338224
rect 435416 338212 435422 338224
rect 447134 338212 447140 338224
rect 435416 338184 447140 338212
rect 435416 338172 435422 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 385770 338104 385776 338156
rect 385828 338144 385834 338156
rect 447226 338144 447232 338156
rect 385828 338116 447232 338144
rect 385828 338104 385834 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 513190 338104 513196 338156
rect 513248 338144 513254 338156
rect 520458 338144 520464 338156
rect 513248 338116 520464 338144
rect 513248 338104 513254 338116
rect 520458 338104 520464 338116
rect 520516 338104 520522 338156
rect 513190 337424 513196 337476
rect 513248 337464 513254 337476
rect 518342 337464 518348 337476
rect 513248 337436 518348 337464
rect 513248 337424 513254 337436
rect 518342 337424 518348 337436
rect 518400 337424 518406 337476
rect 416774 336880 416780 336932
rect 416832 336920 416838 336932
rect 431402 336920 431408 336932
rect 416832 336892 431408 336920
rect 416832 336880 416838 336892
rect 431402 336880 431408 336892
rect 431460 336880 431466 336932
rect 424134 336812 424140 336864
rect 424192 336852 424198 336864
rect 429930 336852 429936 336864
rect 424192 336824 429936 336852
rect 424192 336812 424198 336824
rect 429930 336812 429936 336824
rect 429988 336812 429994 336864
rect 443822 336812 443828 336864
rect 443880 336852 443886 336864
rect 447226 336852 447232 336864
rect 443880 336824 447232 336852
rect 443880 336812 443886 336824
rect 447226 336812 447232 336824
rect 447284 336812 447290 336864
rect 513282 336812 513288 336864
rect 513340 336852 513346 336864
rect 520642 336852 520648 336864
rect 513340 336824 520648 336852
rect 513340 336812 513346 336824
rect 520642 336812 520648 336824
rect 520700 336812 520706 336864
rect 420454 336744 420460 336796
rect 420512 336784 420518 336796
rect 439774 336784 439780 336796
rect 420512 336756 439780 336784
rect 420512 336744 420518 336756
rect 439774 336744 439780 336756
rect 439832 336744 439838 336796
rect 440970 336744 440976 336796
rect 441028 336784 441034 336796
rect 447134 336784 447140 336796
rect 441028 336756 447140 336784
rect 441028 336744 441034 336756
rect 447134 336744 447140 336756
rect 447192 336744 447198 336796
rect 513190 336744 513196 336796
rect 513248 336784 513254 336796
rect 522206 336784 522212 336796
rect 513248 336756 522212 336784
rect 513248 336744 513254 336756
rect 522206 336744 522212 336756
rect 522264 336744 522270 336796
rect 432690 336676 432696 336728
rect 432748 336716 432754 336728
rect 433978 336716 433984 336728
rect 432748 336688 433984 336716
rect 432748 336676 432754 336688
rect 433978 336676 433984 336688
rect 434036 336676 434042 336728
rect 418982 336268 418988 336320
rect 419040 336308 419046 336320
rect 442534 336308 442540 336320
rect 419040 336280 442540 336308
rect 419040 336268 419046 336280
rect 442534 336268 442540 336280
rect 442592 336268 442598 336320
rect 416038 336200 416044 336252
rect 416096 336240 416102 336252
rect 439682 336240 439688 336252
rect 416096 336212 439688 336240
rect 416096 336200 416102 336212
rect 439682 336200 439688 336212
rect 439740 336200 439746 336252
rect 418890 336132 418896 336184
rect 418948 336172 418954 336184
rect 442626 336172 442632 336184
rect 418948 336144 442632 336172
rect 418948 336132 418954 336144
rect 442626 336132 442632 336144
rect 442684 336132 442690 336184
rect 418798 336064 418804 336116
rect 418856 336104 418862 336116
rect 442718 336104 442724 336116
rect 418856 336076 442724 336104
rect 418856 336064 418862 336076
rect 442718 336064 442724 336076
rect 442776 336064 442782 336116
rect 362218 335996 362224 336048
rect 362276 336036 362282 336048
rect 444098 336036 444104 336048
rect 362276 336008 444104 336036
rect 362276 335996 362282 336008
rect 444098 335996 444104 336008
rect 444156 335996 444162 336048
rect 513190 335792 513196 335844
rect 513248 335832 513254 335844
rect 516962 335832 516968 335844
rect 513248 335804 516968 335832
rect 513248 335792 513254 335804
rect 516962 335792 516968 335804
rect 517020 335792 517026 335844
rect 442258 335452 442264 335504
rect 442316 335492 442322 335504
rect 447318 335492 447324 335504
rect 442316 335464 447324 335492
rect 442316 335452 442322 335464
rect 447318 335452 447324 335464
rect 447376 335452 447382 335504
rect 409414 335384 409420 335436
rect 409472 335424 409478 335436
rect 431310 335424 431316 335436
rect 409472 335396 431316 335424
rect 409472 335384 409478 335396
rect 431310 335384 431316 335396
rect 431368 335384 431374 335436
rect 413094 335316 413100 335368
rect 413152 335356 413158 335368
rect 435542 335356 435548 335368
rect 413152 335328 435548 335356
rect 413152 335316 413158 335328
rect 435542 335316 435548 335328
rect 435600 335316 435606 335368
rect 439498 335316 439504 335368
rect 439556 335356 439562 335368
rect 447226 335356 447232 335368
rect 439556 335328 447232 335356
rect 439556 335316 439562 335328
rect 447226 335316 447232 335328
rect 447284 335316 447290 335368
rect 513282 335316 513288 335368
rect 513340 335356 513346 335368
rect 522298 335356 522304 335368
rect 513340 335328 522304 335356
rect 513340 335316 513346 335328
rect 522298 335316 522304 335328
rect 522356 335316 522362 335368
rect 420362 335044 420368 335096
rect 420420 335044 420426 335096
rect 420546 335044 420552 335096
rect 420604 335084 420610 335096
rect 442166 335084 442172 335096
rect 420604 335056 442172 335084
rect 420604 335044 420610 335056
rect 442166 335044 442172 335056
rect 442224 335044 442230 335096
rect 420380 334948 420408 335044
rect 420638 334976 420644 335028
rect 420696 335016 420702 335028
rect 444926 335016 444932 335028
rect 420696 334988 444932 335016
rect 420696 334976 420702 334988
rect 444926 334976 444932 334988
rect 444984 334976 444990 335028
rect 446950 334948 446956 334960
rect 420380 334920 446956 334948
rect 446950 334908 446956 334920
rect 447008 334908 447014 334960
rect 420270 334840 420276 334892
rect 420328 334880 420334 334892
rect 446858 334880 446864 334892
rect 420328 334852 446864 334880
rect 420328 334840 420334 334852
rect 446858 334840 446864 334852
rect 446916 334840 446922 334892
rect 420822 334772 420828 334824
rect 420880 334812 420886 334824
rect 449434 334812 449440 334824
rect 420880 334784 449440 334812
rect 420880 334772 420886 334784
rect 449434 334772 449440 334784
rect 449492 334772 449498 334824
rect 420730 334704 420736 334756
rect 420788 334744 420794 334756
rect 449526 334744 449532 334756
rect 420788 334716 449532 334744
rect 420788 334704 420794 334716
rect 449526 334704 449532 334716
rect 449584 334704 449590 334756
rect 420178 334636 420184 334688
rect 420236 334676 420242 334688
rect 449066 334676 449072 334688
rect 420236 334648 449072 334676
rect 420236 334636 420242 334648
rect 449066 334636 449072 334648
rect 449124 334636 449130 334688
rect 420086 334568 420092 334620
rect 420144 334608 420150 334620
rect 449342 334608 449348 334620
rect 420144 334580 449348 334608
rect 420144 334568 420150 334580
rect 449342 334568 449348 334580
rect 449400 334568 449406 334620
rect 428090 334364 428096 334416
rect 428148 334404 428154 334416
rect 437014 334404 437020 334416
rect 428148 334376 437020 334404
rect 428148 334364 428154 334376
rect 437014 334364 437020 334376
rect 437072 334364 437078 334416
rect 513190 334296 513196 334348
rect 513248 334336 513254 334348
rect 520734 334336 520740 334348
rect 513248 334308 520740 334336
rect 513248 334296 513254 334308
rect 520734 334296 520740 334308
rect 520792 334296 520798 334348
rect 443730 334024 443736 334076
rect 443788 334064 443794 334076
rect 447318 334064 447324 334076
rect 443788 334036 447324 334064
rect 443788 334024 443794 334036
rect 447318 334024 447324 334036
rect 447376 334024 447382 334076
rect 364058 333956 364064 334008
rect 364116 333996 364122 334008
rect 447226 333996 447232 334008
rect 364116 333968 447232 333996
rect 364116 333956 364122 333968
rect 447226 333956 447232 333968
rect 447284 333956 447290 334008
rect 513282 333956 513288 334008
rect 513340 333996 513346 334008
rect 522390 333996 522396 334008
rect 513340 333968 522396 333996
rect 513340 333956 513346 333968
rect 522390 333956 522396 333968
rect 522448 333956 522454 334008
rect 440878 332664 440884 332716
rect 440936 332704 440942 332716
rect 447318 332704 447324 332716
rect 440936 332676 447324 332704
rect 440936 332664 440942 332676
rect 447318 332664 447324 332676
rect 447376 332664 447382 332716
rect 429838 332596 429844 332648
rect 429896 332636 429902 332648
rect 447226 332636 447232 332648
rect 429896 332608 447232 332636
rect 429896 332596 429902 332608
rect 447226 332596 447232 332608
rect 447284 332596 447290 332648
rect 432874 331848 432880 331900
rect 432932 331888 432938 331900
rect 442442 331888 442448 331900
rect 432932 331860 442448 331888
rect 432932 331848 432938 331860
rect 442442 331848 442448 331860
rect 442500 331848 442506 331900
rect 436738 331304 436744 331356
rect 436796 331344 436802 331356
rect 447502 331344 447508 331356
rect 436796 331316 447508 331344
rect 436796 331304 436802 331316
rect 447502 331304 447508 331316
rect 447560 331304 447566 331356
rect 443638 331236 443644 331288
rect 443696 331276 443702 331288
rect 447226 331276 447232 331288
rect 443696 331248 447232 331276
rect 443696 331236 443702 331248
rect 447226 331236 447232 331248
rect 447284 331236 447290 331288
rect 445938 331168 445944 331220
rect 445996 331208 446002 331220
rect 447318 331208 447324 331220
rect 445996 331180 447324 331208
rect 445996 331168 446002 331180
rect 447318 331168 447324 331180
rect 447376 331168 447382 331220
rect 440142 330556 440148 330608
rect 440200 330596 440206 330608
rect 445938 330596 445944 330608
rect 440200 330568 445944 330596
rect 440200 330556 440206 330568
rect 445938 330556 445944 330568
rect 445996 330556 446002 330608
rect 432598 330216 432604 330268
rect 432656 330256 432662 330268
rect 441062 330256 441068 330268
rect 432656 330228 441068 330256
rect 432656 330216 432662 330228
rect 441062 330216 441068 330228
rect 441120 330216 441126 330268
rect 442902 330080 442908 330132
rect 442960 330120 442966 330132
rect 445846 330120 445852 330132
rect 442960 330092 445852 330120
rect 442960 330080 442966 330092
rect 445846 330080 445852 330092
rect 445904 330120 445910 330132
rect 447226 330120 447232 330132
rect 445904 330092 447232 330120
rect 445904 330080 445910 330092
rect 447226 330080 447232 330092
rect 447284 330080 447290 330132
rect 512730 330080 512736 330132
rect 512788 330120 512794 330132
rect 514754 330120 514760 330132
rect 512788 330092 514760 330120
rect 512788 330080 512794 330092
rect 514754 330080 514760 330092
rect 514812 330080 514818 330132
rect 438762 329060 438768 329112
rect 438820 329100 438826 329112
rect 445754 329100 445760 329112
rect 438820 329072 445760 329100
rect 438820 329060 438826 329072
rect 445754 329060 445760 329072
rect 445812 329100 445818 329112
rect 447226 329100 447232 329112
rect 445812 329072 447232 329100
rect 445812 329060 445818 329072
rect 447226 329060 447232 329072
rect 447284 329060 447290 329112
rect 432966 328652 432972 328704
rect 433024 328692 433030 328704
rect 435450 328692 435456 328704
rect 433024 328664 435456 328692
rect 433024 328652 433030 328664
rect 435450 328652 435456 328664
rect 435508 328652 435514 328704
rect 436002 328448 436008 328500
rect 436060 328488 436066 328500
rect 447226 328488 447232 328500
rect 436060 328460 447232 328488
rect 436060 328448 436066 328460
rect 447226 328448 447232 328460
rect 447284 328448 447290 328500
rect 433978 328380 433984 328432
rect 434036 328420 434042 328432
rect 436922 328420 436928 328432
rect 434036 328392 436928 328420
rect 434036 328380 434042 328392
rect 436922 328380 436928 328392
rect 436980 328380 436986 328432
rect 437014 328380 437020 328432
rect 437072 328420 437078 328432
rect 447318 328420 447324 328432
rect 437072 328392 447324 328420
rect 437072 328380 437078 328392
rect 447318 328380 447324 328392
rect 447376 328420 447382 328432
rect 448330 328420 448336 328432
rect 447376 328392 448336 328420
rect 447376 328380 447382 328392
rect 448330 328380 448336 328392
rect 448388 328380 448394 328432
rect 431218 327088 431224 327140
rect 431276 327128 431282 327140
rect 447226 327128 447232 327140
rect 431276 327100 447232 327128
rect 431276 327088 431282 327100
rect 447226 327088 447232 327100
rect 447284 327088 447290 327140
rect 439774 327020 439780 327072
rect 439832 327060 439838 327072
rect 447318 327060 447324 327072
rect 439832 327032 447324 327060
rect 439832 327020 439838 327032
rect 447318 327020 447324 327032
rect 447376 327060 447382 327072
rect 448054 327060 448060 327072
rect 447376 327032 448060 327060
rect 447376 327020 447382 327032
rect 448054 327020 448060 327032
rect 448112 327020 448118 327072
rect 429930 326340 429936 326392
rect 429988 326380 429994 326392
rect 440326 326380 440332 326392
rect 429988 326352 440332 326380
rect 429988 326340 429994 326352
rect 440326 326340 440332 326352
rect 440384 326380 440390 326392
rect 447226 326380 447232 326392
rect 440384 326352 447232 326380
rect 440384 326340 440390 326352
rect 447226 326340 447232 326352
rect 447284 326340 447290 326392
rect 431402 325592 431408 325644
rect 431460 325632 431466 325644
rect 448146 325632 448152 325644
rect 431460 325604 448152 325632
rect 431460 325592 431466 325604
rect 448146 325592 448152 325604
rect 448204 325592 448210 325644
rect 435542 325456 435548 325508
rect 435600 325496 435606 325508
rect 447962 325496 447968 325508
rect 435600 325468 447968 325496
rect 435600 325456 435606 325468
rect 447962 325456 447968 325468
rect 448020 325456 448026 325508
rect 436922 324980 436928 325032
rect 436980 325020 436986 325032
rect 440234 325020 440240 325032
rect 436980 324992 440240 325020
rect 436980 324980 436986 324992
rect 440234 324980 440240 324992
rect 440292 324980 440298 325032
rect 511902 324300 511908 324352
rect 511960 324340 511966 324352
rect 580166 324340 580172 324352
rect 511960 324312 580172 324340
rect 511960 324300 511966 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 440234 323620 440240 323672
rect 440292 323660 440298 323672
rect 447226 323660 447232 323672
rect 440292 323632 447232 323660
rect 440292 323620 440298 323632
rect 447226 323620 447232 323632
rect 447284 323620 447290 323672
rect 431310 323552 431316 323604
rect 431368 323592 431374 323604
rect 449250 323592 449256 323604
rect 431368 323564 449256 323592
rect 431368 323552 431374 323564
rect 449250 323552 449256 323564
rect 449308 323552 449314 323604
rect 510522 323552 510528 323604
rect 510580 323592 510586 323604
rect 580258 323592 580264 323604
rect 510580 323564 580264 323592
rect 510580 323552 510586 323564
rect 580258 323552 580264 323564
rect 580316 323552 580322 323604
rect 507486 322532 507492 322584
rect 507544 322572 507550 322584
rect 509602 322572 509608 322584
rect 507544 322544 509608 322572
rect 507544 322532 507550 322544
rect 509602 322532 509608 322544
rect 509660 322532 509666 322584
rect 442810 322396 442816 322448
rect 442868 322436 442874 322448
rect 449986 322436 449992 322448
rect 442868 322408 449992 322436
rect 442868 322396 442874 322408
rect 449986 322396 449992 322408
rect 450044 322396 450050 322448
rect 446582 322328 446588 322380
rect 446640 322368 446646 322380
rect 470134 322368 470140 322380
rect 446640 322340 470140 322368
rect 446640 322328 446646 322340
rect 470134 322328 470140 322340
rect 470192 322328 470198 322380
rect 446950 322260 446956 322312
rect 447008 322300 447014 322312
rect 483106 322300 483112 322312
rect 447008 322272 483112 322300
rect 447008 322260 447014 322272
rect 483106 322260 483112 322272
rect 483164 322260 483170 322312
rect 447226 322192 447232 322244
rect 447284 322232 447290 322244
rect 449894 322232 449900 322244
rect 447284 322204 449900 322232
rect 447284 322192 447290 322204
rect 449894 322192 449900 322204
rect 449952 322192 449958 322244
rect 449986 322192 449992 322244
rect 450044 322232 450050 322244
rect 479794 322232 479800 322244
rect 450044 322204 479800 322232
rect 450044 322192 450050 322204
rect 479794 322192 479800 322204
rect 479852 322192 479858 322244
rect 507210 322192 507216 322244
rect 507268 322232 507274 322244
rect 514754 322232 514760 322244
rect 507268 322204 514760 322232
rect 507268 322192 507274 322204
rect 514754 322192 514760 322204
rect 514812 322192 514818 322244
rect 445662 322124 445668 322176
rect 445720 322164 445726 322176
rect 471790 322164 471796 322176
rect 445720 322136 471796 322164
rect 445720 322124 445726 322136
rect 471790 322124 471796 322136
rect 471848 322124 471854 322176
rect 477862 322124 477868 322176
rect 477920 322164 477926 322176
rect 514018 322164 514024 322176
rect 477920 322136 514024 322164
rect 477920 322124 477926 322136
rect 514018 322124 514024 322136
rect 514076 322124 514082 322176
rect 444926 322056 444932 322108
rect 444984 322096 444990 322108
rect 482554 322096 482560 322108
rect 444984 322068 482560 322096
rect 444984 322056 444990 322068
rect 482554 322056 482560 322068
rect 482612 322056 482618 322108
rect 504082 322056 504088 322108
rect 504140 322096 504146 322108
rect 511258 322096 511264 322108
rect 504140 322068 511264 322096
rect 504140 322056 504146 322068
rect 511258 322056 511264 322068
rect 511316 322056 511322 322108
rect 439682 321988 439688 322040
rect 439740 322028 439746 322040
rect 470686 322028 470692 322040
rect 439740 322000 470692 322028
rect 439740 321988 439746 322000
rect 470686 321988 470692 322000
rect 470744 321988 470750 322040
rect 478414 321988 478420 322040
rect 478472 322028 478478 322040
rect 518158 322028 518164 322040
rect 478472 322000 518164 322028
rect 478472 321988 478478 322000
rect 518158 321988 518164 322000
rect 518216 321988 518222 322040
rect 450630 321920 450636 321972
rect 450688 321960 450694 321972
rect 460750 321960 460756 321972
rect 450688 321932 460756 321960
rect 450688 321920 450694 321932
rect 460750 321920 460756 321932
rect 460808 321920 460814 321972
rect 467650 321920 467656 321972
rect 467708 321960 467714 321972
rect 467708 321932 504404 321960
rect 467708 321920 467714 321932
rect 446766 321852 446772 321904
rect 446824 321892 446830 321904
rect 461946 321892 461952 321904
rect 446824 321864 461952 321892
rect 446824 321852 446830 321864
rect 461946 321852 461952 321864
rect 462004 321852 462010 321904
rect 468294 321852 468300 321904
rect 468352 321892 468358 321904
rect 504082 321892 504088 321904
rect 468352 321864 504088 321892
rect 468352 321852 468358 321864
rect 504082 321852 504088 321864
rect 504140 321852 504146 321904
rect 504376 321892 504404 321932
rect 507394 321920 507400 321972
rect 507452 321960 507458 321972
rect 509786 321960 509792 321972
rect 507452 321932 509792 321960
rect 507452 321920 507458 321932
rect 509786 321920 509792 321932
rect 509844 321920 509850 321972
rect 509878 321892 509884 321904
rect 504376 321864 509884 321892
rect 509878 321852 509884 321864
rect 509936 321852 509942 321904
rect 442166 321784 442172 321836
rect 442224 321824 442230 321836
rect 462498 321824 462504 321836
rect 442224 321796 462504 321824
rect 442224 321784 442230 321796
rect 462498 321784 462504 321796
rect 462556 321784 462562 321836
rect 467742 321784 467748 321836
rect 467800 321824 467806 321836
rect 516778 321824 516784 321836
rect 467800 321796 516784 321824
rect 467800 321784 467806 321796
rect 516778 321784 516784 321796
rect 516836 321784 516842 321836
rect 457530 321716 457536 321768
rect 457588 321756 457594 321768
rect 567838 321756 567844 321768
rect 457588 321728 567844 321756
rect 457588 321716 457594 321728
rect 567838 321716 567844 321728
rect 567896 321716 567902 321768
rect 458082 321648 458088 321700
rect 458140 321688 458146 321700
rect 580350 321688 580356 321700
rect 458140 321660 580356 321688
rect 458140 321648 458146 321660
rect 580350 321648 580356 321660
rect 580408 321648 580414 321700
rect 457806 321580 457812 321632
rect 457864 321620 457870 321632
rect 580442 321620 580448 321632
rect 457864 321592 580448 321620
rect 457864 321580 457870 321592
rect 580442 321580 580448 321592
rect 580500 321580 580506 321632
rect 456702 321512 456708 321564
rect 456760 321552 456766 321564
rect 580718 321552 580724 321564
rect 456760 321524 580724 321552
rect 456760 321512 456766 321524
rect 580718 321512 580724 321524
rect 580776 321512 580782 321564
rect 456978 321444 456984 321496
rect 457036 321484 457042 321496
rect 580626 321484 580632 321496
rect 457036 321456 580632 321484
rect 457036 321444 457042 321456
rect 580626 321444 580632 321456
rect 580684 321444 580690 321496
rect 458358 321376 458364 321428
rect 458416 321416 458422 321428
rect 569218 321416 569224 321428
rect 458416 321388 569224 321416
rect 458416 321376 458422 321388
rect 569218 321376 569224 321388
rect 569276 321376 569282 321428
rect 445478 321308 445484 321360
rect 445536 321348 445542 321360
rect 461394 321348 461400 321360
rect 445536 321320 461400 321348
rect 445536 321308 445542 321320
rect 461394 321308 461400 321320
rect 461452 321308 461458 321360
rect 468570 321308 468576 321360
rect 468628 321348 468634 321360
rect 576118 321348 576124 321360
rect 468628 321320 576124 321348
rect 468628 321308 468634 321320
rect 576118 321308 576124 321320
rect 576176 321308 576182 321360
rect 445018 321240 445024 321292
rect 445076 321280 445082 321292
rect 459462 321280 459468 321292
rect 445076 321252 459468 321280
rect 445076 321240 445082 321252
rect 459462 321240 459468 321252
rect 459520 321240 459526 321292
rect 467190 321240 467196 321292
rect 467248 321280 467254 321292
rect 570598 321280 570604 321292
rect 467248 321252 570604 321280
rect 467248 321240 467254 321252
rect 570598 321240 570604 321252
rect 570656 321240 570662 321292
rect 446398 321172 446404 321224
rect 446456 321212 446462 321224
rect 459186 321212 459192 321224
rect 446456 321184 459192 321212
rect 446456 321172 446462 321184
rect 459186 321172 459192 321184
rect 459244 321172 459250 321224
rect 477954 321172 477960 321224
rect 478012 321212 478018 321224
rect 574738 321212 574744 321224
rect 478012 321184 574744 321212
rect 478012 321172 478018 321184
rect 574738 321172 574744 321184
rect 574796 321172 574802 321224
rect 479334 321104 479340 321156
rect 479392 321144 479398 321156
rect 573358 321144 573364 321156
rect 479392 321116 573364 321144
rect 479392 321104 479398 321116
rect 573358 321104 573364 321116
rect 573416 321104 573422 321156
rect 445570 321036 445576 321088
rect 445628 321076 445634 321088
rect 461118 321076 461124 321088
rect 445628 321048 461124 321076
rect 445628 321036 445634 321048
rect 461118 321036 461124 321048
rect 461176 321036 461182 321088
rect 468018 321036 468024 321088
rect 468076 321076 468082 321088
rect 511350 321076 511356 321088
rect 468076 321048 511356 321076
rect 468076 321036 468082 321048
rect 511350 321036 511356 321048
rect 511408 321036 511414 321088
rect 450538 320968 450544 321020
rect 450596 321008 450602 321020
rect 481266 321008 481272 321020
rect 450596 320980 481272 321008
rect 450596 320968 450602 320980
rect 481266 320968 481272 320980
rect 481324 320968 481330 321020
rect 507026 320968 507032 321020
rect 507084 321008 507090 321020
rect 516870 321008 516876 321020
rect 507084 320980 516876 321008
rect 507084 320968 507090 320980
rect 516870 320968 516876 320980
rect 516928 320968 516934 321020
rect 445110 320900 445116 320952
rect 445168 320940 445174 320952
rect 460014 320940 460020 320952
rect 445168 320912 460020 320940
rect 445168 320900 445174 320912
rect 460014 320900 460020 320912
rect 460072 320900 460078 320952
rect 460198 320900 460204 320952
rect 460256 320940 460262 320952
rect 518250 320940 518256 320952
rect 460256 320912 518256 320940
rect 460256 320900 460262 320912
rect 518250 320900 518256 320912
rect 518308 320900 518314 320952
rect 449894 320832 449900 320884
rect 449952 320872 449958 320884
rect 456794 320872 456800 320884
rect 449952 320844 456800 320872
rect 449952 320832 449958 320844
rect 456794 320832 456800 320844
rect 456852 320832 456858 320884
rect 459554 320832 459560 320884
rect 459612 320872 459618 320884
rect 580534 320872 580540 320884
rect 459612 320844 580540 320872
rect 459612 320832 459618 320844
rect 580534 320832 580540 320844
rect 580592 320832 580598 320884
rect 446490 320764 446496 320816
rect 446548 320804 446554 320816
rect 480162 320804 480168 320816
rect 446548 320776 480168 320804
rect 446548 320764 446554 320776
rect 480162 320764 480168 320776
rect 480220 320764 480226 320816
rect 507578 320764 507584 320816
rect 507636 320804 507642 320816
rect 513374 320804 513380 320816
rect 507636 320776 513380 320804
rect 507636 320764 507642 320776
rect 513374 320764 513380 320776
rect 513432 320764 513438 320816
rect 442626 320696 442632 320748
rect 442684 320736 442690 320748
rect 482094 320736 482100 320748
rect 442684 320708 482100 320736
rect 442684 320696 442690 320708
rect 482094 320696 482100 320708
rect 482152 320696 482158 320748
rect 507762 320696 507768 320748
rect 507820 320736 507826 320748
rect 510062 320736 510068 320748
rect 507820 320708 510068 320736
rect 507820 320696 507826 320708
rect 510062 320696 510068 320708
rect 510120 320696 510126 320748
rect 442534 320628 442540 320680
rect 442592 320668 442598 320680
rect 480714 320668 480720 320680
rect 442592 320640 480720 320668
rect 442592 320628 442598 320640
rect 480714 320628 480720 320640
rect 480772 320628 480778 320680
rect 457254 320084 457260 320136
rect 457312 320124 457318 320136
rect 459554 320124 459560 320136
rect 457312 320096 459560 320124
rect 457312 320084 457318 320096
rect 459554 320084 459560 320096
rect 459612 320084 459618 320136
rect 479058 320084 479064 320136
rect 479116 320124 479122 320136
rect 578878 320124 578884 320136
rect 479116 320096 578884 320124
rect 479116 320084 479122 320096
rect 578878 320084 578884 320096
rect 578936 320084 578942 320136
rect 456794 320016 456800 320068
rect 456852 320056 456858 320068
rect 472986 320056 472992 320068
rect 456852 320028 472992 320056
rect 456852 320016 456858 320028
rect 472986 320016 472992 320028
rect 473044 320016 473050 320068
rect 478782 320016 478788 320068
rect 478840 320056 478846 320068
rect 571978 320056 571984 320068
rect 478840 320028 571984 320056
rect 478840 320016 478846 320028
rect 571978 320016 571984 320028
rect 572036 320016 572042 320068
rect 446858 319948 446864 320000
rect 446916 319988 446922 320000
rect 462222 319988 462228 320000
rect 446916 319960 462228 319988
rect 446916 319948 446922 319960
rect 462222 319948 462228 319960
rect 462280 319948 462286 320000
rect 469122 319948 469128 320000
rect 469180 319988 469186 320000
rect 515398 319988 515404 320000
rect 469180 319960 515404 319988
rect 469180 319948 469186 319960
rect 515398 319948 515404 319960
rect 515456 319948 515462 320000
rect 450446 319880 450452 319932
rect 450504 319920 450510 319932
rect 461670 319920 461676 319932
rect 450504 319892 461676 319920
rect 450504 319880 450510 319892
rect 461670 319880 461676 319892
rect 461728 319880 461734 319932
rect 478506 319880 478512 319932
rect 478564 319920 478570 319932
rect 519538 319920 519544 319932
rect 478564 319892 519544 319920
rect 478564 319880 478570 319892
rect 519538 319880 519544 319892
rect 519596 319880 519602 319932
rect 444190 319812 444196 319864
rect 444248 319852 444254 319864
rect 458910 319852 458916 319864
rect 444248 319824 458916 319852
rect 444248 319812 444254 319824
rect 458910 319812 458916 319824
rect 458968 319812 458974 319864
rect 468846 319812 468852 319864
rect 468904 319852 468910 319864
rect 510522 319852 510528 319864
rect 468904 319824 510528 319852
rect 468904 319812 468910 319824
rect 510522 319812 510528 319824
rect 510580 319812 510586 319864
rect 449066 319744 449072 319796
rect 449124 319784 449130 319796
rect 472434 319784 472440 319796
rect 449124 319756 472440 319784
rect 449124 319744 449130 319756
rect 472434 319744 472440 319756
rect 472492 319744 472498 319796
rect 477402 319744 477408 319796
rect 477460 319784 477466 319796
rect 511902 319784 511908 319796
rect 477460 319756 511908 319784
rect 477460 319744 477466 319756
rect 511902 319744 511908 319756
rect 511960 319744 511966 319796
rect 446674 319676 446680 319728
rect 446732 319716 446738 319728
rect 469950 319716 469956 319728
rect 446732 319688 469956 319716
rect 446732 319676 446738 319688
rect 469950 319676 469956 319688
rect 470008 319676 470014 319728
rect 501414 319676 501420 319728
rect 501472 319716 501478 319728
rect 501472 319688 509234 319716
rect 501472 319676 501478 319688
rect 449526 319608 449532 319660
rect 449584 319648 449590 319660
rect 472710 319648 472716 319660
rect 449584 319620 472716 319648
rect 449584 319608 449590 319620
rect 472710 319608 472716 319620
rect 472768 319608 472774 319660
rect 445294 319540 445300 319592
rect 445352 319580 445358 319592
rect 480990 319580 480996 319592
rect 445352 319552 480996 319580
rect 445352 319540 445358 319552
rect 480990 319540 480996 319552
rect 481048 319540 481054 319592
rect 500310 319540 500316 319592
rect 500368 319580 500374 319592
rect 509206 319580 509234 319688
rect 534718 319580 534724 319592
rect 500368 319552 509096 319580
rect 509206 319552 534724 319580
rect 500368 319540 500374 319552
rect 445386 319472 445392 319524
rect 445444 319512 445450 319524
rect 482922 319512 482928 319524
rect 445444 319484 482928 319512
rect 445444 319472 445450 319484
rect 482922 319472 482928 319484
rect 482980 319472 482986 319524
rect 502518 319472 502524 319524
rect 502576 319472 502582 319524
rect 509068 319512 509096 319552
rect 534718 319540 534724 319552
rect 534776 319540 534782 319592
rect 538858 319512 538864 319524
rect 509068 319484 538864 319512
rect 538858 319472 538864 319484
rect 538916 319472 538922 319524
rect 445202 319404 445208 319456
rect 445260 319444 445266 319456
rect 470502 319444 470508 319456
rect 445260 319416 470508 319444
rect 445260 319404 445266 319416
rect 470502 319404 470508 319416
rect 470560 319404 470566 319456
rect 502536 319444 502564 319472
rect 543734 319444 543740 319456
rect 502536 319416 543740 319444
rect 543734 319404 543740 319416
rect 543792 319404 543798 319456
rect 449434 319336 449440 319388
rect 449492 319376 449498 319388
rect 482370 319376 482376 319388
rect 449492 319348 482376 319376
rect 449492 319336 449498 319348
rect 482370 319336 482376 319348
rect 482428 319336 482434 319388
rect 449342 319268 449348 319320
rect 449400 319308 449406 319320
rect 472158 319308 472164 319320
rect 449400 319280 472164 319308
rect 449400 319268 449406 319280
rect 472158 319268 472164 319280
rect 472216 319268 472222 319320
rect 449158 319200 449164 319252
rect 449216 319240 449222 319252
rect 469674 319240 469680 319252
rect 449216 319212 469680 319240
rect 449216 319200 449222 319212
rect 469674 319200 469680 319212
rect 469732 319200 469738 319252
rect 473446 319200 473452 319252
rect 473504 319240 473510 319252
rect 473722 319240 473728 319252
rect 473504 319212 473728 319240
rect 473504 319200 473510 319212
rect 473722 319200 473728 319212
rect 473780 319200 473786 319252
rect 496906 319200 496912 319252
rect 496964 319240 496970 319252
rect 497458 319240 497464 319252
rect 496964 319212 497464 319240
rect 496964 319200 496970 319212
rect 497458 319200 497464 319212
rect 497516 319200 497522 319252
rect 501046 319200 501052 319252
rect 501104 319240 501110 319252
rect 501598 319240 501604 319252
rect 501104 319212 501604 319240
rect 501104 319200 501110 319212
rect 501598 319200 501604 319212
rect 501656 319200 501662 319252
rect 454034 319132 454040 319184
rect 454092 319172 454098 319184
rect 455230 319172 455236 319184
rect 454092 319144 455236 319172
rect 454092 319132 454098 319144
rect 455230 319132 455236 319144
rect 455288 319132 455294 319184
rect 454218 319064 454224 319116
rect 454276 319104 454282 319116
rect 454678 319104 454684 319116
rect 454276 319076 454684 319104
rect 454276 319064 454282 319076
rect 454678 319064 454684 319076
rect 454736 319064 454742 319116
rect 455506 319064 455512 319116
rect 455564 319104 455570 319116
rect 456058 319104 456064 319116
rect 455564 319076 456064 319104
rect 455564 319064 455570 319076
rect 456058 319064 456064 319076
rect 456116 319064 456122 319116
rect 462682 319064 462688 319116
rect 462740 319104 462746 319116
rect 463510 319104 463516 319116
rect 462740 319076 463516 319104
rect 462740 319064 462746 319076
rect 463510 319064 463516 319076
rect 463568 319064 463574 319116
rect 463786 319064 463792 319116
rect 463844 319104 463850 319116
rect 464890 319104 464896 319116
rect 463844 319076 464896 319104
rect 463844 319064 463850 319076
rect 464890 319064 464896 319076
rect 464948 319064 464954 319116
rect 465442 319064 465448 319116
rect 465500 319104 465506 319116
rect 465994 319104 466000 319116
rect 465500 319076 466000 319104
rect 465500 319064 465506 319076
rect 465994 319064 466000 319076
rect 466052 319064 466058 319116
rect 475102 319064 475108 319116
rect 475160 319104 475166 319116
rect 475930 319104 475936 319116
rect 475160 319076 475936 319104
rect 475160 319064 475166 319076
rect 475930 319064 475936 319076
rect 475988 319064 475994 319116
rect 476206 319064 476212 319116
rect 476264 319104 476270 319116
rect 476758 319104 476764 319116
rect 476264 319076 476764 319104
rect 476264 319064 476270 319076
rect 476758 319064 476764 319076
rect 476816 319064 476822 319116
rect 483106 319064 483112 319116
rect 483164 319104 483170 319116
rect 483934 319104 483940 319116
rect 483164 319076 483940 319104
rect 483164 319064 483170 319076
rect 483934 319064 483940 319076
rect 483992 319064 483998 319116
rect 484486 319064 484492 319116
rect 484544 319104 484550 319116
rect 485590 319104 485596 319116
rect 484544 319076 485596 319104
rect 484544 319064 484550 319076
rect 485590 319064 485596 319076
rect 485648 319064 485654 319116
rect 495526 319064 495532 319116
rect 495584 319104 495590 319116
rect 496354 319104 496360 319116
rect 495584 319076 496360 319104
rect 495584 319064 495590 319076
rect 496354 319064 496360 319076
rect 496412 319064 496418 319116
rect 499666 319064 499672 319116
rect 499724 319104 499730 319116
rect 500770 319104 500776 319116
rect 499724 319076 500776 319104
rect 499724 319064 499730 319076
rect 500770 319064 500776 319076
rect 500828 319064 500834 319116
rect 504082 319064 504088 319116
rect 504140 319104 504146 319116
rect 504910 319104 504916 319116
rect 504140 319076 504916 319104
rect 504140 319064 504146 319076
rect 504910 319064 504916 319076
rect 504968 319064 504974 319116
rect 454126 318996 454132 319048
rect 454184 319036 454190 319048
rect 454954 319036 454960 319048
rect 454184 319008 454960 319036
rect 454184 318996 454190 319008
rect 454954 318996 454960 319008
rect 455012 318996 455018 319048
rect 462406 318996 462412 319048
rect 462464 319036 462470 319048
rect 463234 319036 463240 319048
rect 462464 319008 463240 319036
rect 462464 318996 462470 319008
rect 463234 318996 463240 319008
rect 463292 318996 463298 319048
rect 465166 318996 465172 319048
rect 465224 319036 465230 319048
rect 466270 319036 466276 319048
rect 465224 319008 466276 319036
rect 465224 318996 465230 319008
rect 466270 318996 466276 319008
rect 466328 318996 466334 319048
rect 474826 318996 474832 319048
rect 474884 319036 474890 319048
rect 475654 319036 475660 319048
rect 474884 319008 475660 319036
rect 474884 318996 474890 319008
rect 475654 318996 475660 319008
rect 475712 318996 475718 319048
rect 480898 318996 480904 319048
rect 480956 319036 480962 319048
rect 483750 319036 483756 319048
rect 480956 319008 483756 319036
rect 480956 318996 480962 319008
rect 483750 318996 483756 319008
rect 483808 318996 483814 319048
rect 498562 318928 498568 318980
rect 498620 318968 498626 318980
rect 499390 318968 499396 318980
rect 498620 318940 499396 318968
rect 498620 318928 498626 318940
rect 499390 318928 499396 318940
rect 499448 318928 499454 318980
rect 485038 318792 485044 318844
rect 485096 318832 485102 318844
rect 485314 318832 485320 318844
rect 485096 318804 485320 318832
rect 485096 318792 485102 318804
rect 485314 318792 485320 318804
rect 485372 318792 485378 318844
rect 444282 318724 444288 318776
rect 444340 318764 444346 318776
rect 469398 318764 469404 318776
rect 444340 318736 469404 318764
rect 444340 318724 444346 318736
rect 469398 318724 469404 318736
rect 469456 318724 469462 318776
rect 477126 318316 477132 318368
rect 477184 318356 477190 318368
rect 479518 318356 479524 318368
rect 477184 318328 479524 318356
rect 477184 318316 477190 318328
rect 479518 318316 479524 318328
rect 479576 318316 479582 318368
rect 432138 318112 432144 318164
rect 432196 318152 432202 318164
rect 439590 318152 439596 318164
rect 432196 318124 439596 318152
rect 432196 318112 432202 318124
rect 439590 318112 439596 318124
rect 439648 318112 439654 318164
rect 456426 318112 456432 318164
rect 456484 318152 456490 318164
rect 456484 318124 458680 318152
rect 456484 318112 456490 318124
rect 449618 318044 449624 318096
rect 449676 318084 449682 318096
rect 456886 318084 456892 318096
rect 449676 318056 456892 318084
rect 449676 318044 449682 318056
rect 456886 318044 456892 318056
rect 456944 318044 456950 318096
rect 458652 318084 458680 318124
rect 458818 318112 458824 318164
rect 458876 318152 458882 318164
rect 487338 318152 487344 318164
rect 458876 318124 487344 318152
rect 458876 318112 458882 318124
rect 487338 318112 487344 318124
rect 487396 318112 487402 318164
rect 494790 318112 494796 318164
rect 494848 318152 494854 318164
rect 540974 318152 540980 318164
rect 494848 318124 540980 318152
rect 494848 318112 494854 318124
rect 540974 318112 540980 318124
rect 541032 318112 541038 318164
rect 461578 318084 461584 318096
rect 458652 318056 461584 318084
rect 461578 318044 461584 318056
rect 461636 318044 461642 318096
rect 493962 318084 493968 318096
rect 470566 318056 493968 318084
rect 459094 317976 459100 318028
rect 459152 318016 459158 318028
rect 470566 318016 470594 318056
rect 493962 318044 493968 318056
rect 494020 318044 494026 318096
rect 495618 318044 495624 318096
rect 495676 318084 495682 318096
rect 543274 318084 543280 318096
rect 495676 318056 543280 318084
rect 495676 318044 495682 318056
rect 543274 318044 543280 318056
rect 543332 318044 543338 318096
rect 459152 317988 470594 318016
rect 459152 317976 459158 317988
rect 448422 317024 448428 317076
rect 448480 317064 448486 317076
rect 457806 317064 457812 317076
rect 448480 317036 457812 317064
rect 448480 317024 448486 317036
rect 457806 317024 457812 317036
rect 457864 317024 457870 317076
rect 447778 316956 447784 317008
rect 447836 316996 447842 317008
rect 462774 316996 462780 317008
rect 447836 316968 462780 316996
rect 447836 316956 447842 316968
rect 462774 316956 462780 316968
rect 462832 316956 462838 317008
rect 500034 316956 500040 317008
rect 500092 316996 500098 317008
rect 542630 316996 542636 317008
rect 500092 316968 542636 316996
rect 500092 316956 500098 316968
rect 542630 316956 542636 316968
rect 542688 316956 542694 317008
rect 457438 316888 457444 316940
rect 457496 316928 457502 316940
rect 490926 316928 490932 316940
rect 457496 316900 490932 316928
rect 457496 316888 457502 316900
rect 490926 316888 490932 316900
rect 490984 316888 490990 316940
rect 498378 316888 498384 316940
rect 498436 316928 498442 316940
rect 541066 316928 541072 316940
rect 498436 316900 541072 316928
rect 498436 316888 498442 316900
rect 541066 316888 541072 316900
rect 541124 316888 541130 316940
rect 453298 316820 453304 316872
rect 453356 316860 453362 316872
rect 489546 316860 489552 316872
rect 453356 316832 489552 316860
rect 453356 316820 453362 316832
rect 489546 316820 489552 316832
rect 489604 316820 489610 316872
rect 490006 316820 490012 316872
rect 490064 316860 490070 316872
rect 490282 316860 490288 316872
rect 490064 316832 490288 316860
rect 490064 316820 490070 316832
rect 490282 316820 490288 316832
rect 490340 316820 490346 316872
rect 493134 316820 493140 316872
rect 493192 316860 493198 316872
rect 493318 316860 493324 316872
rect 493192 316832 493324 316860
rect 493192 316820 493198 316832
rect 493318 316820 493324 316832
rect 493376 316820 493382 316872
rect 495894 316820 495900 316872
rect 495952 316860 495958 316872
rect 542446 316860 542452 316872
rect 495952 316832 542452 316860
rect 495952 316820 495958 316832
rect 542446 316820 542452 316832
rect 542504 316820 542510 316872
rect 454678 316752 454684 316804
rect 454736 316792 454742 316804
rect 502334 316792 502340 316804
rect 454736 316764 502340 316792
rect 454736 316752 454742 316764
rect 502334 316752 502340 316764
rect 502392 316752 502398 316804
rect 450538 316684 450544 316736
rect 450596 316724 450602 316736
rect 504726 316724 504732 316736
rect 450596 316696 504732 316724
rect 450596 316684 450602 316696
rect 504726 316684 504732 316696
rect 504784 316684 504790 316736
rect 486142 316616 486148 316668
rect 486200 316656 486206 316668
rect 486694 316656 486700 316668
rect 486200 316628 486700 316656
rect 486200 316616 486206 316628
rect 486694 316616 486700 316628
rect 486752 316616 486758 316668
rect 487798 316616 487804 316668
rect 487856 316656 487862 316668
rect 488350 316656 488356 316668
rect 487856 316628 488356 316656
rect 487856 316616 487862 316628
rect 488350 316616 488356 316628
rect 488408 316616 488414 316668
rect 488626 316616 488632 316668
rect 488684 316656 488690 316668
rect 489730 316656 489736 316668
rect 488684 316628 489736 316656
rect 488684 316616 488690 316628
rect 489730 316616 489736 316628
rect 489788 316616 489794 316668
rect 492766 316616 492772 316668
rect 492824 316656 492830 316668
rect 493594 316656 493600 316668
rect 492824 316628 493600 316656
rect 492824 316616 492830 316628
rect 493594 316616 493600 316628
rect 493652 316616 493658 316668
rect 494146 316616 494152 316668
rect 494204 316656 494210 316668
rect 495250 316656 495256 316668
rect 494204 316628 495256 316656
rect 494204 316616 494210 316628
rect 495250 316616 495256 316628
rect 495308 316616 495314 316668
rect 485866 316548 485872 316600
rect 485924 316588 485930 316600
rect 486418 316588 486424 316600
rect 485924 316560 486424 316588
rect 485924 316548 485930 316560
rect 486418 316548 486424 316560
rect 486476 316548 486482 316600
rect 490282 316548 490288 316600
rect 490340 316588 490346 316600
rect 491110 316588 491116 316600
rect 490340 316560 491116 316588
rect 490340 316548 490346 316560
rect 491110 316548 491116 316560
rect 491168 316548 491174 316600
rect 464246 316004 464252 316056
rect 464304 316044 464310 316056
rect 464430 316044 464436 316056
rect 464304 316016 464436 316044
rect 464304 316004 464310 316016
rect 464430 316004 464436 316016
rect 464488 316004 464494 316056
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 399478 315976 399484 315988
rect 361816 315948 399484 315976
rect 361816 315936 361822 315948
rect 399478 315936 399484 315948
rect 399536 315936 399542 315988
rect 499758 315460 499764 315512
rect 499816 315500 499822 315512
rect 539686 315500 539692 315512
rect 499816 315472 539692 315500
rect 499816 315460 499822 315472
rect 539686 315460 539692 315472
rect 539744 315460 539750 315512
rect 458910 315392 458916 315444
rect 458968 315432 458974 315444
rect 491386 315432 491392 315444
rect 458968 315404 491392 315432
rect 458968 315392 458974 315404
rect 491386 315392 491392 315404
rect 491444 315392 491450 315444
rect 496078 315392 496084 315444
rect 496136 315432 496142 315444
rect 539594 315432 539600 315444
rect 496136 315404 539600 315432
rect 496136 315392 496142 315404
rect 539594 315392 539600 315404
rect 539652 315392 539658 315444
rect 450722 315324 450728 315376
rect 450780 315364 450786 315376
rect 502978 315364 502984 315376
rect 450780 315336 502984 315364
rect 450780 315324 450786 315336
rect 502978 315324 502984 315336
rect 503036 315324 503042 315376
rect 450630 315256 450636 315308
rect 450688 315296 450694 315308
rect 504358 315296 504364 315308
rect 450688 315268 504364 315296
rect 450688 315256 450694 315268
rect 504358 315256 504364 315268
rect 504416 315256 504422 315308
rect 469858 314644 469864 314696
rect 469916 314684 469922 314696
rect 472342 314684 472348 314696
rect 469916 314656 472348 314684
rect 469916 314644 469922 314656
rect 472342 314644 472348 314656
rect 472400 314644 472406 314696
rect 501598 314032 501604 314084
rect 501656 314072 501662 314084
rect 538950 314072 538956 314084
rect 501656 314044 538956 314072
rect 501656 314032 501662 314044
rect 538950 314032 538956 314044
rect 539008 314032 539014 314084
rect 459002 313964 459008 314016
rect 459060 314004 459066 314016
rect 492306 314004 492312 314016
rect 459060 313976 492312 314004
rect 459060 313964 459066 313976
rect 492306 313964 492312 313976
rect 492364 313964 492370 314016
rect 495802 313964 495808 314016
rect 495860 314004 495866 314016
rect 542538 314004 542544 314016
rect 495860 313976 542544 314004
rect 495860 313964 495866 313976
rect 542538 313964 542544 313976
rect 542596 313964 542602 314016
rect 450814 313896 450820 313948
rect 450872 313936 450878 313948
rect 503898 313936 503904 313948
rect 450872 313908 503904 313936
rect 450872 313896 450878 313908
rect 503898 313896 503904 313908
rect 503956 313896 503962 313948
rect 466822 313216 466828 313268
rect 466880 313256 466886 313268
rect 580166 313256 580172 313268
rect 466880 313228 580172 313256
rect 466880 313216 466886 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 465258 312536 465264 312588
rect 465316 312576 465322 312588
rect 547138 312576 547144 312588
rect 465316 312548 547144 312576
rect 465316 312536 465322 312548
rect 547138 312536 547144 312548
rect 547196 312536 547202 312588
rect 487246 312128 487252 312180
rect 487304 312168 487310 312180
rect 488074 312168 488080 312180
rect 487304 312140 488080 312168
rect 487304 312128 487310 312140
rect 488074 312128 488080 312140
rect 488132 312128 488138 312180
rect 451918 311244 451924 311296
rect 451976 311284 451982 311296
rect 487890 311284 487896 311296
rect 451976 311256 487896 311284
rect 451976 311244 451982 311256
rect 487890 311244 487896 311256
rect 487948 311244 487954 311296
rect 501138 311244 501144 311296
rect 501196 311284 501202 311296
rect 540330 311284 540336 311296
rect 501196 311256 540336 311284
rect 501196 311244 501202 311256
rect 540330 311244 540336 311256
rect 540388 311244 540394 311296
rect 456058 311176 456064 311228
rect 456116 311216 456122 311228
rect 504174 311216 504180 311228
rect 456116 311188 504180 311216
rect 456116 311176 456122 311188
rect 504174 311176 504180 311188
rect 504232 311176 504238 311228
rect 455598 311108 455604 311160
rect 455656 311148 455662 311160
rect 533338 311148 533344 311160
rect 455656 311120 533344 311148
rect 455656 311108 455662 311120
rect 533338 311108 533344 311120
rect 533396 311108 533402 311160
rect 452010 309816 452016 309868
rect 452068 309856 452074 309868
rect 488810 309856 488816 309868
rect 452068 309828 488816 309856
rect 452068 309816 452074 309828
rect 488810 309816 488816 309828
rect 488868 309816 488874 309868
rect 475378 309748 475384 309800
rect 475436 309788 475442 309800
rect 565078 309788 565084 309800
rect 475436 309760 565084 309788
rect 475436 309748 475442 309760
rect 565078 309748 565084 309760
rect 565136 309748 565142 309800
rect 446398 308456 446404 308508
rect 446456 308496 446462 308508
rect 462958 308496 462964 308508
rect 446456 308468 462964 308496
rect 446456 308456 446462 308468
rect 462958 308456 462964 308468
rect 463016 308456 463022 308508
rect 453390 308388 453396 308440
rect 453448 308428 453454 308440
rect 489178 308428 489184 308440
rect 453448 308400 489184 308428
rect 453448 308388 453454 308400
rect 489178 308388 489184 308400
rect 489236 308388 489242 308440
rect 478138 307776 478144 307828
rect 478196 307816 478202 307828
rect 480898 307816 480904 307828
rect 478196 307788 480904 307816
rect 478196 307776 478202 307788
rect 480898 307776 480904 307788
rect 480956 307776 480962 307828
rect 432230 307708 432236 307760
rect 432288 307748 432294 307760
rect 436830 307748 436836 307760
rect 432288 307720 436836 307748
rect 432288 307708 432294 307720
rect 436830 307708 436836 307720
rect 436888 307708 436894 307760
rect 485958 307096 485964 307148
rect 486016 307136 486022 307148
rect 529934 307136 529940 307148
rect 486016 307108 529940 307136
rect 486016 307096 486022 307108
rect 529934 307096 529940 307108
rect 529992 307096 529998 307148
rect 475102 307028 475108 307080
rect 475160 307068 475166 307080
rect 569218 307068 569224 307080
rect 475160 307040 569224 307068
rect 475160 307028 475166 307040
rect 569218 307028 569224 307040
rect 569276 307028 569282 307080
rect 384298 306280 384304 306332
rect 384356 306320 384362 306332
rect 464062 306320 464068 306332
rect 384356 306292 464068 306320
rect 384356 306280 384362 306292
rect 464062 306280 464068 306292
rect 464120 306280 464126 306332
rect 386046 306212 386052 306264
rect 386104 306252 386110 306264
rect 474274 306252 474280 306264
rect 386104 306224 474280 306252
rect 386104 306212 386110 306224
rect 474274 306212 474280 306224
rect 474332 306212 474338 306264
rect 384482 306144 384488 306196
rect 384540 306184 384546 306196
rect 473998 306184 474004 306196
rect 384540 306156 474004 306184
rect 384540 306144 384546 306156
rect 473998 306144 474004 306156
rect 474056 306144 474062 306196
rect 384574 306076 384580 306128
rect 384632 306116 384638 306128
rect 474918 306116 474924 306128
rect 384632 306088 474924 306116
rect 384632 306076 384638 306088
rect 474918 306076 474924 306088
rect 474976 306076 474982 306128
rect 381722 306008 381728 306060
rect 381780 306048 381786 306060
rect 473722 306048 473728 306060
rect 381780 306020 473728 306048
rect 381780 306008 381786 306020
rect 473722 306008 473728 306020
rect 473780 306008 473786 306060
rect 384942 305940 384948 305992
rect 385000 305980 385006 305992
rect 484762 305980 484768 305992
rect 385000 305952 484768 305980
rect 385000 305940 385006 305952
rect 484762 305940 484768 305952
rect 484820 305940 484826 305992
rect 384666 305872 384672 305924
rect 384724 305912 384730 305924
rect 485130 305912 485136 305924
rect 384724 305884 485136 305912
rect 384724 305872 384730 305884
rect 485130 305872 485136 305884
rect 485188 305872 485194 305924
rect 381538 305804 381544 305856
rect 381596 305844 381602 305856
rect 484578 305844 484584 305856
rect 381596 305816 484584 305844
rect 381596 305804 381602 305816
rect 484578 305804 484584 305816
rect 484636 305804 484642 305856
rect 426342 305736 426348 305788
rect 426400 305776 426406 305788
rect 440234 305776 440240 305788
rect 426400 305748 440240 305776
rect 426400 305736 426406 305748
rect 440234 305736 440240 305748
rect 440292 305736 440298 305788
rect 455782 305736 455788 305788
rect 455840 305776 455846 305788
rect 574738 305776 574744 305788
rect 455840 305748 574744 305776
rect 455840 305736 455846 305748
rect 574738 305736 574744 305748
rect 574796 305736 574802 305788
rect 360838 305668 360844 305720
rect 360896 305708 360902 305720
rect 512270 305708 512276 305720
rect 360896 305680 512276 305708
rect 360896 305668 360902 305680
rect 512270 305668 512276 305680
rect 512328 305668 512334 305720
rect 360930 305600 360936 305652
rect 360988 305640 360994 305652
rect 512546 305640 512552 305652
rect 360988 305612 512552 305640
rect 360988 305600 360994 305612
rect 512546 305600 512552 305612
rect 512604 305600 512610 305652
rect 384390 305532 384396 305584
rect 384448 305572 384454 305584
rect 464430 305572 464436 305584
rect 384448 305544 464436 305572
rect 384448 305532 384454 305544
rect 464430 305532 464436 305544
rect 464488 305532 464494 305584
rect 385954 305464 385960 305516
rect 386012 305504 386018 305516
rect 464154 305504 464160 305516
rect 386012 305476 464160 305504
rect 386012 305464 386018 305476
rect 464154 305464 464160 305476
rect 464212 305464 464218 305516
rect 452194 305396 452200 305448
rect 452252 305436 452258 305448
rect 492950 305436 492956 305448
rect 452252 305408 492956 305436
rect 452252 305396 452258 305408
rect 492950 305396 492956 305408
rect 493008 305396 493014 305448
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 4798 305028 4804 305040
rect 3476 305000 4804 305028
rect 3476 304988 3482 305000
rect 4798 304988 4804 305000
rect 4856 304988 4862 305040
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 442350 304960 442356 304972
rect 361816 304932 442356 304960
rect 361816 304920 361822 304932
rect 442350 304920 442356 304932
rect 442408 304920 442414 304972
rect 486234 304444 486240 304496
rect 486292 304484 486298 304496
rect 530026 304484 530032 304496
rect 486292 304456 530032 304484
rect 486292 304444 486298 304456
rect 530026 304444 530032 304456
rect 530084 304444 530090 304496
rect 385862 304376 385868 304428
rect 385920 304416 385926 304428
rect 507026 304416 507032 304428
rect 385920 304388 507032 304416
rect 385920 304376 385926 304388
rect 507026 304376 507032 304388
rect 507084 304376 507090 304428
rect 362218 304308 362224 304360
rect 362276 304348 362282 304360
rect 512730 304348 512736 304360
rect 362276 304320 512736 304348
rect 362276 304308 362282 304320
rect 512730 304308 512736 304320
rect 512788 304308 512794 304360
rect 361022 304240 361028 304292
rect 361080 304280 361086 304292
rect 512178 304280 512184 304292
rect 361080 304252 512184 304280
rect 361080 304240 361086 304252
rect 512178 304240 512184 304252
rect 512236 304240 512242 304292
rect 463786 303560 463792 303612
rect 463844 303600 463850 303612
rect 562318 303600 562324 303612
rect 463844 303572 562324 303600
rect 463844 303560 463850 303572
rect 562318 303560 562324 303572
rect 562376 303560 562382 303612
rect 379330 303492 379336 303544
rect 379388 303532 379394 303544
rect 483658 303532 483664 303544
rect 379388 303504 483664 303532
rect 379388 303492 379394 303504
rect 483658 303492 483664 303504
rect 483716 303492 483722 303544
rect 486142 303492 486148 303544
rect 486200 303532 486206 303544
rect 528554 303532 528560 303544
rect 486200 303504 528560 303532
rect 486200 303492 486206 303504
rect 528554 303492 528560 303504
rect 528612 303492 528618 303544
rect 376478 303424 376484 303476
rect 376536 303464 376542 303476
rect 510890 303464 510896 303476
rect 376536 303436 510896 303464
rect 376536 303424 376542 303436
rect 510890 303424 510896 303436
rect 510948 303424 510954 303476
rect 376294 303356 376300 303408
rect 376352 303396 376358 303408
rect 510982 303396 510988 303408
rect 376352 303368 510988 303396
rect 376352 303356 376358 303368
rect 510982 303356 510988 303368
rect 511040 303356 511046 303408
rect 379146 303288 379152 303340
rect 379204 303328 379210 303340
rect 513926 303328 513932 303340
rect 379204 303300 513932 303328
rect 379204 303288 379210 303300
rect 513926 303288 513932 303300
rect 513984 303288 513990 303340
rect 379054 303220 379060 303272
rect 379112 303260 379118 303272
rect 514110 303260 514116 303272
rect 379112 303232 514116 303260
rect 379112 303220 379118 303232
rect 514110 303220 514116 303232
rect 514168 303220 514174 303272
rect 378962 303152 378968 303204
rect 379020 303192 379026 303204
rect 515306 303192 515312 303204
rect 379020 303164 515312 303192
rect 379020 303152 379026 303164
rect 515306 303152 515312 303164
rect 515364 303152 515370 303204
rect 376386 303084 376392 303136
rect 376444 303124 376450 303136
rect 515214 303124 515220 303136
rect 376444 303096 515220 303124
rect 376444 303084 376450 303096
rect 515214 303084 515220 303096
rect 515272 303084 515278 303136
rect 376202 303016 376208 303068
rect 376260 303056 376266 303068
rect 515122 303056 515128 303068
rect 376260 303028 515128 303056
rect 376260 303016 376266 303028
rect 515122 303016 515128 303028
rect 515180 303016 515186 303068
rect 373626 302948 373632 303000
rect 373684 302988 373690 303000
rect 513834 302988 513840 303000
rect 373684 302960 513840 302988
rect 373684 302948 373690 302960
rect 513834 302948 513840 302960
rect 513892 302948 513898 303000
rect 361114 302880 361120 302932
rect 361172 302920 361178 302932
rect 512362 302920 512368 302932
rect 361172 302892 512368 302920
rect 361172 302880 361178 302892
rect 512362 302880 512368 302892
rect 512420 302880 512426 302932
rect 379422 302812 379428 302864
rect 379480 302852 379486 302864
rect 473446 302852 473452 302864
rect 379480 302824 473452 302852
rect 379480 302812 379486 302824
rect 473446 302812 473452 302824
rect 473504 302812 473510 302864
rect 378686 302744 378692 302796
rect 378744 302784 378750 302796
rect 462406 302784 462412 302796
rect 378744 302756 462412 302784
rect 378744 302744 378750 302756
rect 462406 302744 462412 302756
rect 462464 302744 462470 302796
rect 382090 302676 382096 302728
rect 382148 302716 382154 302728
rect 462682 302716 462688 302728
rect 382148 302688 462688 302716
rect 382148 302676 382154 302688
rect 462682 302676 462688 302688
rect 462740 302676 462746 302728
rect 378778 302608 378784 302660
rect 378836 302648 378842 302660
rect 464338 302648 464344 302660
rect 378836 302620 464344 302648
rect 378836 302608 378842 302620
rect 464338 302608 464344 302620
rect 464396 302608 464402 302660
rect 3510 301928 3516 301980
rect 3568 301968 3574 301980
rect 4890 301968 4896 301980
rect 3568 301940 4896 301968
rect 3568 301928 3574 301940
rect 4890 301928 4896 301940
rect 4948 301928 4954 301980
rect 476298 301588 476304 301640
rect 476356 301628 476362 301640
rect 548518 301628 548524 301640
rect 476356 301600 548524 301628
rect 476356 301588 476362 301600
rect 548518 301588 548524 301600
rect 548576 301588 548582 301640
rect 407114 301520 407120 301572
rect 407172 301560 407178 301572
rect 502426 301560 502432 301572
rect 407172 301532 502432 301560
rect 407172 301520 407178 301532
rect 502426 301520 502432 301532
rect 502484 301520 502490 301572
rect 371878 301452 371884 301504
rect 371936 301492 371942 301504
rect 512454 301492 512460 301504
rect 371936 301464 512460 301492
rect 371936 301452 371942 301464
rect 512454 301452 512460 301464
rect 512512 301452 512518 301504
rect 373442 300772 373448 300824
rect 373500 300812 373506 300824
rect 509418 300812 509424 300824
rect 373500 300784 509424 300812
rect 373500 300772 373506 300784
rect 509418 300772 509424 300784
rect 509476 300772 509482 300824
rect 370682 300704 370688 300756
rect 370740 300744 370746 300756
rect 509326 300744 509332 300756
rect 370740 300716 509332 300744
rect 370740 300704 370746 300716
rect 509326 300704 509332 300716
rect 509384 300704 509390 300756
rect 370958 300636 370964 300688
rect 371016 300676 371022 300688
rect 510798 300676 510804 300688
rect 371016 300648 510804 300676
rect 371016 300636 371022 300648
rect 510798 300636 510804 300648
rect 510856 300636 510862 300688
rect 371050 300568 371056 300620
rect 371108 300608 371114 300620
rect 513558 300608 513564 300620
rect 371108 300580 513564 300608
rect 371108 300568 371114 300580
rect 513558 300568 513564 300580
rect 513616 300568 513622 300620
rect 370774 300500 370780 300552
rect 370832 300540 370838 300552
rect 513742 300540 513748 300552
rect 370832 300512 513748 300540
rect 370832 300500 370838 300512
rect 513742 300500 513748 300512
rect 513800 300500 513806 300552
rect 367738 300432 367744 300484
rect 367796 300472 367802 300484
rect 510706 300472 510712 300484
rect 367796 300444 510712 300472
rect 367796 300432 367802 300444
rect 510706 300432 510712 300444
rect 510764 300432 510770 300484
rect 370866 300364 370872 300416
rect 370924 300404 370930 300416
rect 515030 300404 515036 300416
rect 370924 300376 515036 300404
rect 370924 300364 370930 300376
rect 515030 300364 515036 300376
rect 515088 300364 515094 300416
rect 368014 300296 368020 300348
rect 368072 300336 368078 300348
rect 514938 300336 514944 300348
rect 368072 300308 514944 300336
rect 368072 300296 368078 300308
rect 514938 300296 514944 300308
rect 514996 300296 515002 300348
rect 365070 300228 365076 300280
rect 365128 300268 365134 300280
rect 513466 300268 513472 300280
rect 365128 300240 513472 300268
rect 365128 300228 365134 300240
rect 513466 300228 513472 300240
rect 513524 300228 513530 300280
rect 367922 300160 367928 300212
rect 367980 300200 367986 300212
rect 517698 300200 517704 300212
rect 367980 300172 517704 300200
rect 367980 300160 367986 300172
rect 517698 300160 517704 300172
rect 517756 300160 517762 300212
rect 367830 300092 367836 300144
rect 367888 300132 367894 300144
rect 517606 300132 517612 300144
rect 367888 300104 517612 300132
rect 367888 300092 367894 300104
rect 517606 300092 517612 300104
rect 517664 300092 517670 300144
rect 375926 300024 375932 300076
rect 375984 300064 375990 300076
rect 483106 300064 483112 300076
rect 375984 300036 483112 300064
rect 375984 300024 375990 300036
rect 483106 300024 483112 300036
rect 483164 300024 483170 300076
rect 465534 299956 465540 300008
rect 465592 299996 465598 300008
rect 566458 299996 566464 300008
rect 465592 299968 566464 299996
rect 465592 299956 465598 299968
rect 566458 299956 566464 299968
rect 566516 299956 566522 300008
rect 376662 299888 376668 299940
rect 376720 299928 376726 299940
rect 473538 299928 473544 299940
rect 376720 299900 473544 299928
rect 376720 299888 376726 299900
rect 473538 299888 473544 299900
rect 473596 299888 473602 299940
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 454770 297984 454776 298036
rect 454828 298024 454834 298036
rect 502702 298024 502708 298036
rect 454828 297996 502708 298024
rect 454828 297984 454834 297996
rect 502702 297984 502708 297996
rect 502760 297984 502766 298036
rect 454310 297916 454316 297968
rect 454368 297956 454374 297968
rect 563698 297956 563704 297968
rect 454368 297928 563704 297956
rect 454368 297916 454374 297928
rect 563698 297916 563704 297928
rect 563756 297916 563762 297968
rect 385678 297848 385684 297900
rect 385736 297888 385742 297900
rect 516594 297888 516600 297900
rect 385736 297860 516600 297888
rect 385736 297848 385742 297860
rect 516594 297848 516600 297860
rect 516652 297848 516658 297900
rect 384850 297780 384856 297832
rect 384908 297820 384914 297832
rect 516686 297820 516692 297832
rect 384908 297792 516692 297820
rect 384908 297780 384914 297792
rect 516686 297780 516692 297792
rect 516744 297780 516750 297832
rect 362494 297712 362500 297764
rect 362552 297752 362558 297764
rect 507762 297752 507768 297764
rect 362552 297724 507768 297752
rect 362552 297712 362558 297724
rect 507762 297712 507768 297724
rect 507820 297712 507826 297764
rect 364978 297644 364984 297696
rect 365036 297684 365042 297696
rect 511534 297684 511540 297696
rect 365036 297656 511540 297684
rect 365036 297644 365042 297656
rect 511534 297644 511540 297656
rect 511592 297644 511598 297696
rect 366542 297576 366548 297628
rect 366600 297616 366606 297628
rect 517974 297616 517980 297628
rect 366600 297588 517980 297616
rect 366600 297576 366606 297588
rect 517974 297576 517980 297588
rect 518032 297576 518038 297628
rect 365254 297508 365260 297560
rect 365312 297548 365318 297560
rect 517514 297548 517520 297560
rect 365312 297520 517520 297548
rect 365312 297508 365318 297520
rect 517514 297508 517520 297520
rect 517572 297508 517578 297560
rect 363690 297440 363696 297492
rect 363748 297480 363754 297492
rect 516962 297480 516968 297492
rect 363748 297452 516968 297480
rect 363748 297440 363754 297452
rect 516962 297440 516968 297452
rect 517020 297440 517026 297492
rect 363782 297372 363788 297424
rect 363840 297412 363846 297424
rect 518066 297412 518072 297424
rect 363840 297384 518072 297412
rect 363840 297372 363846 297384
rect 518066 297372 518072 297384
rect 518124 297372 518130 297424
rect 454218 295944 454224 295996
rect 454276 295984 454282 295996
rect 573358 295984 573364 295996
rect 454276 295956 573364 295984
rect 454276 295944 454282 295956
rect 573358 295944 573364 295956
rect 573416 295944 573422 295996
rect 374730 295264 374736 295316
rect 374788 295304 374794 295316
rect 514846 295304 514852 295316
rect 374788 295276 514852 295304
rect 374788 295264 374794 295276
rect 514846 295264 514852 295276
rect 514904 295264 514910 295316
rect 366726 295196 366732 295248
rect 366784 295236 366790 295248
rect 509510 295236 509516 295248
rect 366784 295208 509516 295236
rect 366784 295196 366790 295208
rect 509510 295196 509516 295208
rect 509568 295196 509574 295248
rect 370590 295128 370596 295180
rect 370648 295168 370654 295180
rect 513650 295168 513656 295180
rect 370648 295140 513656 295168
rect 370648 295128 370654 295140
rect 513650 295128 513656 295140
rect 513708 295128 513714 295180
rect 375006 295060 375012 295112
rect 375064 295100 375070 295112
rect 518986 295100 518992 295112
rect 375064 295072 518992 295100
rect 375064 295060 375070 295072
rect 518986 295060 518992 295072
rect 519044 295060 519050 295112
rect 373350 294992 373356 295044
rect 373408 295032 373414 295044
rect 519170 295032 519176 295044
rect 373408 295004 519176 295032
rect 373408 294992 373414 295004
rect 519170 294992 519176 295004
rect 519228 294992 519234 295044
rect 372246 294924 372252 294976
rect 372304 294964 372310 294976
rect 520366 294964 520372 294976
rect 372304 294936 520372 294964
rect 372304 294924 372310 294936
rect 520366 294924 520372 294936
rect 520424 294924 520430 294976
rect 368106 294856 368112 294908
rect 368164 294896 368170 294908
rect 516502 294896 516508 294908
rect 368164 294868 516508 294896
rect 368164 294856 368170 294868
rect 516502 294856 516508 294868
rect 516560 294856 516566 294908
rect 366450 294788 366456 294840
rect 366508 294828 366514 294840
rect 516318 294828 516324 294840
rect 366508 294800 516324 294828
rect 366508 294788 366514 294800
rect 516318 294788 516324 294800
rect 516376 294788 516382 294840
rect 369302 294720 369308 294772
rect 369360 294760 369366 294772
rect 519262 294760 519268 294772
rect 369360 294732 519268 294760
rect 369360 294720 369366 294732
rect 519262 294720 519268 294732
rect 519320 294720 519326 294772
rect 369210 294652 369216 294704
rect 369268 294692 369274 294704
rect 519446 294692 519452 294704
rect 369268 294664 519452 294692
rect 369268 294652 369274 294664
rect 519446 294652 519452 294664
rect 519504 294652 519510 294704
rect 365438 294584 365444 294636
rect 365496 294624 365502 294636
rect 517882 294624 517888 294636
rect 365496 294596 517888 294624
rect 365496 294584 365502 294596
rect 517882 294584 517888 294596
rect 517940 294584 517946 294636
rect 374822 294516 374828 294568
rect 374880 294556 374886 294568
rect 515582 294556 515588 294568
rect 374880 294528 515588 294556
rect 374880 294516 374886 294528
rect 515582 294516 515588 294528
rect 515640 294516 515646 294568
rect 454126 294448 454132 294500
rect 454184 294488 454190 294500
rect 578878 294488 578884 294500
rect 454184 294460 578884 294488
rect 454184 294448 454190 294460
rect 578878 294448 578884 294460
rect 578936 294448 578942 294500
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 385770 293944 385776 293956
rect 361816 293916 385776 293944
rect 361816 293904 361822 293916
rect 385770 293904 385776 293916
rect 385828 293904 385834 293956
rect 476482 293224 476488 293276
rect 476540 293264 476546 293276
rect 537478 293264 537484 293276
rect 476540 293236 537484 293264
rect 476540 293224 476546 293236
rect 537478 293224 537484 293236
rect 537536 293224 537542 293276
rect 383286 292476 383292 292528
rect 383344 292516 383350 292528
rect 507578 292516 507584 292528
rect 383344 292488 507584 292516
rect 383344 292476 383350 292488
rect 507578 292476 507584 292488
rect 507636 292476 507642 292528
rect 380526 292408 380532 292460
rect 380584 292448 380590 292460
rect 507670 292448 507676 292460
rect 380584 292420 507676 292448
rect 380584 292408 380590 292420
rect 507670 292408 507676 292420
rect 507728 292408 507734 292460
rect 378594 292340 378600 292392
rect 378652 292380 378658 292392
rect 507486 292380 507492 292392
rect 378652 292352 507492 292380
rect 378652 292340 378658 292352
rect 507486 292340 507492 292352
rect 507544 292340 507550 292392
rect 386322 292272 386328 292324
rect 386380 292312 386386 292324
rect 520734 292312 520740 292324
rect 386380 292284 520740 292312
rect 386380 292272 386386 292284
rect 520734 292272 520740 292284
rect 520792 292272 520798 292324
rect 377674 292204 377680 292256
rect 377732 292244 377738 292256
rect 514202 292244 514208 292256
rect 377732 292216 514208 292244
rect 377732 292204 377738 292216
rect 514202 292204 514208 292216
rect 514260 292204 514266 292256
rect 377582 292136 377588 292188
rect 377640 292176 377646 292188
rect 516134 292176 516140 292188
rect 377640 292148 516140 292176
rect 377640 292136 377646 292148
rect 516134 292136 516140 292148
rect 516192 292136 516198 292188
rect 381998 292068 382004 292120
rect 382056 292108 382062 292120
rect 520642 292108 520648 292120
rect 382056 292080 520648 292108
rect 382056 292068 382062 292080
rect 520642 292068 520648 292080
rect 520700 292068 520706 292120
rect 376570 292000 376576 292052
rect 376628 292040 376634 292052
rect 520274 292040 520280 292052
rect 376628 292012 520280 292040
rect 376628 292000 376634 292012
rect 520274 292000 520280 292012
rect 520332 292000 520338 292052
rect 375098 291932 375104 291984
rect 375156 291972 375162 291984
rect 518894 291972 518900 291984
rect 375156 291944 518900 291972
rect 375156 291932 375162 291944
rect 518894 291932 518900 291944
rect 518952 291932 518958 291984
rect 362310 291864 362316 291916
rect 362368 291904 362374 291916
rect 519722 291904 519728 291916
rect 362368 291876 519728 291904
rect 362368 291864 362374 291876
rect 519722 291864 519728 291876
rect 519780 291864 519786 291916
rect 361206 291796 361212 291848
rect 361264 291836 361270 291848
rect 520550 291836 520556 291848
rect 361264 291808 520556 291836
rect 361264 291796 361270 291808
rect 520550 291796 520556 291808
rect 520608 291796 520614 291848
rect 385770 291728 385776 291780
rect 385828 291768 385834 291780
rect 507394 291768 507400 291780
rect 385828 291740 507400 291768
rect 385828 291728 385834 291740
rect 507394 291728 507400 291740
rect 507452 291728 507458 291780
rect 362586 291660 362592 291712
rect 362644 291700 362650 291712
rect 443822 291700 443828 291712
rect 362644 291672 443828 291700
rect 362644 291660 362650 291672
rect 443822 291660 443828 291672
rect 443880 291660 443886 291712
rect 457530 291660 457536 291712
rect 457588 291700 457594 291712
rect 490190 291700 490196 291712
rect 457588 291672 490196 291700
rect 457588 291660 457594 291672
rect 490190 291660 490196 291672
rect 490248 291660 490254 291712
rect 499114 291660 499120 291712
rect 499172 291700 499178 291712
rect 541158 291700 541164 291712
rect 499172 291672 541164 291700
rect 499172 291660 499178 291672
rect 541158 291660 541164 291672
rect 541216 291660 541222 291712
rect 478230 291592 478236 291644
rect 478288 291632 478294 291644
rect 483382 291632 483388 291644
rect 478288 291604 483388 291632
rect 478288 291592 478294 291604
rect 483382 291592 483388 291604
rect 483440 291592 483446 291644
rect 465350 291184 465356 291236
rect 465408 291224 465414 291236
rect 469858 291224 469864 291236
rect 465408 291196 469864 291224
rect 465408 291184 465414 291196
rect 469858 291184 469864 291196
rect 469916 291184 469922 291236
rect 455506 290436 455512 290488
rect 455564 290476 455570 290488
rect 571978 290476 571984 290488
rect 455564 290448 571984 290476
rect 455564 290436 455570 290448
rect 571978 290436 571984 290448
rect 572036 290436 572042 290488
rect 380434 289756 380440 289808
rect 380492 289796 380498 289808
rect 519078 289796 519084 289808
rect 380492 289768 519084 289796
rect 380492 289756 380498 289768
rect 519078 289756 519084 289768
rect 519136 289756 519142 289808
rect 383194 289688 383200 289740
rect 383252 289728 383258 289740
rect 521930 289728 521936 289740
rect 383252 289700 521936 289728
rect 383252 289688 383258 289700
rect 521930 289688 521936 289700
rect 521988 289688 521994 289740
rect 363966 289620 363972 289672
rect 364024 289660 364030 289672
rect 507302 289660 507308 289672
rect 364024 289632 507308 289660
rect 364024 289620 364030 289632
rect 507302 289620 507308 289632
rect 507360 289620 507366 289672
rect 372062 289552 372068 289604
rect 372120 289592 372126 289604
rect 516226 289592 516232 289604
rect 372120 289564 516232 289592
rect 372120 289552 372126 289564
rect 516226 289552 516232 289564
rect 516284 289552 516290 289604
rect 366358 289484 366364 289536
rect 366416 289524 366422 289536
rect 510614 289524 510620 289536
rect 366416 289496 510620 289524
rect 366416 289484 366422 289496
rect 510614 289484 510620 289496
rect 510672 289484 510678 289536
rect 374914 289416 374920 289468
rect 374972 289456 374978 289468
rect 519354 289456 519360 289468
rect 374972 289428 519360 289456
rect 374972 289416 374978 289428
rect 519354 289416 519360 289428
rect 519412 289416 519418 289468
rect 377490 289348 377496 289400
rect 377548 289388 377554 289400
rect 522022 289388 522028 289400
rect 377548 289360 522028 289388
rect 377548 289348 377554 289360
rect 522022 289348 522028 289360
rect 522080 289348 522086 289400
rect 369394 289280 369400 289332
rect 369452 289320 369458 289332
rect 517790 289320 517796 289332
rect 369452 289292 517796 289320
rect 369452 289280 369458 289292
rect 517790 289280 517796 289292
rect 517848 289280 517854 289332
rect 366634 289212 366640 289264
rect 366692 289252 366698 289264
rect 516410 289252 516416 289264
rect 366692 289224 516416 289252
rect 366692 289212 366698 289224
rect 516410 289212 516416 289224
rect 516468 289212 516474 289264
rect 369118 289144 369124 289196
rect 369176 289184 369182 289196
rect 521746 289184 521752 289196
rect 369176 289156 521752 289184
rect 369176 289144 369182 289156
rect 521746 289144 521752 289156
rect 521804 289144 521810 289196
rect 363874 289076 363880 289128
rect 363932 289116 363938 289128
rect 519630 289116 519636 289128
rect 363932 289088 519636 289116
rect 363932 289076 363938 289088
rect 519630 289076 519636 289088
rect 519688 289076 519694 289128
rect 386230 289008 386236 289060
rect 386288 289048 386294 289060
rect 521838 289048 521844 289060
rect 386288 289020 521844 289048
rect 386288 289008 386294 289020
rect 521838 289008 521844 289020
rect 521896 289008 521902 289060
rect 441062 288940 441068 288992
rect 441120 288980 441126 288992
rect 446398 288980 446404 288992
rect 441120 288952 446404 288980
rect 441120 288940 441126 288952
rect 446398 288940 446404 288952
rect 446456 288940 446462 288992
rect 454126 288940 454132 288992
rect 454184 288980 454190 288992
rect 465350 288980 465356 288992
rect 454184 288952 465356 288980
rect 454184 288940 454190 288952
rect 465350 288940 465356 288952
rect 465408 288940 465414 288992
rect 474826 288940 474832 288992
rect 474884 288980 474890 288992
rect 544378 288980 544384 288992
rect 474884 288952 544384 288980
rect 474884 288940 474890 288952
rect 544378 288940 544384 288952
rect 544436 288940 544442 288992
rect 454034 287648 454040 287700
rect 454092 287688 454098 287700
rect 576118 287688 576124 287700
rect 454092 287660 576124 287688
rect 454092 287648 454098 287660
rect 576118 287648 576124 287660
rect 576176 287648 576182 287700
rect 485866 286832 485872 286884
rect 485924 286872 485930 286884
rect 530118 286872 530124 286884
rect 485924 286844 530124 286872
rect 485924 286832 485930 286844
rect 530118 286832 530124 286844
rect 530176 286832 530182 286884
rect 383102 286764 383108 286816
rect 383160 286804 383166 286816
rect 507118 286804 507124 286816
rect 383160 286776 507124 286804
rect 383160 286764 383166 286776
rect 507118 286764 507124 286776
rect 507176 286764 507182 286816
rect 377398 286696 377404 286748
rect 377456 286736 377462 286748
rect 507210 286736 507216 286748
rect 377456 286708 507216 286736
rect 377456 286696 377462 286708
rect 507210 286696 507216 286708
rect 507268 286696 507274 286748
rect 386138 286628 386144 286680
rect 386196 286668 386202 286680
rect 522390 286668 522396 286680
rect 386196 286640 522396 286668
rect 386196 286628 386202 286640
rect 522390 286628 522396 286640
rect 522448 286628 522454 286680
rect 381906 286560 381912 286612
rect 381964 286600 381970 286612
rect 522298 286600 522304 286612
rect 381964 286572 522304 286600
rect 381964 286560 381970 286572
rect 522298 286560 522304 286572
rect 522356 286560 522362 286612
rect 378870 286492 378876 286544
rect 378928 286532 378934 286544
rect 522206 286532 522212 286544
rect 378928 286504 522212 286532
rect 378928 286492 378934 286504
rect 522206 286492 522212 286504
rect 522264 286492 522270 286544
rect 376110 286424 376116 286476
rect 376168 286464 376174 286476
rect 520458 286464 520464 286476
rect 376168 286436 520464 286464
rect 376168 286424 376174 286436
rect 520458 286424 520464 286436
rect 520516 286424 520522 286476
rect 373258 286356 373264 286408
rect 373316 286396 373322 286408
rect 522114 286396 522120 286408
rect 373316 286368 522120 286396
rect 373316 286356 373322 286368
rect 522114 286356 522120 286368
rect 522172 286356 522178 286408
rect 372338 286288 372344 286340
rect 372396 286328 372402 286340
rect 521654 286328 521660 286340
rect 372396 286300 521660 286328
rect 372396 286288 372402 286300
rect 521654 286288 521660 286300
rect 521712 286288 521718 286340
rect 475378 285676 475384 285728
rect 475436 285716 475442 285728
rect 478138 285716 478144 285728
rect 475436 285688 478144 285716
rect 475436 285676 475442 285688
rect 478138 285676 478144 285688
rect 478196 285676 478202 285728
rect 453482 284996 453488 285048
rect 453540 285036 453546 285048
rect 487798 285036 487804 285048
rect 453540 285008 487804 285036
rect 453540 284996 453546 285008
rect 487798 284996 487804 285008
rect 487856 284996 487862 285048
rect 501322 284996 501328 285048
rect 501380 285036 501386 285048
rect 539042 285036 539048 285048
rect 501380 285008 539048 285036
rect 501380 284996 501386 285008
rect 539042 284996 539048 285008
rect 539100 284996 539106 285048
rect 476206 284928 476212 284980
rect 476264 284968 476270 284980
rect 570598 284968 570604 284980
rect 476264 284940 570604 284968
rect 476264 284928 476270 284940
rect 570598 284928 570604 284940
rect 570656 284928 570662 284980
rect 452102 283636 452108 283688
rect 452160 283676 452166 283688
rect 487246 283676 487252 283688
rect 452160 283648 487252 283676
rect 452160 283636 452166 283648
rect 487246 283636 487252 283648
rect 487304 283636 487310 283688
rect 496998 283636 497004 283688
rect 497056 283676 497062 283688
rect 539778 283676 539784 283688
rect 497056 283648 539784 283676
rect 497056 283636 497062 283648
rect 539778 283636 539784 283648
rect 539836 283636 539842 283688
rect 449158 283568 449164 283620
rect 449216 283608 449222 283620
rect 454126 283608 454132 283620
rect 449216 283580 454132 283608
rect 449216 283568 449222 283580
rect 454126 283568 454132 283580
rect 454184 283568 454190 283620
rect 465718 283568 465724 283620
rect 465776 283608 465782 283620
rect 554038 283608 554044 283620
rect 465776 283580 554044 283608
rect 465776 283568 465782 283580
rect 554038 283568 554044 283580
rect 554096 283568 554102 283620
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 435358 282860 435364 282872
rect 361816 282832 435364 282860
rect 361816 282820 361822 282832
rect 435358 282820 435364 282832
rect 435416 282820 435422 282872
rect 459278 282208 459284 282260
rect 459336 282248 459342 282260
rect 494238 282248 494244 282260
rect 459336 282220 494244 282248
rect 459336 282208 459342 282220
rect 494238 282208 494244 282220
rect 494296 282208 494302 282260
rect 465442 282140 465448 282192
rect 465500 282180 465506 282192
rect 555418 282180 555424 282192
rect 465500 282152 555424 282180
rect 465500 282140 465506 282152
rect 555418 282140 555424 282152
rect 555476 282140 555482 282192
rect 445018 281868 445024 281920
rect 445076 281908 445082 281920
rect 447778 281908 447784 281920
rect 445076 281880 447784 281908
rect 445076 281868 445082 281880
rect 447778 281868 447784 281880
rect 447836 281868 447842 281920
rect 452378 280848 452384 280900
rect 452436 280888 452442 280900
rect 493134 280888 493140 280900
rect 452436 280860 493140 280888
rect 452436 280848 452442 280860
rect 493134 280848 493140 280860
rect 493192 280848 493198 280900
rect 465166 280780 465172 280832
rect 465224 280820 465230 280832
rect 559558 280820 559564 280832
rect 465224 280792 559564 280820
rect 465224 280780 465230 280792
rect 559558 280780 559564 280792
rect 559616 280780 559622 280832
rect 454954 279420 454960 279472
rect 455012 279460 455018 279472
rect 487522 279460 487528 279472
rect 455012 279432 487528 279460
rect 455012 279420 455018 279432
rect 487522 279420 487528 279432
rect 487580 279420 487586 279472
rect 501046 279420 501052 279472
rect 501104 279460 501110 279472
rect 541526 279460 541532 279472
rect 501104 279432 541532 279460
rect 501104 279420 501110 279432
rect 541526 279420 541532 279432
rect 541584 279420 541590 279472
rect 453574 277992 453580 278044
rect 453632 278032 453638 278044
rect 492766 278032 492772 278044
rect 453632 278004 492772 278032
rect 453632 277992 453638 278004
rect 492766 277992 492772 278004
rect 492824 277992 492830 278044
rect 499942 277992 499948 278044
rect 500000 278032 500006 278044
rect 540238 278032 540244 278044
rect 500000 278004 540244 278032
rect 500000 277992 500006 278004
rect 540238 277992 540244 278004
rect 540296 277992 540302 278044
rect 456334 276768 456340 276820
rect 456392 276808 456398 276820
rect 492214 276808 492220 276820
rect 456392 276780 492220 276808
rect 456392 276768 456398 276780
rect 492214 276768 492220 276780
rect 492272 276768 492278 276820
rect 498838 276768 498844 276820
rect 498896 276808 498902 276820
rect 539962 276808 539968 276820
rect 498896 276780 539968 276808
rect 498896 276768 498902 276780
rect 539962 276768 539968 276780
rect 540020 276768 540026 276820
rect 449802 276700 449808 276752
rect 449860 276740 449866 276752
rect 536834 276740 536840 276752
rect 449860 276712 536840 276740
rect 449860 276700 449866 276712
rect 536834 276700 536840 276712
rect 536892 276700 536898 276752
rect 359458 276632 359464 276684
rect 359516 276672 359522 276684
rect 511994 276672 512000 276684
rect 359516 276644 512000 276672
rect 359516 276632 359522 276644
rect 511994 276632 512000 276644
rect 512052 276632 512058 276684
rect 465718 275476 465724 275528
rect 465776 275516 465782 275528
rect 478230 275516 478236 275528
rect 465776 275488 478236 275516
rect 465776 275476 465782 275488
rect 478230 275476 478236 275488
rect 478288 275476 478294 275528
rect 457622 275408 457628 275460
rect 457680 275448 457686 275460
rect 488626 275448 488632 275460
rect 457680 275420 488632 275448
rect 457680 275408 457686 275420
rect 488626 275408 488632 275420
rect 488684 275408 488690 275460
rect 457714 275340 457720 275392
rect 457772 275380 457778 275392
rect 491938 275380 491944 275392
rect 457772 275352 491944 275380
rect 457772 275340 457778 275352
rect 491938 275340 491944 275352
rect 491996 275340 492002 275392
rect 383378 275272 383384 275324
rect 383436 275312 383442 275324
rect 475194 275312 475200 275324
rect 383436 275284 475200 275312
rect 383436 275272 383442 275284
rect 475194 275272 475200 275284
rect 475252 275272 475258 275324
rect 497458 275272 497464 275324
rect 497516 275312 497522 275324
rect 541434 275312 541440 275324
rect 497516 275284 541440 275312
rect 497516 275272 497522 275284
rect 541434 275272 541440 275284
rect 541492 275272 541498 275324
rect 443822 274660 443828 274712
rect 443880 274700 443886 274712
rect 449158 274700 449164 274712
rect 443880 274672 449164 274700
rect 443880 274660 443886 274672
rect 449158 274660 449164 274672
rect 449216 274660 449222 274712
rect 460290 274048 460296 274100
rect 460348 274088 460354 274100
rect 494514 274088 494520 274100
rect 460348 274060 494520 274088
rect 460348 274048 460354 274060
rect 494514 274048 494520 274060
rect 494572 274048 494578 274100
rect 455046 273980 455052 274032
rect 455104 274020 455110 274032
rect 491662 274020 491668 274032
rect 455104 273992 491668 274020
rect 455104 273980 455110 273992
rect 491662 273980 491668 273992
rect 491720 273980 491726 274032
rect 368198 273912 368204 273964
rect 368256 273952 368262 273964
rect 485038 273952 485044 273964
rect 368256 273924 485044 273952
rect 368256 273912 368262 273924
rect 485038 273912 485044 273924
rect 485096 273912 485102 273964
rect 497182 273912 497188 273964
rect 497240 273952 497246 273964
rect 541250 273952 541256 273964
rect 497240 273924 541256 273952
rect 497240 273912 497246 273924
rect 541250 273912 541256 273924
rect 541308 273912 541314 273964
rect 479518 273164 479524 273216
rect 479576 273204 479582 273216
rect 580166 273204 580172 273216
rect 479576 273176 580172 273204
rect 479576 273164 479582 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 459186 272552 459192 272604
rect 459244 272592 459250 272604
rect 490558 272592 490564 272604
rect 459244 272564 490564 272592
rect 459244 272552 459250 272564
rect 490558 272552 490564 272564
rect 490616 272552 490622 272604
rect 433978 272484 433984 272536
rect 434036 272524 434042 272536
rect 445018 272524 445024 272536
rect 434036 272496 445024 272524
rect 434036 272484 434042 272496
rect 445018 272484 445024 272496
rect 445076 272484 445082 272536
rect 453666 272484 453672 272536
rect 453724 272524 453730 272536
rect 493042 272524 493048 272536
rect 453724 272496 493048 272524
rect 453724 272484 453730 272496
rect 493042 272484 493048 272496
rect 493100 272484 493106 272536
rect 498562 272484 498568 272536
rect 498620 272524 498626 272536
rect 540146 272524 540152 272536
rect 498620 272496 540152 272524
rect 498620 272484 498626 272496
rect 540146 272484 540152 272496
rect 540204 272484 540210 272536
rect 456242 271260 456248 271312
rect 456300 271300 456306 271312
rect 490282 271300 490288 271312
rect 456300 271272 490288 271300
rect 456300 271260 456306 271272
rect 490282 271260 490288 271272
rect 490340 271260 490346 271312
rect 456150 271192 456156 271244
rect 456208 271232 456214 271244
rect 490006 271232 490012 271244
rect 456208 271204 490012 271232
rect 456208 271192 456214 271204
rect 490006 271192 490012 271204
rect 490064 271192 490070 271244
rect 498286 271192 498292 271244
rect 498344 271232 498350 271244
rect 540054 271232 540060 271244
rect 498344 271204 540060 271232
rect 498344 271192 498350 271204
rect 540054 271192 540060 271204
rect 540112 271192 540118 271244
rect 452286 271124 452292 271176
rect 452344 271164 452350 271176
rect 488902 271164 488908 271176
rect 452344 271136 488908 271164
rect 452344 271124 452350 271136
rect 488902 271124 488908 271136
rect 488960 271124 488966 271176
rect 496906 271124 496912 271176
rect 496964 271164 496970 271176
rect 541342 271164 541348 271176
rect 496964 271136 541348 271164
rect 496964 271124 496970 271136
rect 541342 271124 541348 271136
rect 541400 271124 541406 271176
rect 455138 269900 455144 269952
rect 455196 269940 455202 269952
rect 486418 269940 486424 269952
rect 455196 269912 486424 269940
rect 455196 269900 455202 269912
rect 486418 269900 486424 269912
rect 486476 269900 486482 269952
rect 494146 269900 494152 269952
rect 494204 269940 494210 269952
rect 542722 269940 542728 269952
rect 494204 269912 542728 269940
rect 494204 269900 494210 269912
rect 542722 269900 542728 269912
rect 542780 269900 542786 269952
rect 466546 269832 466552 269884
rect 466604 269872 466610 269884
rect 580258 269872 580264 269884
rect 466604 269844 580264 269872
rect 466604 269832 466610 269844
rect 580258 269832 580264 269844
rect 580316 269832 580322 269884
rect 359550 269764 359556 269816
rect 359608 269804 359614 269816
rect 512086 269804 512092 269816
rect 359608 269776 512092 269804
rect 359608 269764 359614 269776
rect 512086 269764 512092 269776
rect 512144 269764 512150 269816
rect 459370 268540 459376 268592
rect 459428 268580 459434 268592
rect 465718 268580 465724 268592
rect 459428 268552 465724 268580
rect 459428 268540 459434 268552
rect 465718 268540 465724 268552
rect 465776 268540 465782 268592
rect 499666 268540 499672 268592
rect 499724 268580 499730 268592
rect 542906 268580 542912 268592
rect 499724 268552 542912 268580
rect 499724 268540 499730 268552
rect 542906 268540 542912 268552
rect 542964 268540 542970 268592
rect 445018 268472 445024 268524
rect 445076 268512 445082 268524
rect 475378 268512 475384 268524
rect 445076 268484 475384 268512
rect 445076 268472 445082 268484
rect 475378 268472 475384 268484
rect 475436 268472 475442 268524
rect 495526 268472 495532 268524
rect 495584 268512 495590 268524
rect 542814 268512 542820 268524
rect 495584 268484 542820 268512
rect 495584 268472 495590 268484
rect 542814 268472 542820 268484
rect 542872 268472 542878 268524
rect 457070 268404 457076 268456
rect 457128 268444 457134 268456
rect 505186 268444 505192 268456
rect 457128 268416 505192 268444
rect 457128 268404 457134 268416
rect 505186 268404 505192 268416
rect 505244 268404 505250 268456
rect 454862 268336 454868 268388
rect 454920 268376 454926 268388
rect 504082 268376 504088 268388
rect 454920 268348 504088 268376
rect 454920 268336 454926 268348
rect 504082 268336 504088 268348
rect 504140 268336 504146 268388
rect 424318 266976 424324 267028
rect 424376 267016 424382 267028
rect 433978 267016 433984 267028
rect 424376 266988 433984 267016
rect 424376 266976 424382 266988
rect 433978 266976 433984 266988
rect 434036 266976 434042 267028
rect 449710 263508 449716 263560
rect 449768 263548 449774 263560
rect 456794 263548 456800 263560
rect 449768 263520 456800 263548
rect 449768 263508 449774 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 440970 260828 440976 260840
rect 361816 260800 440976 260828
rect 361816 260788 361822 260800
rect 440970 260788 440976 260800
rect 441028 260788 441034 260840
rect 433978 260108 433984 260160
rect 434036 260148 434042 260160
rect 443822 260148 443828 260160
rect 434036 260120 443828 260148
rect 434036 260108 434042 260120
rect 443822 260108 443828 260120
rect 443880 260108 443886 260160
rect 3602 259360 3608 259412
rect 3660 259400 3666 259412
rect 4982 259400 4988 259412
rect 3660 259372 4988 259400
rect 3660 259360 3666 259372
rect 4982 259360 4988 259372
rect 5040 259360 5046 259412
rect 433702 255280 433708 255332
rect 433760 255320 433766 255332
rect 441062 255320 441068 255332
rect 433760 255292 441068 255320
rect 433760 255280 433766 255292
rect 441062 255280 441068 255292
rect 441120 255280 441126 255332
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 439498 249744 439504 249756
rect 361816 249716 439504 249744
rect 361816 249704 361822 249716
rect 439498 249704 439504 249716
rect 439556 249704 439562 249756
rect 446398 249024 446404 249076
rect 446456 249064 446462 249076
rect 456794 249064 456800 249076
rect 446456 249036 456800 249064
rect 446456 249024 446462 249036
rect 456794 249024 456800 249036
rect 456852 249024 456858 249076
rect 431310 248412 431316 248464
rect 431368 248452 431374 248464
rect 433702 248452 433708 248464
rect 431368 248424 433708 248452
rect 431368 248412 431374 248424
rect 433702 248412 433708 248424
rect 433760 248412 433766 248464
rect 571978 245556 571984 245608
rect 572036 245596 572042 245608
rect 580166 245596 580172 245608
rect 572036 245568 580172 245596
rect 572036 245556 572042 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3878 241408 3884 241460
rect 3936 241448 3942 241460
rect 5074 241448 5080 241460
rect 3936 241420 5080 241448
rect 3936 241408 3942 241420
rect 5074 241408 5080 241420
rect 5132 241408 5138 241460
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 442258 238728 442264 238740
rect 361816 238700 442264 238728
rect 361816 238688 361822 238700
rect 442258 238688 442264 238700
rect 442316 238688 442322 238740
rect 570598 233180 570604 233232
rect 570656 233220 570662 233232
rect 579982 233220 579988 233232
rect 570656 233192 579988 233220
rect 570656 233180 570662 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 421558 230460 421564 230512
rect 421616 230500 421622 230512
rect 424318 230500 424324 230512
rect 421616 230472 424324 230500
rect 421616 230460 421622 230472
rect 424318 230460 424324 230472
rect 424376 230460 424382 230512
rect 453850 227740 453856 227792
rect 453908 227780 453914 227792
rect 459370 227780 459376 227792
rect 453908 227752 459376 227780
rect 453908 227740 453914 227752
rect 459370 227740 459376 227752
rect 459428 227740 459434 227792
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 443730 227712 443736 227724
rect 361816 227684 443736 227712
rect 361816 227672 361822 227684
rect 443730 227672 443736 227684
rect 443788 227672 443794 227724
rect 432598 221416 432604 221468
rect 432656 221456 432662 221468
rect 453850 221456 453856 221468
rect 432656 221428 453856 221456
rect 432656 221416 432662 221428
rect 453850 221416 453856 221428
rect 453908 221416 453914 221468
rect 425698 220804 425704 220856
rect 425756 220844 425762 220856
rect 433978 220844 433984 220856
rect 425756 220816 433984 220844
rect 425756 220804 425762 220816
rect 433978 220804 433984 220816
rect 434036 220804 434042 220856
rect 414658 220056 414664 220108
rect 414716 220096 414722 220108
rect 447962 220096 447968 220108
rect 414716 220068 447968 220096
rect 414716 220056 414722 220068
rect 447962 220056 447968 220068
rect 448020 220096 448026 220108
rect 459462 220096 459468 220108
rect 448020 220068 459468 220096
rect 448020 220056 448026 220068
rect 459462 220056 459468 220068
rect 459520 220056 459526 220108
rect 559558 219376 559564 219428
rect 559616 219416 559622 219428
rect 580166 219416 580172 219428
rect 559616 219388 580172 219416
rect 559616 219376 559622 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3970 218016 3976 218068
rect 4028 218056 4034 218068
rect 5166 218056 5172 218068
rect 4028 218028 5172 218056
rect 4028 218016 4034 218028
rect 5166 218016 5172 218028
rect 5224 218016 5230 218068
rect 413278 218016 413284 218068
rect 413336 218056 413342 218068
rect 421558 218056 421564 218068
rect 413336 218028 421564 218056
rect 413336 218016 413342 218028
rect 421558 218016 421564 218028
rect 421616 218016 421622 218068
rect 361666 216316 361672 216368
rect 361724 216356 361730 216368
rect 364058 216356 364064 216368
rect 361724 216328 364064 216356
rect 361724 216316 361730 216328
rect 364058 216316 364064 216328
rect 364116 216316 364122 216368
rect 425790 213188 425796 213240
rect 425848 213228 425854 213240
rect 445018 213228 445024 213240
rect 425848 213200 445024 213228
rect 425848 213188 425854 213200
rect 445018 213188 445024 213200
rect 445076 213188 445082 213240
rect 424318 209040 424324 209092
rect 424376 209080 424382 209092
rect 432598 209080 432604 209092
rect 424376 209052 432604 209080
rect 424376 209040 424382 209052
rect 432598 209040 432604 209052
rect 432656 209040 432662 209092
rect 406286 207612 406292 207664
rect 406344 207652 406350 207664
rect 425790 207652 425796 207664
rect 406344 207624 425796 207652
rect 406344 207612 406350 207624
rect 425790 207612 425796 207624
rect 425848 207612 425854 207664
rect 574738 206932 574744 206984
rect 574796 206972 574802 206984
rect 579798 206972 579804 206984
rect 574796 206944 579804 206972
rect 574796 206932 574802 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 411254 206252 411260 206304
rect 411312 206292 411318 206304
rect 450906 206292 450912 206304
rect 411312 206264 450912 206292
rect 411312 206252 411318 206264
rect 450906 206252 450912 206264
rect 450964 206292 450970 206304
rect 456794 206292 456800 206304
rect 450964 206264 456800 206292
rect 450964 206252 450970 206264
rect 456794 206252 456800 206264
rect 456852 206252 456858 206304
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 440878 205612 440884 205624
rect 361816 205584 440884 205612
rect 361816 205572 361822 205584
rect 440878 205572 440884 205584
rect 440936 205572 440942 205624
rect 401594 200744 401600 200796
rect 401652 200784 401658 200796
rect 406286 200784 406292 200796
rect 401652 200756 406292 200784
rect 401652 200744 401658 200756
rect 406286 200744 406292 200756
rect 406344 200744 406350 200796
rect 421558 200744 421564 200796
rect 421616 200784 421622 200796
rect 431310 200784 431316 200796
rect 421616 200756 431316 200784
rect 421616 200744 421622 200756
rect 431310 200744 431316 200756
rect 431368 200744 431374 200796
rect 456794 200744 456800 200796
rect 456852 200784 456858 200796
rect 479518 200784 479524 200796
rect 456852 200756 479524 200784
rect 456852 200744 456858 200756
rect 479518 200744 479524 200756
rect 479576 200744 479582 200796
rect 459462 199384 459468 199436
rect 459520 199424 459526 199436
rect 485774 199424 485780 199436
rect 459520 199396 485780 199424
rect 459520 199384 459526 199396
rect 485774 199384 485780 199396
rect 485832 199384 485838 199436
rect 406378 195236 406384 195288
rect 406436 195276 406442 195288
rect 424318 195276 424324 195288
rect 406436 195248 424324 195276
rect 406436 195236 406442 195248
rect 424318 195236 424324 195248
rect 424376 195236 424382 195288
rect 422846 194692 422852 194744
rect 422904 194732 422910 194744
rect 425698 194732 425704 194744
rect 422904 194704 425704 194732
rect 422904 194692 422910 194704
rect 425698 194692 425704 194704
rect 425756 194692 425762 194744
rect 361758 194488 361764 194540
rect 361816 194528 361822 194540
rect 429838 194528 429844 194540
rect 361816 194500 429844 194528
rect 361816 194488 361822 194500
rect 429838 194488 429844 194500
rect 429896 194488 429902 194540
rect 388438 193808 388444 193860
rect 388496 193848 388502 193860
rect 401594 193848 401600 193860
rect 388496 193820 401600 193848
rect 388496 193808 388502 193820
rect 401594 193808 401600 193820
rect 401652 193808 401658 193860
rect 537478 193128 537484 193180
rect 537536 193168 537542 193180
rect 580166 193168 580172 193180
rect 537536 193140 580172 193168
rect 537536 193128 537542 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 411346 191088 411352 191140
rect 411404 191128 411410 191140
rect 422846 191128 422852 191140
rect 411404 191100 422852 191128
rect 411404 191088 411410 191100
rect 422846 191088 422852 191100
rect 422904 191088 422910 191140
rect 402238 188368 402244 188420
rect 402296 188408 402302 188420
rect 406378 188408 406384 188420
rect 402296 188380 406384 188408
rect 402296 188368 402302 188380
rect 406378 188368 406384 188380
rect 406436 188368 406442 188420
rect 398834 188300 398840 188352
rect 398892 188340 398898 188352
rect 411346 188340 411352 188352
rect 398892 188312 411352 188340
rect 398892 188300 398898 188312
rect 411346 188300 411352 188312
rect 411404 188300 411410 188352
rect 410518 186260 410524 186312
rect 410576 186300 410582 186312
rect 413278 186300 413284 186312
rect 410576 186272 413284 186300
rect 410576 186260 410582 186272
rect 413278 186260 413284 186272
rect 413336 186260 413342 186312
rect 366818 185580 366824 185632
rect 366876 185620 366882 185632
rect 388438 185620 388444 185632
rect 366876 185592 388444 185620
rect 366876 185580 366882 185592
rect 388438 185580 388444 185592
rect 388496 185580 388502 185632
rect 361758 183472 361764 183524
rect 361816 183512 361822 183524
rect 436738 183512 436744 183524
rect 361816 183484 436744 183512
rect 361816 183472 361822 183484
rect 436738 183472 436744 183484
rect 436796 183472 436802 183524
rect 391106 181432 391112 181484
rect 391164 181472 391170 181484
rect 398834 181472 398840 181484
rect 391164 181444 398840 181472
rect 391164 181432 391170 181444
rect 398834 181432 398840 181444
rect 398892 181432 398898 181484
rect 416038 179392 416044 179444
rect 416096 179432 416102 179444
rect 421558 179432 421564 179444
rect 416096 179404 421564 179432
rect 416096 179392 416102 179404
rect 421558 179392 421564 179404
rect 421616 179392 421622 179444
rect 555418 179324 555424 179376
rect 555476 179364 555482 179376
rect 580166 179364 580172 179376
rect 555476 179336 580172 179364
rect 555476 179324 555482 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 396718 178644 396724 178696
rect 396776 178684 396782 178696
rect 410518 178684 410524 178696
rect 396776 178656 410524 178684
rect 396776 178644 396782 178656
rect 410518 178644 410524 178656
rect 410576 178644 410582 178696
rect 398098 178032 398104 178084
rect 398156 178072 398162 178084
rect 402238 178072 402244 178084
rect 398156 178044 402244 178072
rect 398156 178032 398162 178044
rect 402238 178032 402244 178044
rect 402296 178032 402302 178084
rect 361298 175924 361304 175976
rect 361356 175964 361362 175976
rect 391106 175964 391112 175976
rect 361356 175936 391112 175964
rect 361356 175924 361362 175936
rect 391106 175924 391112 175936
rect 391164 175924 391170 175976
rect 364058 172524 364064 172576
rect 364116 172564 364122 172576
rect 366818 172564 366824 172576
rect 364116 172536 366824 172564
rect 364116 172524 364122 172536
rect 366818 172524 366824 172536
rect 366876 172524 366882 172576
rect 361758 171776 361764 171828
rect 361816 171816 361822 171828
rect 443638 171816 443644 171828
rect 361816 171788 443644 171816
rect 361816 171776 361822 171788
rect 443638 171776 443644 171788
rect 443696 171816 443702 171828
rect 524414 171816 524420 171828
rect 443696 171788 524420 171816
rect 443696 171776 443702 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 393958 167016 393964 167068
rect 394016 167056 394022 167068
rect 396718 167056 396724 167068
rect 394016 167028 396724 167056
rect 394016 167016 394022 167028
rect 396718 167016 396724 167028
rect 396776 167016 396782 167068
rect 533338 166948 533344 167000
rect 533396 166988 533402 167000
rect 580166 166988 580172 167000
rect 533396 166960 580172 166988
rect 533396 166948 533402 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 410242 164840 410248 164892
rect 410300 164880 410306 164892
rect 416038 164880 416044 164892
rect 410300 164852 416044 164880
rect 410300 164840 410306 164852
rect 416038 164840 416044 164852
rect 416096 164840 416102 164892
rect 447410 163548 447416 163600
rect 447468 163588 447474 163600
rect 461578 163588 461584 163600
rect 447468 163560 461584 163588
rect 447468 163548 447474 163560
rect 461578 163548 461584 163560
rect 461636 163548 461642 163600
rect 445662 163480 445668 163532
rect 445720 163520 445726 163532
rect 446398 163520 446404 163532
rect 445720 163492 446404 163520
rect 445720 163480 445726 163492
rect 446398 163480 446404 163492
rect 446456 163480 446462 163532
rect 447502 163480 447508 163532
rect 447560 163520 447566 163532
rect 528554 163520 528560 163532
rect 447560 163492 528560 163520
rect 447560 163480 447566 163492
rect 528554 163480 528560 163492
rect 528612 163480 528618 163532
rect 359642 163004 359648 163056
rect 359700 163044 359706 163056
rect 364058 163044 364064 163056
rect 359700 163016 364064 163044
rect 359700 163004 359706 163016
rect 364058 163004 364064 163016
rect 364116 163004 364122 163056
rect 407758 162256 407764 162308
rect 407816 162296 407822 162308
rect 410242 162296 410248 162308
rect 407816 162268 410248 162296
rect 407816 162256 407822 162268
rect 410242 162256 410248 162268
rect 410300 162256 410306 162308
rect 418706 162120 418712 162172
rect 418764 162160 418770 162172
rect 458082 162160 458088 162172
rect 418764 162132 458088 162160
rect 418764 162120 418770 162132
rect 458082 162120 458088 162132
rect 458140 162160 458146 162172
rect 489914 162160 489920 162172
rect 458140 162132 489920 162160
rect 458140 162120 458146 162132
rect 489914 162120 489920 162132
rect 489972 162120 489978 162172
rect 403618 161712 403624 161764
rect 403676 161752 403682 161764
rect 431218 161752 431224 161764
rect 403676 161724 431224 161752
rect 403676 161712 403682 161724
rect 431218 161712 431224 161724
rect 431276 161712 431282 161764
rect 426342 161644 426348 161696
rect 426400 161684 426406 161696
rect 496814 161684 496820 161696
rect 426400 161656 496820 161684
rect 426400 161644 426406 161656
rect 496814 161644 496820 161656
rect 496872 161644 496878 161696
rect 421558 161576 421564 161628
rect 421616 161616 421622 161628
rect 494054 161616 494060 161628
rect 421616 161588 494060 161616
rect 421616 161576 421622 161588
rect 494054 161576 494060 161588
rect 494112 161576 494118 161628
rect 407850 161508 407856 161560
rect 407908 161548 407914 161560
rect 438762 161548 438768 161560
rect 407908 161520 438768 161548
rect 407908 161508 407914 161520
rect 438762 161508 438768 161520
rect 438820 161548 438826 161560
rect 513374 161548 513380 161560
rect 438820 161520 513380 161548
rect 438820 161508 438826 161520
rect 513374 161508 513380 161520
rect 513432 161508 513438 161560
rect 362586 161440 362592 161492
rect 362644 161480 362650 161492
rect 441614 161480 441620 161492
rect 362644 161452 441620 161480
rect 362644 161440 362650 161452
rect 441614 161440 441620 161452
rect 441672 161480 441678 161492
rect 442902 161480 442908 161492
rect 441672 161452 442908 161480
rect 441672 161440 441678 161452
rect 442902 161440 442908 161452
rect 442960 161480 442966 161492
rect 517514 161480 517520 161492
rect 442960 161452 517520 161480
rect 442960 161440 442966 161452
rect 517514 161440 517520 161452
rect 517572 161440 517578 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 440142 161412 440148 161424
rect 361816 161384 440148 161412
rect 361816 161372 361822 161384
rect 440142 161372 440148 161384
rect 440200 161372 440206 161424
rect 440142 160692 440148 160744
rect 440200 160732 440206 160744
rect 521654 160732 521660 160744
rect 440200 160704 521660 160732
rect 440200 160692 440206 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 383470 160420 383476 160472
rect 383528 160460 383534 160472
rect 418154 160460 418160 160472
rect 383528 160432 418160 160460
rect 383528 160420 383534 160432
rect 418154 160420 418160 160432
rect 418212 160420 418218 160472
rect 410610 160352 410616 160404
rect 410668 160392 410674 160404
rect 410668 160364 431954 160392
rect 410668 160352 410674 160364
rect 385586 160284 385592 160336
rect 385644 160324 385650 160336
rect 414750 160324 414756 160336
rect 385644 160296 414756 160324
rect 385644 160284 385650 160296
rect 414750 160284 414756 160296
rect 414808 160284 414814 160336
rect 431926 160324 431954 160364
rect 435266 160324 435272 160336
rect 431926 160296 435272 160324
rect 435266 160284 435272 160296
rect 435324 160324 435330 160336
rect 436002 160324 436008 160336
rect 435324 160296 436008 160324
rect 435324 160284 435330 160296
rect 436002 160284 436008 160296
rect 436060 160324 436066 160336
rect 450906 160324 450912 160336
rect 436060 160296 450912 160324
rect 436060 160284 436066 160296
rect 450906 160284 450912 160296
rect 450964 160284 450970 160336
rect 410518 160216 410524 160268
rect 410576 160256 410582 160268
rect 427998 160256 428004 160268
rect 410576 160228 428004 160256
rect 410576 160216 410582 160228
rect 427998 160216 428004 160228
rect 428056 160216 428062 160268
rect 428642 160216 428648 160268
rect 428700 160256 428706 160268
rect 461670 160256 461676 160268
rect 428700 160228 461676 160256
rect 428700 160216 428706 160228
rect 461670 160216 461676 160228
rect 461728 160216 461734 160268
rect 395338 160148 395344 160200
rect 395396 160188 395402 160200
rect 398098 160188 398104 160200
rect 395396 160160 398104 160188
rect 395396 160148 395402 160160
rect 398098 160148 398104 160160
rect 398156 160148 398162 160200
rect 406378 160148 406384 160200
rect 406436 160188 406442 160200
rect 445202 160188 445208 160200
rect 406436 160160 445208 160188
rect 406436 160148 406442 160160
rect 445202 160148 445208 160160
rect 445260 160188 445266 160200
rect 445662 160188 445668 160200
rect 445260 160160 445668 160188
rect 445260 160148 445266 160160
rect 445662 160148 445668 160160
rect 445720 160188 445726 160200
rect 483658 160188 483664 160200
rect 445720 160160 483664 160188
rect 445720 160148 445726 160160
rect 483658 160148 483664 160160
rect 483716 160148 483722 160200
rect 381354 160080 381360 160132
rect 381412 160120 381418 160132
rect 425008 160120 425014 160132
rect 381412 160092 425014 160120
rect 381412 160080 381418 160092
rect 425008 160080 425014 160092
rect 425066 160120 425072 160132
rect 426342 160120 426348 160132
rect 425066 160092 426348 160120
rect 425066 160080 425072 160092
rect 426342 160080 426348 160092
rect 426400 160080 426406 160132
rect 431632 160080 431638 160132
rect 431690 160120 431696 160132
rect 504358 160120 504364 160132
rect 431690 160092 504364 160120
rect 431690 160080 431696 160092
rect 504358 160080 504364 160092
rect 504416 160080 504422 160132
rect 398098 159332 398104 159384
rect 398156 159372 398162 159384
rect 407758 159372 407764 159384
rect 398156 159344 407764 159372
rect 398156 159332 398162 159344
rect 407758 159332 407764 159344
rect 407816 159332 407822 159384
rect 421374 159372 421380 159384
rect 412606 159344 421380 159372
rect 364058 158720 364064 158772
rect 364116 158760 364122 158772
rect 412606 158760 412634 159344
rect 421374 159332 421380 159344
rect 421432 159332 421438 159384
rect 364116 158732 412634 158760
rect 364116 158720 364122 158732
rect 451550 158380 451556 158432
rect 451608 158420 451614 158432
rect 455138 158420 455144 158432
rect 451608 158392 455144 158420
rect 451608 158380 451614 158392
rect 455138 158380 455144 158392
rect 455196 158380 455202 158432
rect 365530 157972 365536 158024
rect 365588 158012 365594 158024
rect 393958 158012 393964 158024
rect 365588 157984 393964 158012
rect 365588 157972 365594 157984
rect 393958 157972 393964 157984
rect 394016 157972 394022 158024
rect 451734 157292 451740 157344
rect 451792 157332 451798 157344
rect 460290 157332 460296 157344
rect 451792 157304 460296 157332
rect 451792 157292 451798 157304
rect 460290 157292 460296 157304
rect 460348 157292 460354 157344
rect 452562 155524 452568 155576
rect 452620 155564 452626 155576
rect 459278 155564 459284 155576
rect 452620 155536 459284 155564
rect 452620 155524 452626 155536
rect 459278 155524 459284 155536
rect 459336 155524 459342 155576
rect 451734 154504 451740 154556
rect 451792 154544 451798 154556
rect 459094 154544 459100 154556
rect 451792 154516 459100 154544
rect 451792 154504 451798 154516
rect 459094 154504 459100 154516
rect 459152 154504 459158 154556
rect 451642 153144 451648 153196
rect 451700 153184 451706 153196
rect 453574 153184 453580 153196
rect 451700 153156 453580 153184
rect 451700 153144 451706 153156
rect 453574 153144 453580 153156
rect 453632 153144 453638 153196
rect 548518 153144 548524 153196
rect 548576 153184 548582 153196
rect 580166 153184 580172 153196
rect 548576 153156 580172 153184
rect 548576 153144 548582 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 451458 151444 451464 151496
rect 451516 151484 451522 151496
rect 453666 151484 453672 151496
rect 451516 151456 453672 151484
rect 451516 151444 451522 151456
rect 453666 151444 453672 151456
rect 453724 151444 453730 151496
rect 393958 150424 393964 150476
rect 394016 150464 394022 150476
rect 398098 150464 398104 150476
rect 394016 150436 398104 150464
rect 394016 150424 394022 150436
rect 398098 150424 398104 150436
rect 398156 150424 398162 150476
rect 390186 149336 390192 149388
rect 390244 149376 390250 149388
rect 395338 149376 395344 149388
rect 390244 149348 395344 149376
rect 390244 149336 390250 149348
rect 395338 149336 395344 149348
rect 395396 149336 395402 149388
rect 452562 147500 452568 147552
rect 452620 147540 452626 147552
rect 456334 147540 456340 147552
rect 452620 147512 456340 147540
rect 452620 147500 452626 147512
rect 456334 147500 456340 147512
rect 456392 147500 456398 147552
rect 452562 146004 452568 146056
rect 452620 146044 452626 146056
rect 459002 146044 459008 146056
rect 452620 146016 459008 146044
rect 452620 146004 452626 146016
rect 459002 146004 459008 146016
rect 459060 146004 459066 146056
rect 452562 144644 452568 144696
rect 452620 144684 452626 144696
rect 457714 144684 457720 144696
rect 452620 144656 457720 144684
rect 452620 144644 452626 144656
rect 457714 144644 457720 144656
rect 457772 144644 457778 144696
rect 504358 143488 504364 143540
rect 504416 143528 504422 143540
rect 505646 143528 505652 143540
rect 504416 143500 505652 143528
rect 504416 143488 504422 143500
rect 505646 143488 505652 143500
rect 505704 143488 505710 143540
rect 452562 143284 452568 143336
rect 452620 143324 452626 143336
rect 455046 143324 455052 143336
rect 452620 143296 455052 143324
rect 452620 143284 452626 143296
rect 455046 143284 455052 143296
rect 455104 143284 455110 143336
rect 387058 143080 387064 143132
rect 387116 143120 387122 143132
rect 390186 143120 390192 143132
rect 387116 143092 390192 143120
rect 387116 143080 387122 143092
rect 390186 143080 390192 143092
rect 390244 143080 390250 143132
rect 461670 142944 461676 142996
rect 461728 142984 461734 142996
rect 501690 142984 501696 142996
rect 461728 142956 501696 142984
rect 461728 142944 461734 142956
rect 501690 142944 501696 142956
rect 501748 142944 501754 142996
rect 483658 142876 483664 142928
rect 483716 142916 483722 142928
rect 533982 142916 533988 142928
rect 483716 142888 533988 142916
rect 483716 142876 483722 142888
rect 533982 142876 533988 142888
rect 534040 142876 534046 142928
rect 450906 142808 450912 142860
rect 450964 142848 450970 142860
rect 509602 142848 509608 142860
rect 450964 142820 509608 142848
rect 450964 142808 450970 142820
rect 509602 142808 509608 142820
rect 509660 142808 509666 142860
rect 362586 142128 362592 142180
rect 362644 142168 362650 142180
rect 365530 142168 365536 142180
rect 362644 142140 365536 142168
rect 362644 142128 362650 142140
rect 365530 142128 365536 142140
rect 365588 142128 365594 142180
rect 479518 142128 479524 142180
rect 479576 142168 479582 142180
rect 481910 142168 481916 142180
rect 479576 142140 481916 142168
rect 479576 142128 479582 142140
rect 481910 142128 481916 142140
rect 481968 142128 481974 142180
rect 533982 142128 533988 142180
rect 534040 142168 534046 142180
rect 539870 142168 539876 142180
rect 534040 142140 539876 142168
rect 534040 142128 534046 142140
rect 539870 142128 539876 142140
rect 539928 142128 539934 142180
rect 452562 141924 452568 141976
rect 452620 141964 452626 141976
rect 458910 141964 458916 141976
rect 452620 141936 458916 141964
rect 452620 141924 452626 141936
rect 458910 141924 458916 141936
rect 458968 141924 458974 141976
rect 462958 140768 462964 140820
rect 463016 140808 463022 140820
rect 481910 140808 481916 140820
rect 463016 140780 481916 140808
rect 463016 140768 463022 140780
rect 481910 140768 481916 140780
rect 481968 140768 481974 140820
rect 452562 140632 452568 140684
rect 452620 140672 452626 140684
rect 456242 140672 456248 140684
rect 452620 140644 456248 140672
rect 452620 140632 452626 140644
rect 456242 140632 456248 140644
rect 456300 140632 456306 140684
rect 534718 140020 534724 140072
rect 534776 140060 534782 140072
rect 543182 140060 543188 140072
rect 534776 140032 543188 140060
rect 534776 140020 534782 140032
rect 543182 140020 543188 140032
rect 543240 140020 543246 140072
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 407758 139380 407764 139392
rect 361816 139352 407764 139380
rect 361816 139340 361822 139352
rect 407758 139340 407764 139352
rect 407816 139340 407822 139392
rect 451550 139340 451556 139392
rect 451608 139380 451614 139392
rect 457438 139380 457444 139392
rect 451608 139352 457444 139380
rect 451608 139340 451614 139352
rect 457438 139340 457444 139352
rect 457496 139340 457502 139392
rect 554038 139340 554044 139392
rect 554096 139380 554102 139392
rect 580166 139380 580172 139392
rect 554096 139352 580172 139380
rect 554096 139340 554102 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 538858 138524 538864 138576
rect 538916 138564 538922 138576
rect 543090 138564 543096 138576
rect 538916 138536 543096 138564
rect 538916 138524 538922 138536
rect 543090 138524 543096 138536
rect 543148 138524 543154 138576
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 459186 137884 459192 137896
rect 452620 137856 459192 137884
rect 452620 137844 452626 137856
rect 459186 137844 459192 137856
rect 459244 137844 459250 137896
rect 452562 136484 452568 136536
rect 452620 136524 452626 136536
rect 456150 136524 456156 136536
rect 452620 136496 456156 136524
rect 452620 136484 452626 136496
rect 456150 136484 456156 136496
rect 456208 136484 456214 136536
rect 452562 135124 452568 135176
rect 452620 135164 452626 135176
rect 457530 135164 457536 135176
rect 452620 135136 457536 135164
rect 452620 135124 452626 135136
rect 457530 135124 457536 135136
rect 457588 135124 457594 135176
rect 452562 133764 452568 133816
rect 452620 133804 452626 133816
rect 457622 133804 457628 133816
rect 452620 133776 457628 133804
rect 452620 133764 452626 133776
rect 457622 133764 457628 133776
rect 457680 133764 457686 133816
rect 452194 132404 452200 132456
rect 452252 132444 452258 132456
rect 453298 132444 453304 132456
rect 452252 132416 453304 132444
rect 452252 132404 452258 132416
rect 453298 132404 453304 132416
rect 453356 132404 453362 132456
rect 359734 131112 359740 131164
rect 359792 131152 359798 131164
rect 362586 131152 362592 131164
rect 359792 131124 362592 131152
rect 359792 131112 359798 131124
rect 362586 131112 362592 131124
rect 362644 131112 362650 131164
rect 452378 131044 452384 131096
rect 452436 131084 452442 131096
rect 453390 131084 453396 131096
rect 452436 131056 453396 131084
rect 452436 131044 452442 131056
rect 453390 131044 453396 131056
rect 453448 131044 453454 131096
rect 390554 129752 390560 129804
rect 390612 129792 390618 129804
rect 393958 129792 393964 129804
rect 390612 129764 393964 129792
rect 390612 129752 390618 129764
rect 393958 129752 393964 129764
rect 394016 129752 394022 129804
rect 361758 128256 361764 128308
rect 361816 128296 361822 128308
rect 410610 128296 410616 128308
rect 361816 128268 410616 128296
rect 361816 128256 361822 128268
rect 410610 128256 410616 128268
rect 410668 128256 410674 128308
rect 361390 127576 361396 127628
rect 361448 127616 361454 127628
rect 390554 127616 390560 127628
rect 361448 127588 390560 127616
rect 361448 127576 361454 127588
rect 390554 127576 390560 127588
rect 390612 127576 390618 127628
rect 452378 126896 452384 126948
rect 452436 126936 452442 126948
rect 453482 126936 453488 126948
rect 452436 126908 453488 126936
rect 452436 126896 452442 126908
rect 453482 126896 453488 126908
rect 453540 126896 453546 126948
rect 576118 126896 576124 126948
rect 576176 126936 576182 126948
rect 580166 126936 580172 126948
rect 576176 126908 580172 126936
rect 576176 126896 576182 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 365530 126216 365536 126268
rect 365588 126256 365594 126268
rect 387058 126256 387064 126268
rect 365588 126228 387064 126256
rect 365588 126216 365594 126228
rect 387058 126216 387064 126228
rect 387116 126216 387122 126268
rect 451918 123360 451924 123412
rect 451976 123400 451982 123412
rect 454954 123400 454960 123412
rect 451976 123372 454960 123400
rect 451976 123360 451982 123372
rect 454954 123360 454960 123372
rect 455012 123360 455018 123412
rect 451918 122136 451924 122188
rect 451976 122176 451982 122188
rect 458818 122176 458824 122188
rect 451976 122148 458824 122176
rect 451976 122136 451982 122148
rect 458818 122136 458824 122148
rect 458876 122136 458882 122188
rect 359826 119076 359832 119128
rect 359884 119116 359890 119128
rect 365530 119116 365536 119128
rect 359884 119088 365536 119116
rect 359884 119076 359890 119088
rect 365530 119076 365536 119088
rect 365588 119076 365594 119128
rect 361758 117240 361764 117292
rect 361816 117280 361822 117292
rect 403618 117280 403624 117292
rect 361816 117252 403624 117280
rect 361816 117240 361822 117252
rect 403618 117240 403624 117252
rect 403676 117240 403682 117292
rect 569218 113092 569224 113144
rect 569276 113132 569282 113144
rect 579798 113132 579804 113144
rect 569276 113104 579804 113132
rect 569276 113092 569282 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 451182 107380 451188 107432
rect 451240 107420 451246 107432
rect 454862 107420 454868 107432
rect 451240 107392 454868 107420
rect 451240 107380 451246 107392
rect 454862 107380 454868 107392
rect 454920 107380 454926 107432
rect 439130 107244 439136 107296
rect 439188 107284 439194 107296
rect 450630 107284 450636 107296
rect 439188 107256 450636 107284
rect 439188 107244 439194 107256
rect 450630 107244 450636 107256
rect 450688 107244 450694 107296
rect 432966 107176 432972 107228
rect 433024 107216 433030 107228
rect 456058 107216 456064 107228
rect 433024 107188 456064 107216
rect 433024 107176 433030 107188
rect 456058 107176 456064 107188
rect 456116 107176 456122 107228
rect 426802 107108 426808 107160
rect 426860 107148 426866 107160
rect 450814 107148 450820 107160
rect 426860 107120 450820 107148
rect 426860 107108 426866 107120
rect 450814 107108 450820 107120
rect 450872 107108 450878 107160
rect 420638 107040 420644 107092
rect 420696 107080 420702 107092
rect 450722 107080 450728 107092
rect 420696 107052 450728 107080
rect 420696 107040 420702 107052
rect 450722 107040 450728 107052
rect 450780 107040 450786 107092
rect 389818 106972 389824 107024
rect 389876 107012 389882 107024
rect 406378 107012 406384 107024
rect 389876 106984 406384 107012
rect 389876 106972 389882 106984
rect 406378 106972 406384 106984
rect 406436 106972 406442 107024
rect 414474 106972 414480 107024
rect 414532 107012 414538 107024
rect 454770 107012 454776 107024
rect 414532 106984 454776 107012
rect 414532 106972 414538 106984
rect 454770 106972 454776 106984
rect 454828 106972 454834 107024
rect 402146 106904 402152 106956
rect 402204 106944 402210 106956
rect 454678 106944 454684 106956
rect 402204 106916 454684 106944
rect 402204 106904 402210 106916
rect 454678 106904 454684 106916
rect 454736 106904 454742 106956
rect 445294 106496 445300 106548
rect 445352 106536 445358 106548
rect 450538 106536 450544 106548
rect 445352 106508 450544 106536
rect 445352 106496 445358 106508
rect 450538 106496 450544 106508
rect 450596 106496 450602 106548
rect 361758 106224 361764 106276
rect 361816 106264 361822 106276
rect 410518 106264 410524 106276
rect 361816 106236 410524 106264
rect 361816 106224 361822 106236
rect 410518 106224 410524 106236
rect 410576 106224 410582 106276
rect 566458 100648 566464 100700
rect 566516 100688 566522 100700
rect 580166 100688 580172 100700
rect 566516 100660 580172 100688
rect 566516 100648 566522 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3694 98608 3700 98660
rect 3752 98648 3758 98660
rect 20898 98648 20904 98660
rect 3752 98620 20904 98648
rect 3752 98608 3758 98620
rect 20898 98608 20904 98620
rect 20956 98608 20962 98660
rect 361758 95140 361764 95192
rect 361816 95180 361822 95192
rect 381354 95180 381360 95192
rect 361816 95152 381360 95180
rect 361816 95140 361822 95152
rect 381354 95140 381360 95152
rect 381412 95140 381418 95192
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 20898 84232 20904 84244
rect 3200 84204 20904 84232
rect 3200 84192 3206 84204
rect 20898 84192 20904 84204
rect 20956 84192 20962 84244
rect 361666 84124 361672 84176
rect 361724 84164 361730 84176
rect 364058 84164 364064 84176
rect 361724 84136 364064 84164
rect 361724 84124 361730 84136
rect 364058 84124 364064 84136
rect 364116 84124 364122 84176
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 383470 73148 383476 73160
rect 361816 73120 383476 73148
rect 361816 73108 361822 73120
rect 383470 73108 383476 73120
rect 383528 73108 383534 73160
rect 544378 73108 544384 73160
rect 544436 73148 544442 73160
rect 580166 73148 580172 73160
rect 544436 73120 580172 73148
rect 544436 73108 544442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3142 70388 3148 70440
rect 3200 70428 3206 70440
rect 19978 70428 19984 70440
rect 3200 70400 19984 70428
rect 3200 70388 3206 70400
rect 19978 70388 19984 70400
rect 20036 70388 20042 70440
rect 4982 68960 4988 69012
rect 5040 69000 5046 69012
rect 8202 69000 8208 69012
rect 5040 68972 8208 69000
rect 5040 68960 5046 68972
rect 8202 68960 8208 68972
rect 8260 68960 8266 69012
rect 4890 66172 4896 66224
rect 4948 66212 4954 66224
rect 5534 66212 5540 66224
rect 4948 66184 5540 66212
rect 4948 66172 4954 66184
rect 5534 66172 5540 66184
rect 5592 66172 5598 66224
rect 5534 64132 5540 64184
rect 5592 64172 5598 64184
rect 10962 64172 10968 64184
rect 5592 64144 10968 64172
rect 5592 64132 5598 64144
rect 10962 64132 10968 64144
rect 11020 64132 11026 64184
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 385586 62064 385592 62076
rect 361816 62036 385592 62064
rect 361816 62024 361822 62036
rect 385586 62024 385592 62036
rect 385644 62024 385650 62076
rect 8294 60868 8300 60920
rect 8352 60908 8358 60920
rect 10318 60908 10324 60920
rect 8352 60880 10324 60908
rect 8352 60868 8358 60880
rect 10318 60868 10324 60880
rect 10376 60868 10382 60920
rect 5074 60664 5080 60716
rect 5132 60704 5138 60716
rect 9490 60704 9496 60716
rect 5132 60676 9496 60704
rect 5132 60664 5138 60676
rect 9490 60664 9496 60676
rect 9548 60664 9554 60716
rect 547138 60664 547144 60716
rect 547196 60704 547202 60716
rect 580166 60704 580172 60716
rect 547196 60676 580172 60704
rect 547196 60664 547202 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 11054 59372 11060 59424
rect 11112 59412 11118 59424
rect 11112 59384 12480 59412
rect 11112 59372 11118 59384
rect 12452 59344 12480 59384
rect 13814 59344 13820 59356
rect 12452 59316 13820 59344
rect 13814 59304 13820 59316
rect 13872 59304 13878 59356
rect 9490 59100 9496 59152
rect 9548 59140 9554 59152
rect 11054 59140 11060 59152
rect 9548 59112 11060 59140
rect 9548 59100 9554 59112
rect 11054 59100 11060 59112
rect 11112 59100 11118 59152
rect 3142 57944 3148 57996
rect 3200 57984 3206 57996
rect 20070 57984 20076 57996
rect 3200 57956 20076 57984
rect 3200 57944 3206 57956
rect 20070 57944 20076 57956
rect 20128 57944 20134 57996
rect 11054 57876 11060 57928
rect 11112 57916 11118 57928
rect 13722 57916 13728 57928
rect 11112 57888 13728 57916
rect 11112 57876 11118 57888
rect 13722 57876 13728 57888
rect 13780 57876 13786 57928
rect 4798 57128 4804 57180
rect 4856 57168 4862 57180
rect 7374 57168 7380 57180
rect 4856 57140 7380 57168
rect 4856 57128 4862 57140
rect 7374 57128 7380 57140
rect 7432 57128 7438 57180
rect 13814 56516 13820 56568
rect 13872 56556 13878 56568
rect 16482 56556 16488 56568
rect 13872 56528 16488 56556
rect 13872 56516 13878 56528
rect 16482 56516 16488 56528
rect 16540 56516 16546 56568
rect 7374 56108 7380 56160
rect 7432 56148 7438 56160
rect 10502 56148 10508 56160
rect 7432 56120 10508 56148
rect 7432 56108 7438 56120
rect 10502 56108 10508 56120
rect 10560 56108 10566 56160
rect 5166 54612 5172 54664
rect 5224 54652 5230 54664
rect 8202 54652 8208 54664
rect 5224 54624 8208 54652
rect 5224 54612 5230 54624
rect 8202 54612 8208 54624
rect 8260 54612 8266 54664
rect 13722 54340 13728 54392
rect 13780 54380 13786 54392
rect 15194 54380 15200 54392
rect 13780 54352 15200 54380
rect 13780 54340 13786 54352
rect 15194 54340 15200 54352
rect 15252 54340 15258 54392
rect 10502 53796 10508 53848
rect 10560 53836 10566 53848
rect 10560 53808 12480 53836
rect 10560 53796 10566 53808
rect 12452 53768 12480 53808
rect 17494 53768 17500 53780
rect 12452 53740 17500 53768
rect 17494 53728 17500 53740
rect 17552 53728 17558 53780
rect 16482 53456 16488 53508
rect 16540 53496 16546 53508
rect 18874 53496 18880 53508
rect 16540 53468 18880 53496
rect 16540 53456 16546 53468
rect 18874 53456 18880 53468
rect 18932 53456 18938 53508
rect 361758 51076 361764 51128
rect 361816 51116 361822 51128
rect 385586 51116 385592 51128
rect 361816 51088 385592 51116
rect 361816 51076 361822 51088
rect 385586 51076 385592 51088
rect 385644 51076 385650 51128
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 8202 51008 8208 51060
rect 8260 51048 8266 51060
rect 11698 51048 11704 51060
rect 8260 51020 11704 51048
rect 8260 51008 8266 51020
rect 11698 51008 11704 51020
rect 11756 51008 11762 51060
rect 10318 49716 10324 49768
rect 10376 49756 10382 49768
rect 10376 49728 11100 49756
rect 10376 49716 10382 49728
rect 11072 49688 11100 49728
rect 15286 49688 15292 49700
rect 11072 49660 15292 49688
rect 15286 49648 15292 49660
rect 15344 49648 15350 49700
rect 11698 48968 11704 49020
rect 11756 49008 11762 49020
rect 20622 49008 20628 49020
rect 11756 48980 20628 49008
rect 11756 48968 11762 48980
rect 20622 48968 20628 48980
rect 20680 48968 20686 49020
rect 17494 48288 17500 48340
rect 17552 48328 17558 48340
rect 17552 48300 19380 48328
rect 17552 48288 17558 48300
rect 19352 48260 19380 48300
rect 20714 48260 20720 48272
rect 19352 48232 20720 48260
rect 20714 48220 20720 48232
rect 20772 48220 20778 48272
rect 15286 46996 15292 47048
rect 15344 47036 15350 47048
rect 21266 47036 21272 47048
rect 15344 47008 21272 47036
rect 15344 46996 15350 47008
rect 21266 46996 21272 47008
rect 21324 46996 21330 47048
rect 3694 46860 3700 46912
rect 3752 46900 3758 46912
rect 386046 46900 386052 46912
rect 3752 46872 386052 46900
rect 3752 46860 3758 46872
rect 386046 46860 386052 46872
rect 386104 46860 386110 46912
rect 573358 46860 573364 46912
rect 573416 46900 573422 46912
rect 580166 46900 580172 46912
rect 573416 46872 580172 46900
rect 573416 46860 573422 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3234 46792 3240 46844
rect 3292 46832 3298 46844
rect 384482 46832 384488 46844
rect 3292 46804 384488 46832
rect 3292 46792 3298 46804
rect 384482 46792 384488 46804
rect 384540 46792 384546 46844
rect 3326 46724 3332 46776
rect 3384 46764 3390 46776
rect 384298 46764 384304 46776
rect 3384 46736 384304 46764
rect 3384 46724 3390 46736
rect 384298 46724 384304 46736
rect 384356 46724 384362 46776
rect 3970 46656 3976 46708
rect 4028 46696 4034 46708
rect 381722 46696 381728 46708
rect 4028 46668 381728 46696
rect 4028 46656 4034 46668
rect 381722 46656 381728 46668
rect 381780 46656 381786 46708
rect 4062 46588 4068 46640
rect 4120 46628 4126 46640
rect 381538 46628 381544 46640
rect 4120 46600 381544 46628
rect 4120 46588 4126 46600
rect 381538 46588 381544 46600
rect 381596 46588 381602 46640
rect 3602 46520 3608 46572
rect 3660 46560 3666 46572
rect 379422 46560 379428 46572
rect 3660 46532 379428 46560
rect 3660 46520 3666 46532
rect 379422 46520 379428 46532
rect 379480 46520 379486 46572
rect 3786 46452 3792 46504
rect 3844 46492 3850 46504
rect 379330 46492 379336 46504
rect 3844 46464 379336 46492
rect 3844 46452 3850 46464
rect 379330 46452 379336 46464
rect 379388 46452 379394 46504
rect 3510 46384 3516 46436
rect 3568 46424 3574 46436
rect 378686 46424 378692 46436
rect 3568 46396 378692 46424
rect 3568 46384 3574 46396
rect 378686 46384 378692 46396
rect 378744 46384 378750 46436
rect 3418 46316 3424 46368
rect 3476 46356 3482 46368
rect 375926 46356 375932 46368
rect 3476 46328 375932 46356
rect 3476 46316 3482 46328
rect 375926 46316 375932 46328
rect 375984 46316 375990 46368
rect 19978 46248 19984 46300
rect 20036 46288 20042 46300
rect 384390 46288 384396 46300
rect 20036 46260 384396 46288
rect 20036 46248 20042 46260
rect 384390 46248 384396 46260
rect 384448 46248 384454 46300
rect 21450 46180 21456 46232
rect 21508 46220 21514 46232
rect 384666 46220 384672 46232
rect 21508 46192 384672 46220
rect 21508 46180 21514 46192
rect 384666 46180 384672 46192
rect 384724 46180 384730 46232
rect 21266 46112 21272 46164
rect 21324 46152 21330 46164
rect 361390 46152 361396 46164
rect 21324 46124 361396 46152
rect 21324 46112 21330 46124
rect 361390 46112 361396 46124
rect 361448 46112 361454 46164
rect 20806 46044 20812 46096
rect 20864 46084 20870 46096
rect 359734 46084 359740 46096
rect 20864 46056 359740 46084
rect 20864 46044 20870 46056
rect 359734 46044 359740 46056
rect 359792 46044 359798 46096
rect 358262 45636 358268 45688
rect 358320 45676 358326 45688
rect 361298 45676 361304 45688
rect 358320 45648 361304 45676
rect 358320 45636 358326 45648
rect 361298 45636 361304 45648
rect 361356 45636 361362 45688
rect 3878 45500 3884 45552
rect 3936 45540 3942 45552
rect 382090 45540 382096 45552
rect 3936 45512 382096 45540
rect 3936 45500 3942 45512
rect 382090 45500 382096 45512
rect 382148 45500 382154 45552
rect 3418 45432 3424 45484
rect 3476 45472 3482 45484
rect 368198 45472 368204 45484
rect 3476 45444 368204 45472
rect 3476 45432 3482 45444
rect 368198 45432 368204 45444
rect 368256 45432 368262 45484
rect 21358 45364 21364 45416
rect 21416 45404 21422 45416
rect 376662 45404 376668 45416
rect 21416 45376 376668 45404
rect 21416 45364 21422 45376
rect 376662 45364 376668 45376
rect 376720 45364 376726 45416
rect 20714 45296 20720 45348
rect 20772 45336 20778 45348
rect 358262 45336 358268 45348
rect 20772 45308 358268 45336
rect 20772 45296 20778 45308
rect 358262 45296 358268 45308
rect 358320 45296 358326 45348
rect 69014 45228 69020 45280
rect 69072 45268 69078 45280
rect 376294 45268 376300 45280
rect 69072 45240 376300 45268
rect 69072 45228 69078 45240
rect 376294 45228 376300 45240
rect 376352 45228 376358 45280
rect 64874 45160 64880 45212
rect 64932 45200 64938 45212
rect 376386 45200 376392 45212
rect 64932 45172 376392 45200
rect 64932 45160 64938 45172
rect 376386 45160 376392 45172
rect 376444 45160 376450 45212
rect 60734 45092 60740 45144
rect 60792 45132 60798 45144
rect 379146 45132 379152 45144
rect 60792 45104 379152 45132
rect 60792 45092 60798 45104
rect 379146 45092 379152 45104
rect 379204 45092 379210 45144
rect 57974 45024 57980 45076
rect 58032 45064 58038 45076
rect 378962 45064 378968 45076
rect 58032 45036 378968 45064
rect 58032 45024 58038 45036
rect 378962 45024 378968 45036
rect 379020 45024 379026 45076
rect 53834 44956 53840 45008
rect 53892 44996 53898 45008
rect 379054 44996 379060 45008
rect 53892 44968 379060 44996
rect 53892 44956 53898 44968
rect 379054 44956 379060 44968
rect 379112 44956 379118 45008
rect 51074 44888 51080 44940
rect 51132 44928 51138 44940
rect 379238 44928 379244 44940
rect 51132 44900 379244 44928
rect 51132 44888 51138 44900
rect 379238 44888 379244 44900
rect 379296 44888 379302 44940
rect 46934 44820 46940 44872
rect 46992 44860 46998 44872
rect 381446 44860 381452 44872
rect 46992 44832 381452 44860
rect 46992 44820 46998 44832
rect 381446 44820 381452 44832
rect 381504 44820 381510 44872
rect 71774 44752 71780 44804
rect 71832 44792 71838 44804
rect 376202 44792 376208 44804
rect 71832 44764 376208 44792
rect 71832 44752 71838 44764
rect 376202 44752 376208 44764
rect 376260 44752 376266 44804
rect 75914 44684 75920 44736
rect 75972 44724 75978 44736
rect 376478 44724 376484 44736
rect 75972 44696 376484 44724
rect 75972 44684 75978 44696
rect 376478 44684 376484 44696
rect 376536 44684 376542 44736
rect 78674 44616 78680 44668
rect 78732 44656 78738 44668
rect 373626 44656 373632 44668
rect 78732 44628 373632 44656
rect 78732 44616 78738 44628
rect 373626 44616 373632 44628
rect 373684 44616 373690 44668
rect 114554 42712 114560 42764
rect 114612 42752 114618 42764
rect 367830 42752 367836 42764
rect 114612 42724 367836 42752
rect 114612 42712 114618 42724
rect 367830 42712 367836 42724
rect 367888 42712 367894 42764
rect 110414 42644 110420 42696
rect 110472 42684 110478 42696
rect 367922 42684 367928 42696
rect 110472 42656 367928 42684
rect 110472 42644 110478 42656
rect 367922 42644 367928 42656
rect 367980 42644 367986 42696
rect 107654 42576 107660 42628
rect 107712 42616 107718 42628
rect 368014 42616 368020 42628
rect 107712 42588 368020 42616
rect 107712 42576 107718 42588
rect 368014 42576 368020 42588
rect 368072 42576 368078 42628
rect 103514 42508 103520 42560
rect 103572 42548 103578 42560
rect 367738 42548 367744 42560
rect 103572 42520 367744 42548
rect 103572 42508 103578 42520
rect 367738 42508 367744 42520
rect 367796 42508 367802 42560
rect 100754 42440 100760 42492
rect 100812 42480 100818 42492
rect 370682 42480 370688 42492
rect 100812 42452 370688 42480
rect 100812 42440 100818 42452
rect 370682 42440 370688 42452
rect 370740 42440 370746 42492
rect 96614 42372 96620 42424
rect 96672 42412 96678 42424
rect 371050 42412 371056 42424
rect 96672 42384 371056 42412
rect 96672 42372 96678 42384
rect 371050 42372 371056 42384
rect 371108 42372 371114 42424
rect 93854 42304 93860 42356
rect 93912 42344 93918 42356
rect 370866 42344 370872 42356
rect 93912 42316 370872 42344
rect 93912 42304 93918 42316
rect 370866 42304 370872 42316
rect 370924 42304 370930 42356
rect 89714 42236 89720 42288
rect 89772 42276 89778 42288
rect 370774 42276 370780 42288
rect 89772 42248 370780 42276
rect 89772 42236 89778 42248
rect 370774 42236 370780 42248
rect 370832 42236 370838 42288
rect 85574 42168 85580 42220
rect 85632 42208 85638 42220
rect 370958 42208 370964 42220
rect 85632 42180 370964 42208
rect 85632 42168 85638 42180
rect 370958 42168 370964 42180
rect 371016 42168 371022 42220
rect 82814 42100 82820 42152
rect 82872 42140 82878 42152
rect 373442 42140 373448 42152
rect 82872 42112 373448 42140
rect 82872 42100 82878 42112
rect 373442 42100 373448 42112
rect 373500 42100 373506 42152
rect 11054 42032 11060 42084
rect 11112 42072 11118 42084
rect 373534 42072 373540 42084
rect 11112 42044 373540 42072
rect 11112 42032 11118 42044
rect 373534 42032 373540 42044
rect 373592 42032 373598 42084
rect 118694 41964 118700 42016
rect 118752 42004 118758 42016
rect 365070 42004 365076 42016
rect 118752 41976 365076 42004
rect 118752 41964 118758 41976
rect 365070 41964 365076 41976
rect 365128 41964 365134 42016
rect 461578 41352 461584 41404
rect 461636 41392 461642 41404
rect 536834 41392 536840 41404
rect 461636 41364 536840 41392
rect 461636 41352 461642 41364
rect 536834 41352 536840 41364
rect 536892 41352 536898 41404
rect 66254 39992 66260 40044
rect 66312 40032 66318 40044
rect 365438 40032 365444 40044
rect 66312 40004 365444 40032
rect 66312 39992 66318 40004
rect 365438 39992 365444 40004
rect 365496 39992 365502 40044
rect 62114 39924 62120 39976
rect 62172 39964 62178 39976
rect 366726 39964 366732 39976
rect 62172 39936 366732 39964
rect 62172 39924 62178 39936
rect 366726 39924 366732 39936
rect 366784 39924 366790 39976
rect 59354 39856 59360 39908
rect 59412 39896 59418 39908
rect 368106 39896 368112 39908
rect 59412 39868 368112 39896
rect 59412 39856 59418 39868
rect 368106 39856 368112 39868
rect 368164 39856 368170 39908
rect 55214 39788 55220 39840
rect 55272 39828 55278 39840
rect 366542 39828 366548 39840
rect 55272 39800 366548 39828
rect 55272 39788 55278 39800
rect 366542 39788 366548 39800
rect 366600 39788 366606 39840
rect 52454 39720 52460 39772
rect 52512 39760 52518 39772
rect 363782 39760 363788 39772
rect 52512 39732 363788 39760
rect 52512 39720 52518 39732
rect 363782 39720 363788 39732
rect 363840 39720 363846 39772
rect 33134 39652 33140 39704
rect 33192 39692 33198 39704
rect 363690 39692 363696 39704
rect 33192 39664 363696 39692
rect 33192 39652 33198 39664
rect 363690 39652 363696 39664
rect 363748 39652 363754 39704
rect 28994 39584 29000 39636
rect 29052 39624 29058 39636
rect 362402 39624 362408 39636
rect 29052 39596 362408 39624
rect 29052 39584 29058 39596
rect 362402 39584 362408 39596
rect 362460 39584 362466 39636
rect 26234 39516 26240 39568
rect 26292 39556 26298 39568
rect 362494 39556 362500 39568
rect 26292 39528 362500 39556
rect 26292 39516 26298 39528
rect 362494 39516 362500 39528
rect 362552 39516 362558 39568
rect 20714 39448 20720 39500
rect 20772 39488 20778 39500
rect 365162 39488 365168 39500
rect 20772 39460 365168 39488
rect 20772 39448 20778 39460
rect 365162 39448 365168 39460
rect 365220 39448 365226 39500
rect 40034 39380 40040 39432
rect 40092 39420 40098 39432
rect 384850 39420 384856 39432
rect 40092 39392 384856 39420
rect 40092 39380 40098 39392
rect 384850 39380 384856 39392
rect 384908 39380 384914 39432
rect 2774 39312 2780 39364
rect 2832 39352 2838 39364
rect 365346 39352 365352 39364
rect 2832 39324 365352 39352
rect 2832 39312 2838 39324
rect 365346 39312 365352 39324
rect 365404 39312 365410 39364
rect 121454 39244 121460 39296
rect 121512 39284 121518 39296
rect 365254 39284 365260 39296
rect 121512 39256 365260 39284
rect 121512 39244 121518 39256
rect 365254 39244 365260 39256
rect 365312 39244 365318 39296
rect 109034 37204 109040 37256
rect 109092 37244 109098 37256
rect 377674 37244 377680 37256
rect 109092 37216 377680 37244
rect 109092 37204 109098 37216
rect 377674 37204 377680 37216
rect 377732 37204 377738 37256
rect 104894 37136 104900 37188
rect 104952 37176 104958 37188
rect 375098 37176 375104 37188
rect 104952 37148 375104 37176
rect 104952 37136 104958 37148
rect 375098 37136 375104 37148
rect 375156 37136 375162 37188
rect 102134 37068 102140 37120
rect 102192 37108 102198 37120
rect 376570 37108 376576 37120
rect 102192 37080 376576 37108
rect 102192 37068 102198 37080
rect 376570 37068 376576 37080
rect 376628 37068 376634 37120
rect 97994 37000 98000 37052
rect 98052 37040 98058 37052
rect 374822 37040 374828 37052
rect 98052 37012 374828 37040
rect 98052 37000 98058 37012
rect 374822 37000 374828 37012
rect 374880 37000 374886 37052
rect 93946 36932 93952 36984
rect 94004 36972 94010 36984
rect 374730 36972 374736 36984
rect 94004 36944 374736 36972
rect 94004 36932 94010 36944
rect 374730 36932 374736 36944
rect 374788 36932 374794 36984
rect 91094 36864 91100 36916
rect 91152 36904 91158 36916
rect 375006 36904 375012 36916
rect 91152 36876 375012 36904
rect 91152 36864 91158 36876
rect 375006 36864 375012 36876
rect 375064 36864 375070 36916
rect 86954 36796 86960 36848
rect 87012 36836 87018 36848
rect 372246 36836 372252 36848
rect 87012 36808 372252 36836
rect 87012 36796 87018 36808
rect 372246 36796 372252 36808
rect 372304 36796 372310 36848
rect 84194 36728 84200 36780
rect 84252 36768 84258 36780
rect 373350 36768 373356 36780
rect 84252 36740 373356 36768
rect 84252 36728 84258 36740
rect 373350 36728 373356 36740
rect 373408 36728 373414 36780
rect 80054 36660 80060 36712
rect 80112 36700 80118 36712
rect 369302 36700 369308 36712
rect 80112 36672 369308 36700
rect 80112 36660 80118 36672
rect 369302 36660 369308 36672
rect 369360 36660 369366 36712
rect 73154 36592 73160 36644
rect 73212 36632 73218 36644
rect 369210 36632 369216 36644
rect 73212 36604 369216 36632
rect 73212 36592 73218 36604
rect 369210 36592 369216 36604
rect 369268 36592 369274 36644
rect 69106 36524 69112 36576
rect 69164 36564 69170 36576
rect 366450 36564 366456 36576
rect 69164 36536 366456 36564
rect 69164 36524 69170 36536
rect 366450 36524 366456 36536
rect 366508 36524 366514 36576
rect 111794 36456 111800 36508
rect 111852 36496 111858 36508
rect 378594 36496 378600 36508
rect 111852 36468 378600 36496
rect 111852 36456 111858 36468
rect 378594 36456 378600 36468
rect 378652 36456 378658 36508
rect 118786 34416 118792 34468
rect 118844 34456 118850 34468
rect 380250 34456 380256 34468
rect 118844 34428 380256 34456
rect 118844 34416 118850 34428
rect 380250 34416 380256 34428
rect 380308 34416 380314 34468
rect 115934 34348 115940 34400
rect 115992 34388 115998 34400
rect 377582 34388 377588 34400
rect 115992 34360 377588 34388
rect 115992 34348 115998 34360
rect 377582 34348 377588 34360
rect 377640 34348 377646 34400
rect 56594 34280 56600 34332
rect 56652 34320 56658 34332
rect 369394 34320 369400 34332
rect 56652 34292 369400 34320
rect 56652 34280 56658 34292
rect 369394 34280 369400 34292
rect 369452 34280 369458 34332
rect 49694 34212 49700 34264
rect 49752 34252 49758 34264
rect 366634 34252 366640 34264
rect 49752 34224 366640 34252
rect 49752 34212 49758 34224
rect 366634 34212 366640 34224
rect 366692 34212 366698 34264
rect 44174 34144 44180 34196
rect 44232 34184 44238 34196
rect 363874 34184 363880 34196
rect 44232 34156 363880 34184
rect 44232 34144 44238 34156
rect 363874 34144 363880 34156
rect 363932 34144 363938 34196
rect 41414 34076 41420 34128
rect 41472 34116 41478 34128
rect 361206 34116 361212 34128
rect 41472 34088 361212 34116
rect 41472 34076 41478 34088
rect 361206 34076 361212 34088
rect 361264 34076 361270 34128
rect 34514 34008 34520 34060
rect 34572 34048 34578 34060
rect 381998 34048 382004 34060
rect 34572 34020 382004 34048
rect 34572 34008 34578 34020
rect 381998 34008 382004 34020
rect 382056 34008 382062 34060
rect 9674 33940 9680 33992
rect 9732 33980 9738 33992
rect 363966 33980 363972 33992
rect 9732 33952 363972 33980
rect 9732 33940 9738 33952
rect 363966 33940 363972 33952
rect 364024 33940 364030 33992
rect 30374 33872 30380 33924
rect 30432 33912 30438 33924
rect 386322 33912 386328 33924
rect 30432 33884 386328 33912
rect 30432 33872 30438 33884
rect 386322 33872 386328 33884
rect 386380 33872 386386 33924
rect 22094 33804 22100 33856
rect 22152 33844 22158 33856
rect 383286 33844 383292 33856
rect 22152 33816 383292 33844
rect 22152 33804 22158 33816
rect 383286 33804 383292 33816
rect 383344 33804 383350 33856
rect 17954 33736 17960 33788
rect 18012 33776 18018 33788
rect 380526 33776 380532 33788
rect 18012 33748 380532 33776
rect 18012 33736 18018 33748
rect 380526 33736 380532 33748
rect 380584 33736 380590 33788
rect 122834 33668 122840 33720
rect 122892 33708 122898 33720
rect 382918 33708 382924 33720
rect 122892 33680 382924 33708
rect 122892 33668 122898 33680
rect 382918 33668 382924 33680
rect 382976 33668 382982 33720
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 378778 33096 378784 33108
rect 3568 33068 378784 33096
rect 3568 33056 3574 33068
rect 378778 33056 378784 33068
rect 378836 33056 378842 33108
rect 565078 33056 565084 33108
rect 565136 33096 565142 33108
rect 580166 33096 580172 33108
rect 565136 33068 580172 33096
rect 565136 33056 565142 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 113174 31696 113180 31748
rect 113232 31736 113238 31748
rect 372338 31736 372344 31748
rect 113232 31708 372344 31736
rect 113232 31696 113238 31708
rect 372338 31696 372344 31708
rect 372396 31696 372402 31748
rect 385586 31696 385592 31748
rect 385644 31736 385650 31748
rect 462314 31736 462320 31748
rect 385644 31708 462320 31736
rect 385644 31696 385650 31708
rect 462314 31696 462320 31708
rect 462372 31696 462378 31748
rect 106274 31628 106280 31680
rect 106332 31668 106338 31680
rect 369118 31668 369124 31680
rect 106332 31640 369124 31668
rect 106332 31628 106338 31640
rect 369118 31628 369124 31640
rect 369176 31628 369182 31680
rect 99374 31560 99380 31612
rect 99432 31600 99438 31612
rect 366358 31600 366364 31612
rect 99432 31572 366364 31600
rect 99432 31560 99438 31572
rect 366358 31560 366364 31572
rect 366416 31560 366422 31612
rect 88334 31492 88340 31544
rect 88392 31532 88398 31544
rect 385862 31532 385868 31544
rect 88392 31504 385868 31532
rect 88392 31492 88398 31504
rect 385862 31492 385868 31504
rect 385920 31492 385926 31544
rect 74534 31424 74540 31476
rect 74592 31464 74598 31476
rect 383194 31464 383200 31476
rect 74592 31436 383200 31464
rect 74592 31424 74598 31436
rect 383194 31424 383200 31436
rect 383252 31424 383258 31476
rect 77294 31356 77300 31408
rect 77352 31396 77358 31408
rect 386230 31396 386236 31408
rect 77352 31368 386236 31396
rect 77352 31356 77358 31368
rect 386230 31356 386236 31368
rect 386288 31356 386294 31408
rect 67634 31288 67640 31340
rect 67692 31328 67698 31340
rect 377490 31328 377496 31340
rect 67692 31300 377496 31328
rect 67692 31288 67698 31300
rect 377490 31288 377496 31300
rect 377548 31288 377554 31340
rect 70394 31220 70400 31272
rect 70452 31260 70458 31272
rect 380434 31260 380440 31272
rect 70452 31232 380440 31260
rect 70452 31220 70458 31232
rect 380434 31220 380440 31232
rect 380492 31220 380498 31272
rect 60826 31152 60832 31204
rect 60884 31192 60890 31204
rect 372062 31192 372068 31204
rect 60884 31164 372068 31192
rect 60884 31152 60890 31164
rect 372062 31152 372068 31164
rect 372120 31152 372126 31204
rect 63494 31084 63500 31136
rect 63552 31124 63558 31136
rect 374914 31124 374920 31136
rect 63552 31096 374920 31124
rect 63552 31084 63558 31096
rect 374914 31084 374920 31096
rect 374972 31084 374978 31136
rect 13814 31016 13820 31068
rect 13872 31056 13878 31068
rect 384758 31056 384764 31068
rect 13872 31028 384764 31056
rect 13872 31016 13878 31028
rect 384758 31016 384764 31028
rect 384816 31016 384822 31068
rect 124214 30948 124220 31000
rect 124272 30988 124278 31000
rect 380158 30988 380164 31000
rect 124272 30960 380164 30988
rect 124272 30948 124278 30960
rect 380158 30948 380164 30960
rect 380216 30948 380222 31000
rect 92474 29588 92480 29640
rect 92532 29628 92538 29640
rect 460198 29628 460204 29640
rect 92532 29600 460204 29628
rect 92532 29588 92538 29600
rect 460198 29588 460204 29600
rect 460256 29588 460262 29640
rect 117314 28636 117320 28688
rect 117372 28676 117378 28688
rect 374638 28676 374644 28688
rect 117372 28648 374644 28676
rect 117372 28636 117378 28648
rect 374638 28636 374644 28648
rect 374696 28636 374702 28688
rect 42794 28568 42800 28620
rect 42852 28608 42858 28620
rect 373258 28608 373264 28620
rect 42852 28580 373264 28608
rect 42852 28568 42858 28580
rect 373258 28568 373264 28580
rect 373316 28568 373322 28620
rect 38654 28500 38660 28552
rect 38712 28540 38718 28552
rect 376110 28540 376116 28552
rect 38712 28512 376116 28540
rect 38712 28500 38718 28512
rect 376110 28500 376116 28512
rect 376168 28500 376174 28552
rect 35894 28432 35900 28484
rect 35952 28472 35958 28484
rect 378870 28472 378876 28484
rect 35952 28444 378876 28472
rect 35952 28432 35958 28444
rect 378870 28432 378876 28444
rect 378928 28432 378934 28484
rect 31754 28364 31760 28416
rect 31812 28404 31818 28416
rect 381906 28404 381912 28416
rect 31812 28376 381912 28404
rect 31812 28364 31818 28376
rect 381906 28364 381912 28376
rect 381964 28364 381970 28416
rect 19334 28296 19340 28348
rect 19392 28336 19398 28348
rect 377398 28336 377404 28348
rect 19392 28308 377404 28336
rect 19392 28296 19398 28308
rect 377398 28296 377404 28308
rect 377456 28296 377462 28348
rect 27614 28228 27620 28280
rect 27672 28268 27678 28280
rect 386138 28268 386144 28280
rect 27672 28240 386144 28268
rect 27672 28228 27678 28240
rect 386138 28228 386144 28240
rect 386196 28228 386202 28280
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 383378 20652 383384 20664
rect 3476 20624 383384 20652
rect 3476 20612 3482 20624
rect 383378 20612 383384 20624
rect 383436 20612 383442 20664
rect 562318 20612 562324 20664
rect 562376 20652 562382 20664
rect 579982 20652 579988 20664
rect 562376 20624 579988 20652
rect 562376 20612 562382 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 376018 6848 376024 6860
rect 3476 6820 376024 6848
rect 3476 6808 3482 6820
rect 376018 6808 376024 6820
rect 376076 6808 376082 6860
rect 563698 6808 563704 6860
rect 563756 6848 563762 6860
rect 580166 6848 580172 6860
rect 563756 6820 580172 6848
rect 563756 6808 563762 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 360930 4128 360936 4140
rect 85724 4100 360936 4128
rect 85724 4088 85730 4100
rect 360930 4088 360936 4100
rect 360988 4088 360994 4140
rect 96246 4020 96252 4072
rect 96304 4060 96310 4072
rect 371878 4060 371884 4072
rect 96304 4032 371884 4060
rect 96304 4020 96310 4032
rect 371878 4020 371884 4032
rect 371936 4020 371942 4072
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 359458 3992 359464 4004
rect 82136 3964 359464 3992
rect 82136 3952 82142 3964
rect 359458 3952 359464 3964
rect 359516 3952 359522 4004
rect 77386 3884 77392 3936
rect 77444 3924 77450 3936
rect 370590 3924 370596 3936
rect 77444 3896 370596 3924
rect 77444 3884 77450 3896
rect 370590 3884 370596 3896
rect 370648 3884 370654 3936
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 359550 3856 359556 3868
rect 53800 3828 359556 3856
rect 53800 3816 53806 3828
rect 359550 3816 359556 3828
rect 359608 3816 359614 3868
rect 48958 3748 48964 3800
rect 49016 3788 49022 3800
rect 364978 3788 364984 3800
rect 49016 3760 364984 3788
rect 49016 3748 49022 3760
rect 364978 3748 364984 3760
rect 365036 3748 365042 3800
rect 46658 3680 46664 3732
rect 46716 3720 46722 3732
rect 363598 3720 363604 3732
rect 46716 3692 363604 3720
rect 46716 3680 46722 3692
rect 363598 3680 363604 3692
rect 363656 3680 363662 3732
rect 38378 3612 38384 3664
rect 38436 3652 38442 3664
rect 362310 3652 362316 3664
rect 38436 3624 362316 3652
rect 38436 3612 38442 3624
rect 362310 3612 362316 3624
rect 362368 3612 362374 3664
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 385770 3584 385776 3596
rect 27764 3556 385776 3584
rect 27764 3544 27770 3556
rect 385770 3544 385776 3556
rect 385828 3544 385834 3596
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 383102 3516 383108 3528
rect 24268 3488 383108 3516
rect 24268 3476 24274 3488
rect 383102 3476 383108 3488
rect 383160 3476 383166 3528
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 380342 3448 380348 3460
rect 17092 3420 380348 3448
rect 17092 3408 17098 3420
rect 380342 3408 380348 3420
rect 380400 3408 380406 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 103330 3340 103336 3392
rect 103388 3380 103394 3392
rect 361114 3380 361120 3392
rect 103388 3352 361120 3380
rect 103388 3340 103394 3352
rect 361114 3340 361120 3352
rect 361172 3340 361178 3392
rect 110414 3272 110420 3324
rect 110472 3312 110478 3324
rect 111610 3312 111616 3324
rect 110472 3284 111616 3312
rect 110472 3272 110478 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 360838 3312 360844 3324
rect 113146 3284 360844 3312
rect 110506 3204 110512 3256
rect 110564 3244 110570 3256
rect 113146 3244 113174 3284
rect 360838 3272 360844 3284
rect 360896 3272 360902 3324
rect 110564 3216 113174 3244
rect 110564 3204 110570 3216
rect 121086 3204 121092 3256
rect 121144 3244 121150 3256
rect 361022 3244 361028 3256
rect 121144 3216 361028 3244
rect 121144 3204 121150 3216
rect 361022 3204 361028 3216
rect 361080 3204 361086 3256
rect 44266 2184 44272 2236
rect 44324 2224 44330 2236
rect 385678 2224 385684 2236
rect 44324 2196 385684 2224
rect 44324 2184 44330 2196
rect 385678 2184 385684 2196
rect 385736 2184 385742 2236
rect 37182 2116 37188 2168
rect 37240 2156 37246 2168
rect 383010 2156 383016 2168
rect 37240 2128 383016 2156
rect 37240 2116 37246 2128
rect 383010 2116 383016 2128
rect 383068 2116 383074 2168
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 381630 2088 381636 2100
rect 2924 2060 381636 2088
rect 2924 2048 2930 2060
rect 381630 2048 381636 2060
rect 381688 2048 381694 2100
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 397460 700884 397512 700936
rect 446496 700884 446548 700936
rect 364984 700816 365036 700868
rect 445024 700816 445076 700868
rect 283840 700748 283892 700800
rect 446588 700748 446640 700800
rect 235172 700680 235224 700732
rect 445116 700680 445168 700732
rect 154120 700612 154172 700664
rect 416044 700612 416096 700664
rect 137836 700544 137888 700596
rect 450544 700544 450596 700596
rect 105452 700476 105504 700528
rect 444288 700476 444340 700528
rect 72976 700408 73028 700460
rect 444104 700408 444156 700460
rect 40500 700340 40552 700392
rect 450636 700340 450688 700392
rect 8116 700272 8168 700324
rect 418804 700272 418856 700324
rect 429844 700272 429896 700324
rect 446404 700272 446456 700324
rect 447784 700272 447836 700324
rect 478512 700272 478564 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 573364 696940 573416 696992
rect 580172 696940 580224 696992
rect 218060 686536 218112 686588
rect 445208 686536 445260 686588
rect 201500 686468 201552 686520
rect 445300 686468 445352 686520
rect 347780 685176 347832 685228
rect 446680 685176 446732 685228
rect 266360 685108 266412 685160
rect 418988 685108 419040 685160
rect 19984 684768 20036 684820
rect 418896 684768 418948 684820
rect 3608 684700 3660 684752
rect 420184 684700 420236 684752
rect 3332 684632 3384 684684
rect 420276 684632 420328 684684
rect 3148 684564 3200 684616
rect 420368 684564 420420 684616
rect 3884 684496 3936 684548
rect 445392 684496 445444 684548
rect 17960 683544 18012 683596
rect 359464 683544 359516 683596
rect 21364 683476 21416 683528
rect 420552 683476 420604 683528
rect 4068 683408 4120 683460
rect 420644 683408 420696 683460
rect 3516 683340 3568 683392
rect 420736 683340 420788 683392
rect 3700 683272 3752 683324
rect 445484 683272 445536 683324
rect 3424 683204 3476 683256
rect 445576 683204 445628 683256
rect 3976 683136 4028 683188
rect 446772 683136 446824 683188
rect 2964 682728 3016 682780
rect 420092 682728 420144 682780
rect 2872 682660 2924 682712
rect 450452 682660 450504 682712
rect 12900 680280 12952 680332
rect 17868 680348 17920 680400
rect 361764 678988 361816 679040
rect 364984 678988 365036 679040
rect 3516 678512 3568 678564
rect 3608 678512 3660 678564
rect 3516 678308 3568 678360
rect 3884 678172 3936 678224
rect 10416 676132 10468 676184
rect 12900 676200 12952 676252
rect 569224 670692 569276 670744
rect 580172 670692 580224 670744
rect 8024 667904 8076 667956
rect 10416 667904 10468 667956
rect 361764 667904 361816 667956
rect 381544 667904 381596 667956
rect 4804 665184 4856 665236
rect 8024 665184 8076 665236
rect 3148 658180 3200 658232
rect 19984 658180 20036 658232
rect 361672 656140 361724 656192
rect 406384 656140 406436 656192
rect 361764 645872 361816 645924
rect 378784 645872 378836 645924
rect 361580 634788 361632 634840
rect 407764 634788 407816 634840
rect 3700 631320 3752 631372
rect 20904 631320 20956 631372
rect 576124 630640 576176 630692
rect 579988 630640 580040 630692
rect 361580 623772 361632 623824
rect 376024 623772 376076 623824
rect 361580 612756 361632 612808
rect 410524 612756 410576 612808
rect 359464 601672 359516 601724
rect 361764 601672 361816 601724
rect 374736 601672 374788 601724
rect 366364 601604 366416 601656
rect 457536 600584 457588 600636
rect 461584 600584 461636 600636
rect 457352 599972 457404 600024
rect 462964 599972 463016 600024
rect 460204 599768 460256 599820
rect 463700 599768 463752 599820
rect 458824 599632 458876 599684
rect 466460 599632 466512 599684
rect 457904 599564 457956 599616
rect 469864 599564 469916 599616
rect 459928 598340 459980 598392
rect 463792 598340 463844 598392
rect 457720 598272 457772 598324
rect 464344 598272 464396 598324
rect 488632 598272 488684 598324
rect 494244 598272 494296 598324
rect 457628 598204 457680 598256
rect 468484 598204 468536 598256
rect 482284 598204 482336 598256
rect 494060 598204 494112 598256
rect 493324 597864 493376 597916
rect 494980 597864 495032 597916
rect 458732 596912 458784 596964
rect 465080 596912 465132 596964
rect 459836 596844 459888 596896
rect 466552 596844 466604 596896
rect 459744 596776 459796 596828
rect 470876 596776 470928 596828
rect 457444 596164 457496 596216
rect 461676 596164 461728 596216
rect 361764 590656 361816 590708
rect 371884 590656 371936 590708
rect 571984 590656 572036 590708
rect 579620 590656 579672 590708
rect 366364 590588 366416 590640
rect 367560 590588 367612 590640
rect 367560 586508 367612 586560
rect 372528 586440 372580 586492
rect 361764 579640 361816 579692
rect 370504 579640 370556 579692
rect 372620 577396 372672 577448
rect 374828 577396 374880 577448
rect 511264 576852 511316 576904
rect 579620 576852 579672 576904
rect 374828 571956 374880 572008
rect 376208 571956 376260 572008
rect 361764 568556 361816 568608
rect 367744 568556 367796 568608
rect 376208 568488 376260 568540
rect 377404 568488 377456 568540
rect 377404 564068 377456 564120
rect 380348 564068 380400 564120
rect 380348 559172 380400 559224
rect 384948 559172 385000 559224
rect 361580 557744 361632 557796
rect 363604 557744 363656 557796
rect 385040 551964 385092 552016
rect 387064 551964 387116 552016
rect 361580 546592 361632 546644
rect 363696 546592 363748 546644
rect 457812 542988 457864 543040
rect 468576 542988 468628 543040
rect 459560 541628 459612 541680
rect 470692 541628 470744 541680
rect 387064 540880 387116 540932
rect 388444 540880 388496 540932
rect 519544 536800 519596 536852
rect 580172 536800 580224 536852
rect 361580 535712 361632 535764
rect 363788 535712 363840 535764
rect 448060 526396 448112 526448
rect 500960 526396 501012 526448
rect 457260 525036 457312 525088
rect 465172 525036 465224 525088
rect 361764 524424 361816 524476
rect 411904 524424 411956 524476
rect 511356 524424 511408 524476
rect 580172 524424 580224 524476
rect 448428 523676 448480 523728
rect 506480 523676 506532 523728
rect 448336 522248 448388 522300
rect 493324 522248 493376 522300
rect 474740 521636 474792 521688
rect 475200 521636 475252 521688
rect 494336 521636 494388 521688
rect 458088 520956 458140 521008
rect 465724 520956 465776 521008
rect 449716 520888 449768 520940
rect 475200 520888 475252 520940
rect 482652 520888 482704 520940
rect 520280 520888 520332 520940
rect 461768 520412 461820 520464
rect 488632 520412 488684 520464
rect 467840 520344 467892 520396
rect 469128 520344 469180 520396
rect 494244 520344 494296 520396
rect 477408 520276 477460 520328
rect 482652 520276 482704 520328
rect 457996 519596 458048 519648
rect 468760 519596 468812 519648
rect 447968 519528 448020 519580
rect 467840 519528 467892 519580
rect 449808 518168 449860 518220
rect 462412 518168 462464 518220
rect 388444 517488 388496 517540
rect 389456 517488 389508 517540
rect 459652 517488 459704 517540
rect 462504 517488 462556 517540
rect 491852 516128 491904 516180
rect 448428 516060 448480 516112
rect 494060 515380 494112 515432
rect 538220 515380 538272 515432
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 361764 513340 361816 513392
rect 414664 513340 414716 513392
rect 494060 512592 494112 512644
rect 494428 512592 494480 512644
rect 535460 512592 535512 512644
rect 389456 511980 389508 512032
rect 393228 511912 393280 511964
rect 567844 510620 567896 510672
rect 580172 510620 580224 510672
rect 494336 508512 494388 508564
rect 532700 508512 532752 508564
rect 393320 506744 393372 506796
rect 396724 506744 396776 506796
rect 495072 505724 495124 505776
rect 529940 505724 529992 505776
rect 361764 502324 361816 502376
rect 416136 502324 416188 502376
rect 448520 500216 448572 500268
rect 545120 500216 545172 500268
rect 448520 498788 448572 498840
rect 542452 498788 542504 498840
rect 453304 497428 453356 497480
rect 480260 497428 480312 497480
rect 454040 497020 454092 497072
rect 459560 497020 459612 497072
rect 454132 496952 454184 497004
rect 458088 496952 458140 497004
rect 452844 496884 452896 496936
rect 455144 496884 455196 496936
rect 455420 496884 455472 496936
rect 461032 496884 461084 496936
rect 451372 496816 451424 496868
rect 453672 496816 453724 496868
rect 454684 496816 454736 496868
rect 456616 496816 456668 496868
rect 448428 496068 448480 496120
rect 547880 496068 547932 496120
rect 449992 494708 450044 494760
rect 450728 494708 450780 494760
rect 361764 491308 361816 491360
rect 417424 491308 417476 491360
rect 518164 484372 518216 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 419080 480224 419132 480276
rect 396724 476076 396776 476128
rect 400864 476008 400916 476060
rect 516784 470568 516836 470620
rect 579620 470568 579672 470620
rect 400864 468188 400916 468240
rect 401968 468188 402020 468240
rect 401968 464992 402020 465044
rect 403624 464992 403676 465044
rect 515404 464380 515456 464432
rect 542360 464380 542412 464432
rect 449808 464312 449860 464364
rect 525800 464312 525852 464364
rect 488264 462952 488316 463004
rect 494060 462952 494112 463004
rect 527640 462952 527692 463004
rect 436100 462408 436152 462460
rect 554136 462408 554188 462460
rect 431960 462340 432012 462392
rect 551192 462340 551244 462392
rect 477408 461592 477460 461644
rect 521752 461592 521804 461644
rect 476028 461456 476080 461508
rect 477408 461456 477460 461508
rect 449900 460912 449952 460964
rect 524420 460912 524472 460964
rect 449716 460164 449768 460216
rect 485780 460164 485832 460216
rect 449624 458804 449676 458856
rect 488540 458804 488592 458856
rect 361764 458192 361816 458244
rect 383016 458192 383068 458244
rect 449440 457444 449492 457496
rect 487160 457444 487212 457496
rect 403624 456764 403676 456816
rect 408408 456696 408460 456748
rect 473728 456492 473780 456544
rect 476028 456492 476080 456544
rect 451924 455472 451976 455524
rect 480996 455472 481048 455524
rect 423588 455404 423640 455456
rect 473728 455404 473780 455456
rect 449532 454724 449584 454776
rect 481640 454724 481692 454776
rect 449348 454656 449400 454708
rect 484400 454656 484452 454708
rect 408500 452548 408552 452600
rect 410340 452548 410392 452600
rect 422484 447516 422536 447568
rect 423588 447516 423640 447568
rect 427452 447176 427504 447228
rect 446864 447176 446916 447228
rect 423588 447108 423640 447160
rect 443368 447108 443420 447160
rect 410340 447040 410392 447092
rect 413284 447040 413336 447092
rect 436100 445680 436152 445732
rect 437388 445680 437440 445732
rect 432696 444524 432748 444576
rect 445760 444524 445812 444576
rect 437296 444456 437348 444508
rect 445852 444456 445904 444508
rect 442632 444388 442684 444440
rect 445944 444388 445996 444440
rect 443368 444320 443420 444372
rect 447876 444320 447928 444372
rect 413284 438268 413336 438320
rect 414756 438268 414808 438320
rect 361764 436092 361816 436144
rect 419172 436092 419224 436144
rect 574744 430584 574796 430636
rect 579620 430584 579672 430636
rect 456892 429972 456944 430024
rect 474280 429972 474332 430024
rect 458180 429904 458232 429956
rect 476948 429904 477000 429956
rect 458364 429836 458416 429888
rect 479340 429836 479392 429888
rect 479524 429836 479576 429888
rect 484952 429836 485004 429888
rect 486424 429156 486476 429208
rect 487620 429156 487672 429208
rect 457444 428408 457496 428460
rect 471612 428408 471664 428460
rect 414756 426368 414808 426420
rect 417516 426368 417568 426420
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 502984 423512 503036 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 444196 423376 444248 423428
rect 447784 423376 447836 423428
rect 483020 423376 483072 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 485780 423308 485832 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 487160 423240 487212 423292
rect 528928 423240 528980 423292
rect 488540 423172 488592 423224
rect 531504 423172 531556 423224
rect 496820 423104 496872 423156
rect 545672 423104 545724 423156
rect 498200 423036 498252 423088
rect 548248 423036 548300 423088
rect 499580 422968 499632 423020
rect 550824 422968 550876 423020
rect 501052 422900 501104 422952
rect 553400 422900 553452 422952
rect 483112 421540 483164 421592
rect 521200 421540 521252 421592
rect 417516 420452 417568 420504
rect 424324 420452 424376 420504
rect 494060 420180 494112 420232
rect 541808 420180 541860 420232
rect 362408 418752 362460 418804
rect 443644 418752 443696 418804
rect 509884 418140 509936 418192
rect 579712 418140 579764 418192
rect 421472 417732 421524 417784
rect 503720 417732 503772 417784
rect 425980 417664 426032 417716
rect 507860 417664 507912 417716
rect 425336 417596 425388 417648
rect 507952 417596 508004 417648
rect 424048 417528 424100 417580
rect 506480 417528 506532 417580
rect 424692 417460 424744 417512
rect 506572 417460 506624 417512
rect 422116 417392 422168 417444
rect 503996 417392 504048 417444
rect 362316 416032 362368 416084
rect 440884 416032 440936 416084
rect 361580 413992 361632 414044
rect 442264 413992 442316 414044
rect 362224 413244 362276 413296
rect 436744 413244 436796 413296
rect 361580 402976 361632 403028
rect 439504 402976 439556 403028
rect 502616 402228 502668 402280
rect 557540 402228 557592 402280
rect 497464 400868 497516 400920
rect 546500 400868 546552 400920
rect 494152 399440 494204 399492
rect 539600 399440 539652 399492
rect 492680 398080 492732 398132
rect 538220 398080 538272 398132
rect 492772 396720 492824 396772
rect 536840 396720 536892 396772
rect 460940 395292 460992 395344
rect 490012 395292 490064 395344
rect 491576 395292 491628 395344
rect 535460 395292 535512 395344
rect 461032 393932 461084 393984
rect 486424 393932 486476 393984
rect 491392 393932 491444 393984
rect 534172 393932 534224 393984
rect 463608 392572 463660 392624
rect 481640 392572 481692 392624
rect 490564 392572 490616 392624
rect 534080 392572 534132 392624
rect 361580 391960 361632 392012
rect 440976 391960 441028 392012
rect 450084 391280 450136 391332
rect 491116 391280 491168 391332
rect 496452 391280 496504 391332
rect 543740 391280 543792 391332
rect 422392 391212 422444 391264
rect 506020 391212 506072 391264
rect 460388 389852 460440 389904
rect 479524 389852 479576 389904
rect 495716 389852 495768 389904
rect 542360 389852 542412 389904
rect 422300 389784 422352 389836
rect 505284 389784 505336 389836
rect 449992 389240 450044 389292
rect 450728 389240 450780 389292
rect 454040 389240 454092 389292
rect 454868 389240 454920 389292
rect 460940 389240 460992 389292
rect 461492 389240 461544 389292
rect 483020 389240 483072 389292
rect 483572 389240 483624 389292
rect 492680 389240 492732 389292
rect 493140 389240 493192 389292
rect 494060 389240 494112 389292
rect 494612 389240 494664 389292
rect 507860 389240 507912 389292
rect 508596 389240 508648 389292
rect 453764 389104 453816 389156
rect 454684 389104 454736 389156
rect 456708 389104 456760 389156
rect 457444 389104 457496 389156
rect 468576 389104 468628 389156
rect 469220 389104 469272 389156
rect 469864 388900 469916 388952
rect 478052 388900 478104 388952
rect 484676 388900 484728 388952
rect 502984 388900 503036 388952
rect 499396 388832 499448 388884
rect 522304 388832 522356 388884
rect 468484 388764 468536 388816
rect 478788 388764 478840 388816
rect 500868 388764 500920 388816
rect 523684 388764 523736 388816
rect 459652 388696 459704 388748
rect 463608 388696 463660 388748
rect 468760 388696 468812 388748
rect 480260 388696 480312 388748
rect 502340 388696 502392 388748
rect 526444 388696 526496 388748
rect 461676 388628 461728 388680
rect 468484 388628 468536 388680
rect 468668 388628 468720 388680
rect 482468 388628 482520 388680
rect 485412 388628 485464 388680
rect 524420 388628 524472 388680
rect 461584 388560 461636 388612
rect 476580 388560 476632 388612
rect 486884 388560 486936 388612
rect 527180 388560 527232 388612
rect 465724 388492 465776 388544
rect 481732 388492 481784 388544
rect 489828 388492 489880 388544
rect 530584 388492 530636 388544
rect 448428 388424 448480 388476
rect 461768 388424 461820 388476
rect 464344 388424 464396 388476
rect 480996 388424 481048 388476
rect 488356 388424 488408 388476
rect 529204 388424 529256 388476
rect 462964 388152 463016 388204
rect 469956 388152 470008 388204
rect 466460 387744 466512 387796
rect 467380 387744 467432 387796
rect 450268 387132 450320 387184
rect 491300 387132 491352 387184
rect 449164 387064 449216 387116
rect 513380 387064 513432 387116
rect 447876 386588 447928 386640
rect 553952 386588 554004 386640
rect 382924 386520 382976 386572
rect 512184 386520 512236 386572
rect 380256 386452 380308 386504
rect 512276 386452 512328 386504
rect 380164 386384 380216 386436
rect 512000 386384 512052 386436
rect 447784 385976 447836 386028
rect 451924 385976 451976 386028
rect 447600 385364 447652 385416
rect 453304 385364 453356 385416
rect 447692 385092 447744 385144
rect 563428 385092 563480 385144
rect 374644 385024 374696 385076
rect 512092 385024 512144 385076
rect 364984 384956 365036 385008
rect 447140 384956 447192 385008
rect 512736 383732 512788 383784
rect 534724 383732 534776 383784
rect 513288 383664 513340 383716
rect 548524 383664 548576 383716
rect 381544 383596 381596 383648
rect 447140 383596 447192 383648
rect 406384 383528 406436 383580
rect 447232 383528 447284 383580
rect 513196 382440 513248 382492
rect 518348 382440 518400 382492
rect 513288 382372 513340 382424
rect 519636 382372 519688 382424
rect 512920 382236 512972 382288
rect 522304 382236 522356 382288
rect 378784 382168 378836 382220
rect 447140 382168 447192 382220
rect 407764 382100 407816 382152
rect 447232 382100 447284 382152
rect 512368 381080 512420 381132
rect 515496 381080 515548 381132
rect 361580 380876 361632 380928
rect 442356 380876 442408 380928
rect 513288 380876 513340 380928
rect 548616 380876 548668 380928
rect 376024 380808 376076 380860
rect 447140 380808 447192 380860
rect 410524 380740 410576 380792
rect 447232 380740 447284 380792
rect 512092 380400 512144 380452
rect 512460 380400 512512 380452
rect 512092 380128 512144 380180
rect 514116 380128 514168 380180
rect 512828 379516 512880 379568
rect 544384 379516 544436 379568
rect 371884 379448 371936 379500
rect 447232 379448 447284 379500
rect 374736 379380 374788 379432
rect 447140 379380 447192 379432
rect 512184 378292 512236 378344
rect 523684 378292 523736 378344
rect 513288 378224 513340 378276
rect 547144 378224 547196 378276
rect 514024 378156 514076 378208
rect 579620 378156 579672 378208
rect 367744 378088 367796 378140
rect 447232 378088 447284 378140
rect 370504 378020 370556 378072
rect 447140 378020 447192 378072
rect 513196 376864 513248 376916
rect 517520 376864 517572 376916
rect 363696 376660 363748 376712
rect 447232 376660 447284 376712
rect 363604 376592 363656 376644
rect 447140 376592 447192 376644
rect 512368 375980 512420 376032
rect 549904 375980 549956 376032
rect 363788 375300 363840 375352
rect 447140 375300 447192 375352
rect 411904 375232 411956 375284
rect 447232 375232 447284 375284
rect 512736 374144 512788 374196
rect 516140 374144 516192 374196
rect 414664 373940 414716 373992
rect 447140 373940 447192 373992
rect 416136 373872 416188 373924
rect 447232 373872 447284 373924
rect 512828 372648 512880 372700
rect 517612 372648 517664 372700
rect 513288 372580 513340 372632
rect 521660 372580 521712 372632
rect 417424 372512 417476 372564
rect 447140 372512 447192 372564
rect 419080 372444 419132 372496
rect 447232 372444 447284 372496
rect 512552 371220 512604 371272
rect 517704 371220 517756 371272
rect 383016 371152 383068 371204
rect 447232 371152 447284 371204
rect 436744 371084 436796 371136
rect 447140 371084 447192 371136
rect 512000 370064 512052 370116
rect 514208 370064 514260 370116
rect 513288 369996 513340 370048
rect 521752 369996 521804 370048
rect 512092 369928 512144 369980
rect 514944 369928 514996 369980
rect 361580 369860 361632 369912
rect 444012 369860 444064 369912
rect 419172 369792 419224 369844
rect 447232 369792 447284 369844
rect 440884 369724 440936 369776
rect 447140 369724 447192 369776
rect 513012 368568 513064 368620
rect 518900 368568 518952 368620
rect 443644 368432 443696 368484
rect 447140 368432 447192 368484
rect 442264 368364 442316 368416
rect 447232 368364 447284 368416
rect 512644 367208 512696 367260
rect 520280 367208 520332 367260
rect 439504 367004 439556 367056
rect 447140 367004 447192 367056
rect 440976 366936 441028 366988
rect 447232 366936 447284 366988
rect 512460 365848 512512 365900
rect 515588 365848 515640 365900
rect 444012 365644 444064 365696
rect 447140 365644 447192 365696
rect 442356 365576 442408 365628
rect 447232 365576 447284 365628
rect 512092 364488 512144 364540
rect 514852 364488 514904 364540
rect 570604 364352 570656 364404
rect 580172 364352 580224 364404
rect 513288 363060 513340 363112
rect 518256 363060 518308 363112
rect 442264 362992 442316 363044
rect 447232 362992 447284 363044
rect 512000 362992 512052 363044
rect 515036 362992 515088 363044
rect 432604 362924 432656 362976
rect 447140 362924 447192 362976
rect 512000 362176 512052 362228
rect 513748 362176 513800 362228
rect 513288 362040 513340 362092
rect 518992 362040 519044 362092
rect 513104 361768 513156 361820
rect 516876 361768 516928 361820
rect 443644 361632 443696 361684
rect 447232 361632 447284 361684
rect 435456 361564 435508 361616
rect 447140 361564 447192 361616
rect 442448 360272 442500 360324
rect 447232 360272 447284 360324
rect 513288 360272 513340 360324
rect 520372 360272 520424 360324
rect 439596 360204 439648 360256
rect 447140 360204 447192 360256
rect 547144 359184 547196 359236
rect 552296 359184 552348 359236
rect 548616 359116 548668 359168
rect 558184 359116 558236 359168
rect 544384 359048 544436 359100
rect 553768 359048 553820 359100
rect 548524 358980 548576 359032
rect 565544 358980 565596 359032
rect 523684 358912 523736 358964
rect 550824 358912 550876 358964
rect 441068 358844 441120 358896
rect 447232 358844 447284 358896
rect 513288 358844 513340 358896
rect 519176 358844 519228 358896
rect 534724 358844 534776 358896
rect 567016 358844 567068 358896
rect 436836 358776 436888 358828
rect 447140 358776 447192 358828
rect 514116 358776 514168 358828
rect 555240 358776 555292 358828
rect 549904 358708 549956 358760
rect 556712 358708 556764 358760
rect 519636 358640 519688 358692
rect 562600 358640 562652 358692
rect 518348 358572 518400 358624
rect 561128 358572 561180 358624
rect 522304 358504 522356 358556
rect 564072 358504 564124 358556
rect 515496 358436 515548 358488
rect 559656 358436 559708 358488
rect 512092 357620 512144 357672
rect 519268 357620 519320 357672
rect 512092 357416 512144 357468
rect 513840 357416 513892 357468
rect 512092 356328 512144 356380
rect 513656 356328 513708 356380
rect 512736 356124 512788 356176
rect 521844 356124 521896 356176
rect 513288 354764 513340 354816
rect 519452 354764 519504 354816
rect 513196 354696 513248 354748
rect 521936 354696 521988 354748
rect 512092 353744 512144 353796
rect 515128 353744 515180 353796
rect 513288 353268 513340 353320
rect 519084 353268 519136 353320
rect 512920 352112 512972 352164
rect 516324 352112 516376 352164
rect 424324 352044 424376 352096
rect 426900 352044 426952 352096
rect 394700 351908 394752 351960
rect 447140 351908 447192 351960
rect 513288 351908 513340 351960
rect 522028 351908 522080 351960
rect 512828 351432 512880 351484
rect 517888 351432 517940 351484
rect 512092 350752 512144 350804
rect 515220 350752 515272 350804
rect 405740 350548 405792 350600
rect 447140 350548 447192 350600
rect 513012 349256 513064 349308
rect 519360 349256 519412 349308
rect 512092 349188 512144 349240
rect 513932 349188 513984 349240
rect 446864 349052 446916 349104
rect 447600 349052 447652 349104
rect 432788 348372 432840 348424
rect 442264 348372 442316 348424
rect 512828 347896 512880 347948
rect 516232 347896 516284 347948
rect 361764 347760 361816 347812
rect 402244 347760 402296 347812
rect 512920 347760 512972 347812
rect 516508 347760 516560 347812
rect 362224 347692 362276 347744
rect 447140 347692 447192 347744
rect 426900 347624 426952 347676
rect 430580 347624 430632 347676
rect 513288 346672 513340 346724
rect 517796 346672 517848 346724
rect 512828 346536 512880 346588
rect 517980 346536 518032 346588
rect 512644 346400 512696 346452
rect 515312 346400 515364 346452
rect 512092 345924 512144 345976
rect 514116 345924 514168 345976
rect 432788 344292 432840 344344
rect 443644 344292 443696 344344
rect 512644 344224 512696 344276
rect 515496 344224 515548 344276
rect 513288 343952 513340 344004
rect 518072 343952 518124 344004
rect 512828 343816 512880 343868
rect 516416 343816 516468 343868
rect 402244 342864 402296 342916
rect 402980 342864 403032 342916
rect 447876 342864 447928 342916
rect 430580 342184 430632 342236
rect 432696 342184 432748 342236
rect 513288 341232 513340 341284
rect 519636 341232 519688 341284
rect 444104 340960 444156 341012
rect 447232 340960 447284 341012
rect 513012 340960 513064 341012
rect 516600 340960 516652 341012
rect 361764 340892 361816 340944
rect 447140 340892 447192 340944
rect 513288 339872 513340 339924
rect 520556 339872 520608 339924
rect 442356 339532 442408 339584
rect 447232 339532 447284 339584
rect 513012 339532 513064 339584
rect 516692 339532 516744 339584
rect 399484 339464 399536 339516
rect 447140 339464 447192 339516
rect 513196 339464 513248 339516
rect 522120 339464 522172 339516
rect 401600 339396 401652 339448
rect 402980 339396 403032 339448
rect 412640 338716 412692 338768
rect 449164 338716 449216 338768
rect 513288 338240 513340 338292
rect 519728 338240 519780 338292
rect 435364 338172 435416 338224
rect 447140 338172 447192 338224
rect 385776 338104 385828 338156
rect 447232 338104 447284 338156
rect 513196 338104 513248 338156
rect 520464 338104 520516 338156
rect 513196 337424 513248 337476
rect 518348 337424 518400 337476
rect 416780 336880 416832 336932
rect 431408 336880 431460 336932
rect 424140 336812 424192 336864
rect 429936 336812 429988 336864
rect 443828 336812 443880 336864
rect 447232 336812 447284 336864
rect 513288 336812 513340 336864
rect 520648 336812 520700 336864
rect 420460 336744 420512 336796
rect 439780 336744 439832 336796
rect 440976 336744 441028 336796
rect 447140 336744 447192 336796
rect 513196 336744 513248 336796
rect 522212 336744 522264 336796
rect 432696 336676 432748 336728
rect 433984 336676 434036 336728
rect 418988 336268 419040 336320
rect 442540 336268 442592 336320
rect 416044 336200 416096 336252
rect 439688 336200 439740 336252
rect 418896 336132 418948 336184
rect 442632 336132 442684 336184
rect 418804 336064 418856 336116
rect 442724 336064 442776 336116
rect 362224 335996 362276 336048
rect 444104 335996 444156 336048
rect 513196 335792 513248 335844
rect 516968 335792 517020 335844
rect 442264 335452 442316 335504
rect 447324 335452 447376 335504
rect 409420 335384 409472 335436
rect 431316 335384 431368 335436
rect 413100 335316 413152 335368
rect 435548 335316 435600 335368
rect 439504 335316 439556 335368
rect 447232 335316 447284 335368
rect 513288 335316 513340 335368
rect 522304 335316 522356 335368
rect 420368 335044 420420 335096
rect 420552 335044 420604 335096
rect 442172 335044 442224 335096
rect 420644 334976 420696 335028
rect 444932 334976 444984 335028
rect 446956 334908 447008 334960
rect 420276 334840 420328 334892
rect 446864 334840 446916 334892
rect 420828 334772 420880 334824
rect 449440 334772 449492 334824
rect 420736 334704 420788 334756
rect 449532 334704 449584 334756
rect 420184 334636 420236 334688
rect 449072 334636 449124 334688
rect 420092 334568 420144 334620
rect 449348 334568 449400 334620
rect 428096 334364 428148 334416
rect 437020 334364 437072 334416
rect 513196 334296 513248 334348
rect 520740 334296 520792 334348
rect 443736 334024 443788 334076
rect 447324 334024 447376 334076
rect 364064 333956 364116 334008
rect 447232 333956 447284 334008
rect 513288 333956 513340 334008
rect 522396 333956 522448 334008
rect 440884 332664 440936 332716
rect 447324 332664 447376 332716
rect 429844 332596 429896 332648
rect 447232 332596 447284 332648
rect 432880 331848 432932 331900
rect 442448 331848 442500 331900
rect 436744 331304 436796 331356
rect 447508 331304 447560 331356
rect 443644 331236 443696 331288
rect 447232 331236 447284 331288
rect 445944 331168 445996 331220
rect 447324 331168 447376 331220
rect 440148 330556 440200 330608
rect 445944 330556 445996 330608
rect 432604 330216 432656 330268
rect 441068 330216 441120 330268
rect 442908 330080 442960 330132
rect 445852 330080 445904 330132
rect 447232 330080 447284 330132
rect 512736 330080 512788 330132
rect 514760 330080 514812 330132
rect 438768 329060 438820 329112
rect 445760 329060 445812 329112
rect 447232 329060 447284 329112
rect 432972 328652 433024 328704
rect 435456 328652 435508 328704
rect 436008 328448 436060 328500
rect 447232 328448 447284 328500
rect 433984 328380 434036 328432
rect 436928 328380 436980 328432
rect 437020 328380 437072 328432
rect 447324 328380 447376 328432
rect 448336 328380 448388 328432
rect 431224 327088 431276 327140
rect 447232 327088 447284 327140
rect 439780 327020 439832 327072
rect 447324 327020 447376 327072
rect 448060 327020 448112 327072
rect 429936 326340 429988 326392
rect 440332 326340 440384 326392
rect 447232 326340 447284 326392
rect 431408 325592 431460 325644
rect 448152 325592 448204 325644
rect 435548 325456 435600 325508
rect 447968 325456 448020 325508
rect 436928 324980 436980 325032
rect 440240 324980 440292 325032
rect 511908 324300 511960 324352
rect 580172 324300 580224 324352
rect 440240 323620 440292 323672
rect 447232 323620 447284 323672
rect 431316 323552 431368 323604
rect 449256 323552 449308 323604
rect 510528 323552 510580 323604
rect 580264 323552 580316 323604
rect 507492 322532 507544 322584
rect 509608 322532 509660 322584
rect 442816 322396 442868 322448
rect 449992 322396 450044 322448
rect 446588 322328 446640 322380
rect 470140 322328 470192 322380
rect 446956 322260 447008 322312
rect 483112 322260 483164 322312
rect 447232 322192 447284 322244
rect 449900 322192 449952 322244
rect 449992 322192 450044 322244
rect 479800 322192 479852 322244
rect 507216 322192 507268 322244
rect 514760 322192 514812 322244
rect 445668 322124 445720 322176
rect 471796 322124 471848 322176
rect 477868 322124 477920 322176
rect 514024 322124 514076 322176
rect 444932 322056 444984 322108
rect 482560 322056 482612 322108
rect 504088 322056 504140 322108
rect 511264 322056 511316 322108
rect 439688 321988 439740 322040
rect 470692 321988 470744 322040
rect 478420 321988 478472 322040
rect 518164 321988 518216 322040
rect 450636 321920 450688 321972
rect 460756 321920 460808 321972
rect 467656 321920 467708 321972
rect 446772 321852 446824 321904
rect 461952 321852 462004 321904
rect 468300 321852 468352 321904
rect 504088 321852 504140 321904
rect 507400 321920 507452 321972
rect 509792 321920 509844 321972
rect 509884 321852 509936 321904
rect 442172 321784 442224 321836
rect 462504 321784 462556 321836
rect 467748 321784 467800 321836
rect 516784 321784 516836 321836
rect 457536 321716 457588 321768
rect 567844 321716 567896 321768
rect 458088 321648 458140 321700
rect 580356 321648 580408 321700
rect 457812 321580 457864 321632
rect 580448 321580 580500 321632
rect 456708 321512 456760 321564
rect 580724 321512 580776 321564
rect 456984 321444 457036 321496
rect 580632 321444 580684 321496
rect 458364 321376 458416 321428
rect 569224 321376 569276 321428
rect 445484 321308 445536 321360
rect 461400 321308 461452 321360
rect 468576 321308 468628 321360
rect 576124 321308 576176 321360
rect 445024 321240 445076 321292
rect 459468 321240 459520 321292
rect 467196 321240 467248 321292
rect 570604 321240 570656 321292
rect 446404 321172 446456 321224
rect 459192 321172 459244 321224
rect 477960 321172 478012 321224
rect 574744 321172 574796 321224
rect 479340 321104 479392 321156
rect 573364 321104 573416 321156
rect 445576 321036 445628 321088
rect 461124 321036 461176 321088
rect 468024 321036 468076 321088
rect 511356 321036 511408 321088
rect 450544 320968 450596 321020
rect 481272 320968 481324 321020
rect 507032 320968 507084 321020
rect 516876 320968 516928 321020
rect 445116 320900 445168 320952
rect 460020 320900 460072 320952
rect 460204 320900 460256 320952
rect 518256 320900 518308 320952
rect 449900 320832 449952 320884
rect 456800 320832 456852 320884
rect 459560 320832 459612 320884
rect 580540 320832 580592 320884
rect 446496 320764 446548 320816
rect 480168 320764 480220 320816
rect 507584 320764 507636 320816
rect 513380 320764 513432 320816
rect 442632 320696 442684 320748
rect 482100 320696 482152 320748
rect 507768 320696 507820 320748
rect 510068 320696 510120 320748
rect 442540 320628 442592 320680
rect 480720 320628 480772 320680
rect 457260 320084 457312 320136
rect 459560 320084 459612 320136
rect 479064 320084 479116 320136
rect 578884 320084 578936 320136
rect 456800 320016 456852 320068
rect 472992 320016 473044 320068
rect 478788 320016 478840 320068
rect 571984 320016 572036 320068
rect 446864 319948 446916 320000
rect 462228 319948 462280 320000
rect 469128 319948 469180 320000
rect 515404 319948 515456 320000
rect 450452 319880 450504 319932
rect 461676 319880 461728 319932
rect 478512 319880 478564 319932
rect 519544 319880 519596 319932
rect 444196 319812 444248 319864
rect 458916 319812 458968 319864
rect 468852 319812 468904 319864
rect 510528 319812 510580 319864
rect 449072 319744 449124 319796
rect 472440 319744 472492 319796
rect 477408 319744 477460 319796
rect 511908 319744 511960 319796
rect 446680 319676 446732 319728
rect 469956 319676 470008 319728
rect 501420 319676 501472 319728
rect 449532 319608 449584 319660
rect 472716 319608 472768 319660
rect 445300 319540 445352 319592
rect 480996 319540 481048 319592
rect 500316 319540 500368 319592
rect 445392 319472 445444 319524
rect 482928 319472 482980 319524
rect 502524 319472 502576 319524
rect 534724 319540 534776 319592
rect 538864 319472 538916 319524
rect 445208 319404 445260 319456
rect 470508 319404 470560 319456
rect 543740 319404 543792 319456
rect 449440 319336 449492 319388
rect 482376 319336 482428 319388
rect 449348 319268 449400 319320
rect 472164 319268 472216 319320
rect 449164 319200 449216 319252
rect 469680 319200 469732 319252
rect 473452 319200 473504 319252
rect 473728 319200 473780 319252
rect 496912 319200 496964 319252
rect 497464 319200 497516 319252
rect 501052 319200 501104 319252
rect 501604 319200 501656 319252
rect 454040 319132 454092 319184
rect 455236 319132 455288 319184
rect 454224 319064 454276 319116
rect 454684 319064 454736 319116
rect 455512 319064 455564 319116
rect 456064 319064 456116 319116
rect 462688 319064 462740 319116
rect 463516 319064 463568 319116
rect 463792 319064 463844 319116
rect 464896 319064 464948 319116
rect 465448 319064 465500 319116
rect 466000 319064 466052 319116
rect 475108 319064 475160 319116
rect 475936 319064 475988 319116
rect 476212 319064 476264 319116
rect 476764 319064 476816 319116
rect 483112 319064 483164 319116
rect 483940 319064 483992 319116
rect 484492 319064 484544 319116
rect 485596 319064 485648 319116
rect 495532 319064 495584 319116
rect 496360 319064 496412 319116
rect 499672 319064 499724 319116
rect 500776 319064 500828 319116
rect 504088 319064 504140 319116
rect 504916 319064 504968 319116
rect 454132 318996 454184 319048
rect 454960 318996 455012 319048
rect 462412 318996 462464 319048
rect 463240 318996 463292 319048
rect 465172 318996 465224 319048
rect 466276 318996 466328 319048
rect 474832 318996 474884 319048
rect 475660 318996 475712 319048
rect 480904 318996 480956 319048
rect 483756 318996 483808 319048
rect 498568 318928 498620 318980
rect 499396 318928 499448 318980
rect 485044 318792 485096 318844
rect 485320 318792 485372 318844
rect 444288 318724 444340 318776
rect 469404 318724 469456 318776
rect 477132 318316 477184 318368
rect 479524 318316 479576 318368
rect 432144 318112 432196 318164
rect 439596 318112 439648 318164
rect 456432 318112 456484 318164
rect 449624 318044 449676 318096
rect 456892 318044 456944 318096
rect 458824 318112 458876 318164
rect 487344 318112 487396 318164
rect 494796 318112 494848 318164
rect 540980 318112 541032 318164
rect 461584 318044 461636 318096
rect 459100 317976 459152 318028
rect 493968 318044 494020 318096
rect 495624 318044 495676 318096
rect 543280 318044 543332 318096
rect 448428 317024 448480 317076
rect 457812 317024 457864 317076
rect 447784 316956 447836 317008
rect 462780 316956 462832 317008
rect 500040 316956 500092 317008
rect 542636 316956 542688 317008
rect 457444 316888 457496 316940
rect 490932 316888 490984 316940
rect 498384 316888 498436 316940
rect 541072 316888 541124 316940
rect 453304 316820 453356 316872
rect 489552 316820 489604 316872
rect 490012 316820 490064 316872
rect 490288 316820 490340 316872
rect 493140 316820 493192 316872
rect 493324 316820 493376 316872
rect 495900 316820 495952 316872
rect 542452 316820 542504 316872
rect 454684 316752 454736 316804
rect 502340 316752 502392 316804
rect 450544 316684 450596 316736
rect 504732 316684 504784 316736
rect 486148 316616 486200 316668
rect 486700 316616 486752 316668
rect 487804 316616 487856 316668
rect 488356 316616 488408 316668
rect 488632 316616 488684 316668
rect 489736 316616 489788 316668
rect 492772 316616 492824 316668
rect 493600 316616 493652 316668
rect 494152 316616 494204 316668
rect 495256 316616 495308 316668
rect 485872 316548 485924 316600
rect 486424 316548 486476 316600
rect 490288 316548 490340 316600
rect 491116 316548 491168 316600
rect 464252 316004 464304 316056
rect 464436 316004 464488 316056
rect 361764 315936 361816 315988
rect 399484 315936 399536 315988
rect 499764 315460 499816 315512
rect 539692 315460 539744 315512
rect 458916 315392 458968 315444
rect 491392 315392 491444 315444
rect 496084 315392 496136 315444
rect 539600 315392 539652 315444
rect 450728 315324 450780 315376
rect 502984 315324 503036 315376
rect 450636 315256 450688 315308
rect 504364 315256 504416 315308
rect 469864 314644 469916 314696
rect 472348 314644 472400 314696
rect 501604 314032 501656 314084
rect 538956 314032 539008 314084
rect 459008 313964 459060 314016
rect 492312 313964 492364 314016
rect 495808 313964 495860 314016
rect 542544 313964 542596 314016
rect 450820 313896 450872 313948
rect 503904 313896 503956 313948
rect 466828 313216 466880 313268
rect 580172 313216 580224 313268
rect 465264 312536 465316 312588
rect 547144 312536 547196 312588
rect 487252 312128 487304 312180
rect 488080 312128 488132 312180
rect 451924 311244 451976 311296
rect 487896 311244 487948 311296
rect 501144 311244 501196 311296
rect 540336 311244 540388 311296
rect 456064 311176 456116 311228
rect 504180 311176 504232 311228
rect 455604 311108 455656 311160
rect 533344 311108 533396 311160
rect 452016 309816 452068 309868
rect 488816 309816 488868 309868
rect 475384 309748 475436 309800
rect 565084 309748 565136 309800
rect 446404 308456 446456 308508
rect 462964 308456 463016 308508
rect 453396 308388 453448 308440
rect 489184 308388 489236 308440
rect 478144 307776 478196 307828
rect 480904 307776 480956 307828
rect 432236 307708 432288 307760
rect 436836 307708 436888 307760
rect 485964 307096 486016 307148
rect 529940 307096 529992 307148
rect 475108 307028 475160 307080
rect 569224 307028 569276 307080
rect 384304 306280 384356 306332
rect 464068 306280 464120 306332
rect 386052 306212 386104 306264
rect 474280 306212 474332 306264
rect 384488 306144 384540 306196
rect 474004 306144 474056 306196
rect 384580 306076 384632 306128
rect 474924 306076 474976 306128
rect 381728 306008 381780 306060
rect 473728 306008 473780 306060
rect 384948 305940 385000 305992
rect 484768 305940 484820 305992
rect 384672 305872 384724 305924
rect 485136 305872 485188 305924
rect 381544 305804 381596 305856
rect 484584 305804 484636 305856
rect 426348 305736 426400 305788
rect 440240 305736 440292 305788
rect 455788 305736 455840 305788
rect 574744 305736 574796 305788
rect 360844 305668 360896 305720
rect 512276 305668 512328 305720
rect 360936 305600 360988 305652
rect 512552 305600 512604 305652
rect 384396 305532 384448 305584
rect 464436 305532 464488 305584
rect 385960 305464 386012 305516
rect 464160 305464 464212 305516
rect 452200 305396 452252 305448
rect 492956 305396 493008 305448
rect 3424 304988 3476 305040
rect 4804 304988 4856 305040
rect 361764 304920 361816 304972
rect 442356 304920 442408 304972
rect 486240 304444 486292 304496
rect 530032 304444 530084 304496
rect 385868 304376 385920 304428
rect 507032 304376 507084 304428
rect 362224 304308 362276 304360
rect 512736 304308 512788 304360
rect 361028 304240 361080 304292
rect 512184 304240 512236 304292
rect 463792 303560 463844 303612
rect 562324 303560 562376 303612
rect 379336 303492 379388 303544
rect 483664 303492 483716 303544
rect 486148 303492 486200 303544
rect 528560 303492 528612 303544
rect 376484 303424 376536 303476
rect 510896 303424 510948 303476
rect 376300 303356 376352 303408
rect 510988 303356 511040 303408
rect 379152 303288 379204 303340
rect 513932 303288 513984 303340
rect 379060 303220 379112 303272
rect 514116 303220 514168 303272
rect 378968 303152 379020 303204
rect 515312 303152 515364 303204
rect 376392 303084 376444 303136
rect 515220 303084 515272 303136
rect 376208 303016 376260 303068
rect 515128 303016 515180 303068
rect 373632 302948 373684 303000
rect 513840 302948 513892 303000
rect 361120 302880 361172 302932
rect 512368 302880 512420 302932
rect 379428 302812 379480 302864
rect 473452 302812 473504 302864
rect 378692 302744 378744 302796
rect 462412 302744 462464 302796
rect 382096 302676 382148 302728
rect 462688 302676 462740 302728
rect 378784 302608 378836 302660
rect 464344 302608 464396 302660
rect 3516 301928 3568 301980
rect 4896 301928 4948 301980
rect 476304 301588 476356 301640
rect 548524 301588 548576 301640
rect 407120 301520 407172 301572
rect 502432 301520 502484 301572
rect 371884 301452 371936 301504
rect 512460 301452 512512 301504
rect 373448 300772 373500 300824
rect 509424 300772 509476 300824
rect 370688 300704 370740 300756
rect 509332 300704 509384 300756
rect 370964 300636 371016 300688
rect 510804 300636 510856 300688
rect 371056 300568 371108 300620
rect 513564 300568 513616 300620
rect 370780 300500 370832 300552
rect 513748 300500 513800 300552
rect 367744 300432 367796 300484
rect 510712 300432 510764 300484
rect 370872 300364 370924 300416
rect 515036 300364 515088 300416
rect 368020 300296 368072 300348
rect 514944 300296 514996 300348
rect 365076 300228 365128 300280
rect 513472 300228 513524 300280
rect 367928 300160 367980 300212
rect 517704 300160 517756 300212
rect 367836 300092 367888 300144
rect 517612 300092 517664 300144
rect 375932 300024 375984 300076
rect 483112 300024 483164 300076
rect 465540 299956 465592 300008
rect 566464 299956 566516 300008
rect 376668 299888 376720 299940
rect 473544 299888 473596 299940
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 454776 297984 454828 298036
rect 502708 297984 502760 298036
rect 454316 297916 454368 297968
rect 563704 297916 563756 297968
rect 385684 297848 385736 297900
rect 516600 297848 516652 297900
rect 384856 297780 384908 297832
rect 516692 297780 516744 297832
rect 362500 297712 362552 297764
rect 507768 297712 507820 297764
rect 364984 297644 365036 297696
rect 511540 297644 511592 297696
rect 366548 297576 366600 297628
rect 517980 297576 518032 297628
rect 365260 297508 365312 297560
rect 517520 297508 517572 297560
rect 363696 297440 363748 297492
rect 516968 297440 517020 297492
rect 363788 297372 363840 297424
rect 518072 297372 518124 297424
rect 454224 295944 454276 295996
rect 573364 295944 573416 295996
rect 374736 295264 374788 295316
rect 514852 295264 514904 295316
rect 366732 295196 366784 295248
rect 509516 295196 509568 295248
rect 370596 295128 370648 295180
rect 513656 295128 513708 295180
rect 375012 295060 375064 295112
rect 518992 295060 519044 295112
rect 373356 294992 373408 295044
rect 519176 294992 519228 295044
rect 372252 294924 372304 294976
rect 520372 294924 520424 294976
rect 368112 294856 368164 294908
rect 516508 294856 516560 294908
rect 366456 294788 366508 294840
rect 516324 294788 516376 294840
rect 369308 294720 369360 294772
rect 519268 294720 519320 294772
rect 369216 294652 369268 294704
rect 519452 294652 519504 294704
rect 365444 294584 365496 294636
rect 517888 294584 517940 294636
rect 374828 294516 374880 294568
rect 515588 294516 515640 294568
rect 454132 294448 454184 294500
rect 578884 294448 578936 294500
rect 361764 293904 361816 293956
rect 385776 293904 385828 293956
rect 476488 293224 476540 293276
rect 537484 293224 537536 293276
rect 383292 292476 383344 292528
rect 507584 292476 507636 292528
rect 380532 292408 380584 292460
rect 507676 292408 507728 292460
rect 378600 292340 378652 292392
rect 507492 292340 507544 292392
rect 386328 292272 386380 292324
rect 520740 292272 520792 292324
rect 377680 292204 377732 292256
rect 514208 292204 514260 292256
rect 377588 292136 377640 292188
rect 516140 292136 516192 292188
rect 382004 292068 382056 292120
rect 520648 292068 520700 292120
rect 376576 292000 376628 292052
rect 520280 292000 520332 292052
rect 375104 291932 375156 291984
rect 518900 291932 518952 291984
rect 362316 291864 362368 291916
rect 519728 291864 519780 291916
rect 361212 291796 361264 291848
rect 520556 291796 520608 291848
rect 385776 291728 385828 291780
rect 507400 291728 507452 291780
rect 362592 291660 362644 291712
rect 443828 291660 443880 291712
rect 457536 291660 457588 291712
rect 490196 291660 490248 291712
rect 499120 291660 499172 291712
rect 541164 291660 541216 291712
rect 478236 291592 478288 291644
rect 483388 291592 483440 291644
rect 465356 291184 465408 291236
rect 469864 291184 469916 291236
rect 455512 290436 455564 290488
rect 571984 290436 572036 290488
rect 380440 289756 380492 289808
rect 519084 289756 519136 289808
rect 383200 289688 383252 289740
rect 521936 289688 521988 289740
rect 363972 289620 364024 289672
rect 507308 289620 507360 289672
rect 372068 289552 372120 289604
rect 516232 289552 516284 289604
rect 366364 289484 366416 289536
rect 510620 289484 510672 289536
rect 374920 289416 374972 289468
rect 519360 289416 519412 289468
rect 377496 289348 377548 289400
rect 522028 289348 522080 289400
rect 369400 289280 369452 289332
rect 517796 289280 517848 289332
rect 366640 289212 366692 289264
rect 516416 289212 516468 289264
rect 369124 289144 369176 289196
rect 521752 289144 521804 289196
rect 363880 289076 363932 289128
rect 519636 289076 519688 289128
rect 386236 289008 386288 289060
rect 521844 289008 521896 289060
rect 441068 288940 441120 288992
rect 446404 288940 446456 288992
rect 454132 288940 454184 288992
rect 465356 288940 465408 288992
rect 474832 288940 474884 288992
rect 544384 288940 544436 288992
rect 454040 287648 454092 287700
rect 576124 287648 576176 287700
rect 485872 286832 485924 286884
rect 530124 286832 530176 286884
rect 383108 286764 383160 286816
rect 507124 286764 507176 286816
rect 377404 286696 377456 286748
rect 507216 286696 507268 286748
rect 386144 286628 386196 286680
rect 522396 286628 522448 286680
rect 381912 286560 381964 286612
rect 522304 286560 522356 286612
rect 378876 286492 378928 286544
rect 522212 286492 522264 286544
rect 376116 286424 376168 286476
rect 520464 286424 520516 286476
rect 373264 286356 373316 286408
rect 522120 286356 522172 286408
rect 372344 286288 372396 286340
rect 521660 286288 521712 286340
rect 475384 285676 475436 285728
rect 478144 285676 478196 285728
rect 453488 284996 453540 285048
rect 487804 284996 487856 285048
rect 501328 284996 501380 285048
rect 539048 284996 539100 285048
rect 476212 284928 476264 284980
rect 570604 284928 570656 284980
rect 452108 283636 452160 283688
rect 487252 283636 487304 283688
rect 497004 283636 497056 283688
rect 539784 283636 539836 283688
rect 449164 283568 449216 283620
rect 454132 283568 454184 283620
rect 465724 283568 465776 283620
rect 554044 283568 554096 283620
rect 361764 282820 361816 282872
rect 435364 282820 435416 282872
rect 459284 282208 459336 282260
rect 494244 282208 494296 282260
rect 465448 282140 465500 282192
rect 555424 282140 555476 282192
rect 445024 281868 445076 281920
rect 447784 281868 447836 281920
rect 452384 280848 452436 280900
rect 493140 280848 493192 280900
rect 465172 280780 465224 280832
rect 559564 280780 559616 280832
rect 454960 279420 455012 279472
rect 487528 279420 487580 279472
rect 501052 279420 501104 279472
rect 541532 279420 541584 279472
rect 453580 277992 453632 278044
rect 492772 277992 492824 278044
rect 499948 277992 500000 278044
rect 540244 277992 540296 278044
rect 456340 276768 456392 276820
rect 492220 276768 492272 276820
rect 498844 276768 498896 276820
rect 539968 276768 540020 276820
rect 449808 276700 449860 276752
rect 536840 276700 536892 276752
rect 359464 276632 359516 276684
rect 512000 276632 512052 276684
rect 465724 275476 465776 275528
rect 478236 275476 478288 275528
rect 457628 275408 457680 275460
rect 488632 275408 488684 275460
rect 457720 275340 457772 275392
rect 491944 275340 491996 275392
rect 383384 275272 383436 275324
rect 475200 275272 475252 275324
rect 497464 275272 497516 275324
rect 541440 275272 541492 275324
rect 443828 274660 443880 274712
rect 449164 274660 449216 274712
rect 460296 274048 460348 274100
rect 494520 274048 494572 274100
rect 455052 273980 455104 274032
rect 491668 273980 491720 274032
rect 368204 273912 368256 273964
rect 485044 273912 485096 273964
rect 497188 273912 497240 273964
rect 541256 273912 541308 273964
rect 479524 273164 479576 273216
rect 580172 273164 580224 273216
rect 459192 272552 459244 272604
rect 490564 272552 490616 272604
rect 433984 272484 434036 272536
rect 445024 272484 445076 272536
rect 453672 272484 453724 272536
rect 493048 272484 493100 272536
rect 498568 272484 498620 272536
rect 540152 272484 540204 272536
rect 456248 271260 456300 271312
rect 490288 271260 490340 271312
rect 456156 271192 456208 271244
rect 490012 271192 490064 271244
rect 498292 271192 498344 271244
rect 540060 271192 540112 271244
rect 452292 271124 452344 271176
rect 488908 271124 488960 271176
rect 496912 271124 496964 271176
rect 541348 271124 541400 271176
rect 455144 269900 455196 269952
rect 486424 269900 486476 269952
rect 494152 269900 494204 269952
rect 542728 269900 542780 269952
rect 466552 269832 466604 269884
rect 580264 269832 580316 269884
rect 359556 269764 359608 269816
rect 512092 269764 512144 269816
rect 459376 268540 459428 268592
rect 465724 268540 465776 268592
rect 499672 268540 499724 268592
rect 542912 268540 542964 268592
rect 445024 268472 445076 268524
rect 475384 268472 475436 268524
rect 495532 268472 495584 268524
rect 542820 268472 542872 268524
rect 457076 268404 457128 268456
rect 505192 268404 505244 268456
rect 454868 268336 454920 268388
rect 504088 268336 504140 268388
rect 424324 266976 424376 267028
rect 433984 266976 434036 267028
rect 449716 263508 449768 263560
rect 456800 263508 456852 263560
rect 361764 260788 361816 260840
rect 440976 260788 441028 260840
rect 433984 260108 434036 260160
rect 443828 260108 443880 260160
rect 3608 259360 3660 259412
rect 4988 259360 5040 259412
rect 433708 255280 433760 255332
rect 441068 255280 441120 255332
rect 361764 249704 361816 249756
rect 439504 249704 439556 249756
rect 446404 249024 446456 249076
rect 456800 249024 456852 249076
rect 431316 248412 431368 248464
rect 433708 248412 433760 248464
rect 571984 245556 572036 245608
rect 580172 245556 580224 245608
rect 3884 241408 3936 241460
rect 5080 241408 5132 241460
rect 361764 238688 361816 238740
rect 442264 238688 442316 238740
rect 570604 233180 570656 233232
rect 579988 233180 580040 233232
rect 421564 230460 421616 230512
rect 424324 230460 424376 230512
rect 453856 227740 453908 227792
rect 459376 227740 459428 227792
rect 361764 227672 361816 227724
rect 443736 227672 443788 227724
rect 432604 221416 432656 221468
rect 453856 221416 453908 221468
rect 425704 220804 425756 220856
rect 433984 220804 434036 220856
rect 414664 220056 414716 220108
rect 447968 220056 448020 220108
rect 459468 220056 459520 220108
rect 559564 219376 559616 219428
rect 580172 219376 580224 219428
rect 3976 218016 4028 218068
rect 5172 218016 5224 218068
rect 413284 218016 413336 218068
rect 421564 218016 421616 218068
rect 361672 216316 361724 216368
rect 364064 216316 364116 216368
rect 425796 213188 425848 213240
rect 445024 213188 445076 213240
rect 424324 209040 424376 209092
rect 432604 209040 432656 209092
rect 406292 207612 406344 207664
rect 425796 207612 425848 207664
rect 574744 206932 574796 206984
rect 579804 206932 579856 206984
rect 411260 206252 411312 206304
rect 450912 206252 450964 206304
rect 456800 206252 456852 206304
rect 361764 205572 361816 205624
rect 440884 205572 440936 205624
rect 401600 200744 401652 200796
rect 406292 200744 406344 200796
rect 421564 200744 421616 200796
rect 431316 200744 431368 200796
rect 456800 200744 456852 200796
rect 479524 200744 479576 200796
rect 459468 199384 459520 199436
rect 485780 199384 485832 199436
rect 406384 195236 406436 195288
rect 424324 195236 424376 195288
rect 422852 194692 422904 194744
rect 425704 194692 425756 194744
rect 361764 194488 361816 194540
rect 429844 194488 429896 194540
rect 388444 193808 388496 193860
rect 401600 193808 401652 193860
rect 537484 193128 537536 193180
rect 580172 193128 580224 193180
rect 411352 191088 411404 191140
rect 422852 191088 422904 191140
rect 402244 188368 402296 188420
rect 406384 188368 406436 188420
rect 398840 188300 398892 188352
rect 411352 188300 411404 188352
rect 410524 186260 410576 186312
rect 413284 186260 413336 186312
rect 366824 185580 366876 185632
rect 388444 185580 388496 185632
rect 361764 183472 361816 183524
rect 436744 183472 436796 183524
rect 391112 181432 391164 181484
rect 398840 181432 398892 181484
rect 416044 179392 416096 179444
rect 421564 179392 421616 179444
rect 555424 179324 555476 179376
rect 580172 179324 580224 179376
rect 396724 178644 396776 178696
rect 410524 178644 410576 178696
rect 398104 178032 398156 178084
rect 402244 178032 402296 178084
rect 361304 175924 361356 175976
rect 391112 175924 391164 175976
rect 364064 172524 364116 172576
rect 366824 172524 366876 172576
rect 361764 171776 361816 171828
rect 443644 171776 443696 171828
rect 524420 171776 524472 171828
rect 393964 167016 394016 167068
rect 396724 167016 396776 167068
rect 533344 166948 533396 167000
rect 580172 166948 580224 167000
rect 410248 164840 410300 164892
rect 416044 164840 416096 164892
rect 447416 163548 447468 163600
rect 461584 163548 461636 163600
rect 445668 163480 445720 163532
rect 446404 163480 446456 163532
rect 447508 163480 447560 163532
rect 528560 163480 528612 163532
rect 359648 163004 359700 163056
rect 364064 163004 364116 163056
rect 407764 162256 407816 162308
rect 410248 162256 410300 162308
rect 418712 162120 418764 162172
rect 458088 162120 458140 162172
rect 489920 162120 489972 162172
rect 403624 161712 403676 161764
rect 431224 161712 431276 161764
rect 426348 161644 426400 161696
rect 496820 161644 496872 161696
rect 421564 161576 421616 161628
rect 494060 161576 494112 161628
rect 407856 161508 407908 161560
rect 438768 161508 438820 161560
rect 513380 161508 513432 161560
rect 362592 161440 362644 161492
rect 441620 161440 441672 161492
rect 442908 161440 442960 161492
rect 517520 161440 517572 161492
rect 361764 161372 361816 161424
rect 440148 161372 440200 161424
rect 440148 160692 440200 160744
rect 521660 160692 521712 160744
rect 383476 160420 383528 160472
rect 418160 160420 418212 160472
rect 410616 160352 410668 160404
rect 385592 160284 385644 160336
rect 414756 160284 414808 160336
rect 435272 160284 435324 160336
rect 436008 160284 436060 160336
rect 450912 160284 450964 160336
rect 410524 160216 410576 160268
rect 428004 160216 428056 160268
rect 428648 160216 428700 160268
rect 461676 160216 461728 160268
rect 395344 160148 395396 160200
rect 398104 160148 398156 160200
rect 406384 160148 406436 160200
rect 445208 160148 445260 160200
rect 445668 160148 445720 160200
rect 483664 160148 483716 160200
rect 381360 160080 381412 160132
rect 425014 160080 425066 160132
rect 426348 160080 426400 160132
rect 431638 160080 431690 160132
rect 504364 160080 504416 160132
rect 398104 159332 398156 159384
rect 407764 159332 407816 159384
rect 364064 158720 364116 158772
rect 421380 159332 421432 159384
rect 451556 158380 451608 158432
rect 455144 158380 455196 158432
rect 365536 157972 365588 158024
rect 393964 157972 394016 158024
rect 451740 157292 451792 157344
rect 460296 157292 460348 157344
rect 452568 155524 452620 155576
rect 459284 155524 459336 155576
rect 451740 154504 451792 154556
rect 459100 154504 459152 154556
rect 451648 153144 451700 153196
rect 453580 153144 453632 153196
rect 548524 153144 548576 153196
rect 580172 153144 580224 153196
rect 451464 151444 451516 151496
rect 453672 151444 453724 151496
rect 393964 150424 394016 150476
rect 398104 150424 398156 150476
rect 390192 149336 390244 149388
rect 395344 149336 395396 149388
rect 452568 147500 452620 147552
rect 456340 147500 456392 147552
rect 452568 146004 452620 146056
rect 459008 146004 459060 146056
rect 452568 144644 452620 144696
rect 457720 144644 457772 144696
rect 504364 143488 504416 143540
rect 505652 143488 505704 143540
rect 452568 143284 452620 143336
rect 455052 143284 455104 143336
rect 387064 143080 387116 143132
rect 390192 143080 390244 143132
rect 461676 142944 461728 142996
rect 501696 142944 501748 142996
rect 483664 142876 483716 142928
rect 533988 142876 534040 142928
rect 450912 142808 450964 142860
rect 509608 142808 509660 142860
rect 362592 142128 362644 142180
rect 365536 142128 365588 142180
rect 479524 142128 479576 142180
rect 481916 142128 481968 142180
rect 533988 142128 534040 142180
rect 539876 142128 539928 142180
rect 452568 141924 452620 141976
rect 458916 141924 458968 141976
rect 462964 140768 463016 140820
rect 481916 140768 481968 140820
rect 452568 140632 452620 140684
rect 456248 140632 456300 140684
rect 534724 140020 534776 140072
rect 543188 140020 543240 140072
rect 361764 139340 361816 139392
rect 407764 139340 407816 139392
rect 451556 139340 451608 139392
rect 457444 139340 457496 139392
rect 554044 139340 554096 139392
rect 580172 139340 580224 139392
rect 538864 138524 538916 138576
rect 543096 138524 543148 138576
rect 452568 137844 452620 137896
rect 459192 137844 459244 137896
rect 452568 136484 452620 136536
rect 456156 136484 456208 136536
rect 452568 135124 452620 135176
rect 457536 135124 457588 135176
rect 452568 133764 452620 133816
rect 457628 133764 457680 133816
rect 452200 132404 452252 132456
rect 453304 132404 453356 132456
rect 359740 131112 359792 131164
rect 362592 131112 362644 131164
rect 452384 131044 452436 131096
rect 453396 131044 453448 131096
rect 390560 129752 390612 129804
rect 393964 129752 394016 129804
rect 361764 128256 361816 128308
rect 410616 128256 410668 128308
rect 361396 127576 361448 127628
rect 390560 127576 390612 127628
rect 452384 126896 452436 126948
rect 453488 126896 453540 126948
rect 576124 126896 576176 126948
rect 580172 126896 580224 126948
rect 365536 126216 365588 126268
rect 387064 126216 387116 126268
rect 451924 123360 451976 123412
rect 454960 123360 455012 123412
rect 451924 122136 451976 122188
rect 458824 122136 458876 122188
rect 359832 119076 359884 119128
rect 365536 119076 365588 119128
rect 361764 117240 361816 117292
rect 403624 117240 403676 117292
rect 569224 113092 569276 113144
rect 579804 113092 579856 113144
rect 451188 107380 451240 107432
rect 454868 107380 454920 107432
rect 439136 107244 439188 107296
rect 450636 107244 450688 107296
rect 432972 107176 433024 107228
rect 456064 107176 456116 107228
rect 426808 107108 426860 107160
rect 450820 107108 450872 107160
rect 420644 107040 420696 107092
rect 450728 107040 450780 107092
rect 389824 106972 389876 107024
rect 406384 106972 406436 107024
rect 414480 106972 414532 107024
rect 454776 106972 454828 107024
rect 402152 106904 402204 106956
rect 454684 106904 454736 106956
rect 445300 106496 445352 106548
rect 450544 106496 450596 106548
rect 361764 106224 361816 106276
rect 410524 106224 410576 106276
rect 566464 100648 566516 100700
rect 580172 100648 580224 100700
rect 3700 98608 3752 98660
rect 20904 98608 20956 98660
rect 361764 95140 361816 95192
rect 381360 95140 381412 95192
rect 3148 84192 3200 84244
rect 20904 84192 20956 84244
rect 361672 84124 361724 84176
rect 364064 84124 364116 84176
rect 361764 73108 361816 73160
rect 383476 73108 383528 73160
rect 544384 73108 544436 73160
rect 580172 73108 580224 73160
rect 3148 70388 3200 70440
rect 19984 70388 20036 70440
rect 4988 68960 5040 69012
rect 8208 68960 8260 69012
rect 4896 66172 4948 66224
rect 5540 66172 5592 66224
rect 5540 64132 5592 64184
rect 10968 64132 11020 64184
rect 361764 62024 361816 62076
rect 385592 62024 385644 62076
rect 8300 60868 8352 60920
rect 10324 60868 10376 60920
rect 5080 60664 5132 60716
rect 9496 60664 9548 60716
rect 547144 60664 547196 60716
rect 580172 60664 580224 60716
rect 11060 59372 11112 59424
rect 13820 59304 13872 59356
rect 9496 59100 9548 59152
rect 11060 59100 11112 59152
rect 3148 57944 3200 57996
rect 20076 57944 20128 57996
rect 11060 57876 11112 57928
rect 13728 57876 13780 57928
rect 4804 57128 4856 57180
rect 7380 57128 7432 57180
rect 13820 56516 13872 56568
rect 16488 56516 16540 56568
rect 7380 56108 7432 56160
rect 10508 56108 10560 56160
rect 5172 54612 5224 54664
rect 8208 54612 8260 54664
rect 13728 54340 13780 54392
rect 15200 54340 15252 54392
rect 10508 53796 10560 53848
rect 17500 53728 17552 53780
rect 16488 53456 16540 53508
rect 18880 53456 18932 53508
rect 361764 51076 361816 51128
rect 385592 51076 385644 51128
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 8208 51008 8260 51060
rect 11704 51008 11756 51060
rect 10324 49716 10376 49768
rect 15292 49648 15344 49700
rect 11704 48968 11756 49020
rect 20628 48968 20680 49020
rect 17500 48288 17552 48340
rect 20720 48220 20772 48272
rect 15292 46996 15344 47048
rect 21272 46996 21324 47048
rect 3700 46860 3752 46912
rect 386052 46860 386104 46912
rect 573364 46860 573416 46912
rect 580172 46860 580224 46912
rect 3240 46792 3292 46844
rect 384488 46792 384540 46844
rect 3332 46724 3384 46776
rect 384304 46724 384356 46776
rect 3976 46656 4028 46708
rect 381728 46656 381780 46708
rect 4068 46588 4120 46640
rect 381544 46588 381596 46640
rect 3608 46520 3660 46572
rect 379428 46520 379480 46572
rect 3792 46452 3844 46504
rect 379336 46452 379388 46504
rect 3516 46384 3568 46436
rect 378692 46384 378744 46436
rect 3424 46316 3476 46368
rect 375932 46316 375984 46368
rect 19984 46248 20036 46300
rect 384396 46248 384448 46300
rect 21456 46180 21508 46232
rect 384672 46180 384724 46232
rect 21272 46112 21324 46164
rect 361396 46112 361448 46164
rect 20812 46044 20864 46096
rect 359740 46044 359792 46096
rect 358268 45636 358320 45688
rect 361304 45636 361356 45688
rect 3884 45500 3936 45552
rect 382096 45500 382148 45552
rect 3424 45432 3476 45484
rect 368204 45432 368256 45484
rect 21364 45364 21416 45416
rect 376668 45364 376720 45416
rect 20720 45296 20772 45348
rect 358268 45296 358320 45348
rect 69020 45228 69072 45280
rect 376300 45228 376352 45280
rect 64880 45160 64932 45212
rect 376392 45160 376444 45212
rect 60740 45092 60792 45144
rect 379152 45092 379204 45144
rect 57980 45024 58032 45076
rect 378968 45024 379020 45076
rect 53840 44956 53892 45008
rect 379060 44956 379112 45008
rect 51080 44888 51132 44940
rect 379244 44888 379296 44940
rect 46940 44820 46992 44872
rect 381452 44820 381504 44872
rect 71780 44752 71832 44804
rect 376208 44752 376260 44804
rect 75920 44684 75972 44736
rect 376484 44684 376536 44736
rect 78680 44616 78732 44668
rect 373632 44616 373684 44668
rect 114560 42712 114612 42764
rect 367836 42712 367888 42764
rect 110420 42644 110472 42696
rect 367928 42644 367980 42696
rect 107660 42576 107712 42628
rect 368020 42576 368072 42628
rect 103520 42508 103572 42560
rect 367744 42508 367796 42560
rect 100760 42440 100812 42492
rect 370688 42440 370740 42492
rect 96620 42372 96672 42424
rect 371056 42372 371108 42424
rect 93860 42304 93912 42356
rect 370872 42304 370924 42356
rect 89720 42236 89772 42288
rect 370780 42236 370832 42288
rect 85580 42168 85632 42220
rect 370964 42168 371016 42220
rect 82820 42100 82872 42152
rect 373448 42100 373500 42152
rect 11060 42032 11112 42084
rect 373540 42032 373592 42084
rect 118700 41964 118752 42016
rect 365076 41964 365128 42016
rect 461584 41352 461636 41404
rect 536840 41352 536892 41404
rect 66260 39992 66312 40044
rect 365444 39992 365496 40044
rect 62120 39924 62172 39976
rect 366732 39924 366784 39976
rect 59360 39856 59412 39908
rect 368112 39856 368164 39908
rect 55220 39788 55272 39840
rect 366548 39788 366600 39840
rect 52460 39720 52512 39772
rect 363788 39720 363840 39772
rect 33140 39652 33192 39704
rect 363696 39652 363748 39704
rect 29000 39584 29052 39636
rect 362408 39584 362460 39636
rect 26240 39516 26292 39568
rect 362500 39516 362552 39568
rect 20720 39448 20772 39500
rect 365168 39448 365220 39500
rect 40040 39380 40092 39432
rect 384856 39380 384908 39432
rect 2780 39312 2832 39364
rect 365352 39312 365404 39364
rect 121460 39244 121512 39296
rect 365260 39244 365312 39296
rect 109040 37204 109092 37256
rect 377680 37204 377732 37256
rect 104900 37136 104952 37188
rect 375104 37136 375156 37188
rect 102140 37068 102192 37120
rect 376576 37068 376628 37120
rect 98000 37000 98052 37052
rect 374828 37000 374880 37052
rect 93952 36932 94004 36984
rect 374736 36932 374788 36984
rect 91100 36864 91152 36916
rect 375012 36864 375064 36916
rect 86960 36796 87012 36848
rect 372252 36796 372304 36848
rect 84200 36728 84252 36780
rect 373356 36728 373408 36780
rect 80060 36660 80112 36712
rect 369308 36660 369360 36712
rect 73160 36592 73212 36644
rect 369216 36592 369268 36644
rect 69112 36524 69164 36576
rect 366456 36524 366508 36576
rect 111800 36456 111852 36508
rect 378600 36456 378652 36508
rect 118792 34416 118844 34468
rect 380256 34416 380308 34468
rect 115940 34348 115992 34400
rect 377588 34348 377640 34400
rect 56600 34280 56652 34332
rect 369400 34280 369452 34332
rect 49700 34212 49752 34264
rect 366640 34212 366692 34264
rect 44180 34144 44232 34196
rect 363880 34144 363932 34196
rect 41420 34076 41472 34128
rect 361212 34076 361264 34128
rect 34520 34008 34572 34060
rect 382004 34008 382056 34060
rect 9680 33940 9732 33992
rect 363972 33940 364024 33992
rect 30380 33872 30432 33924
rect 386328 33872 386380 33924
rect 22100 33804 22152 33856
rect 383292 33804 383344 33856
rect 17960 33736 18012 33788
rect 380532 33736 380584 33788
rect 122840 33668 122892 33720
rect 382924 33668 382976 33720
rect 3516 33056 3568 33108
rect 378784 33056 378836 33108
rect 565084 33056 565136 33108
rect 580172 33056 580224 33108
rect 113180 31696 113232 31748
rect 372344 31696 372396 31748
rect 385592 31696 385644 31748
rect 462320 31696 462372 31748
rect 106280 31628 106332 31680
rect 369124 31628 369176 31680
rect 99380 31560 99432 31612
rect 366364 31560 366416 31612
rect 88340 31492 88392 31544
rect 385868 31492 385920 31544
rect 74540 31424 74592 31476
rect 383200 31424 383252 31476
rect 77300 31356 77352 31408
rect 386236 31356 386288 31408
rect 67640 31288 67692 31340
rect 377496 31288 377548 31340
rect 70400 31220 70452 31272
rect 380440 31220 380492 31272
rect 60832 31152 60884 31204
rect 372068 31152 372120 31204
rect 63500 31084 63552 31136
rect 374920 31084 374972 31136
rect 13820 31016 13872 31068
rect 384764 31016 384816 31068
rect 124220 30948 124272 31000
rect 380164 30948 380216 31000
rect 92480 29588 92532 29640
rect 460204 29588 460256 29640
rect 117320 28636 117372 28688
rect 374644 28636 374696 28688
rect 42800 28568 42852 28620
rect 373264 28568 373316 28620
rect 38660 28500 38712 28552
rect 376116 28500 376168 28552
rect 35900 28432 35952 28484
rect 378876 28432 378928 28484
rect 31760 28364 31812 28416
rect 381912 28364 381964 28416
rect 19340 28296 19392 28348
rect 377404 28296 377456 28348
rect 27620 28228 27672 28280
rect 386144 28228 386196 28280
rect 3424 20612 3476 20664
rect 383384 20612 383436 20664
rect 562324 20612 562376 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 376024 6808 376076 6860
rect 563704 6808 563756 6860
rect 580172 6808 580224 6860
rect 85672 4088 85724 4140
rect 360936 4088 360988 4140
rect 96252 4020 96304 4072
rect 371884 4020 371936 4072
rect 82084 3952 82136 4004
rect 359464 3952 359516 4004
rect 77392 3884 77444 3936
rect 370596 3884 370648 3936
rect 53748 3816 53800 3868
rect 359556 3816 359608 3868
rect 48964 3748 49016 3800
rect 364984 3748 365036 3800
rect 46664 3680 46716 3732
rect 363604 3680 363656 3732
rect 38384 3612 38436 3664
rect 362316 3612 362368 3664
rect 27712 3544 27764 3596
rect 385776 3544 385828 3596
rect 24216 3476 24268 3528
rect 383108 3476 383160 3528
rect 17040 3408 17092 3460
rect 380348 3408 380400 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 103336 3340 103388 3392
rect 361120 3340 361172 3392
rect 110420 3272 110472 3324
rect 111616 3272 111668 3324
rect 110512 3204 110564 3256
rect 360844 3272 360896 3324
rect 121092 3204 121144 3256
rect 361028 3204 361080 3256
rect 44272 2184 44324 2236
rect 385684 2184 385736 2236
rect 37188 2116 37240 2168
rect 383016 2116 383068 2168
rect 2872 2048 2924 2100
rect 381636 2048 381688 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 23492 687857 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 23478 687848 23534 687857
rect 23478 687783 23534 687792
rect 88352 685137 88380 702406
rect 105464 700534 105492 703520
rect 137848 700602 137876 703520
rect 154132 700670 154160 703520
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 170324 700369 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170310 700360 170366 700369
rect 170310 700295 170366 700304
rect 201512 686526 201540 702986
rect 218072 686594 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700738 235212 703520
rect 235172 700732 235224 700738
rect 235172 700674 235224 700680
rect 267660 697610 267688 703520
rect 283852 700806 283880 703520
rect 283840 700800 283892 700806
rect 283840 700742 283892 700748
rect 300136 700505 300164 703520
rect 332520 700641 332548 703520
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 332506 700632 332562 700641
rect 332506 700567 332562 700576
rect 300122 700496 300178 700505
rect 300122 700431 300178 700440
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 218060 686588 218112 686594
rect 218060 686530 218112 686536
rect 201500 686520 201552 686526
rect 201500 686462 201552 686468
rect 266372 685166 266400 697546
rect 347792 685234 347820 702406
rect 364996 700874 365024 703520
rect 397472 700942 397500 703520
rect 397460 700936 397512 700942
rect 397460 700878 397512 700884
rect 364984 700868 365036 700874
rect 364984 700810 365036 700816
rect 347780 685228 347832 685234
rect 347780 685170 347832 685176
rect 266360 685160 266412 685166
rect 88338 685128 88394 685137
rect 266360 685102 266412 685108
rect 88338 685063 88394 685072
rect 19984 684820 20036 684826
rect 19984 684762 20036 684768
rect 3608 684752 3660 684758
rect 3608 684694 3660 684700
rect 3332 684684 3384 684690
rect 3332 684626 3384 684632
rect 3148 684616 3200 684622
rect 3148 684558 3200 684564
rect 2964 682780 3016 682786
rect 2964 682722 3016 682728
rect 2872 682712 2924 682718
rect 2872 682654 2924 682660
rect 2884 673454 2912 682654
rect 2976 677770 3004 682722
rect 3160 677906 3188 684558
rect 3344 683114 3372 684626
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3516 683392 3568 683398
rect 3516 683334 3568 683340
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3344 683086 3464 683114
rect 3436 678450 3464 683086
rect 3528 678570 3556 683334
rect 3620 678570 3648 684694
rect 3884 684548 3936 684554
rect 3884 684490 3936 684496
rect 3700 683324 3752 683330
rect 3700 683266 3752 683272
rect 3516 678564 3568 678570
rect 3516 678506 3568 678512
rect 3608 678564 3660 678570
rect 3608 678506 3660 678512
rect 3436 678422 3648 678450
rect 3516 678360 3568 678366
rect 3516 678302 3568 678308
rect 3160 677878 3464 677906
rect 2976 677742 3372 677770
rect 2884 673426 3280 673454
rect 3148 658232 3200 658238
rect 3146 658200 3148 658209
rect 3200 658200 3202 658209
rect 3146 658135 3202 658144
rect 3252 580009 3280 673426
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 677742
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 449585 3464 677878
rect 3528 462641 3556 678302
rect 3620 475697 3648 678422
rect 3712 632097 3740 683266
rect 3896 678314 3924 684490
rect 17960 683596 18012 683602
rect 17960 683538 18012 683544
rect 4068 683460 4120 683466
rect 4068 683402 4120 683408
rect 3976 683188 4028 683194
rect 3976 683130 4028 683136
rect 3804 678286 3924 678314
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3700 631372 3752 631378
rect 3700 631314 3752 631320
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3712 423609 3740 631314
rect 3804 501809 3832 678286
rect 3884 678224 3936 678230
rect 3884 678166 3936 678172
rect 3896 514865 3924 678166
rect 3988 527921 4016 683130
rect 4080 553897 4108 683402
rect 17972 683114 18000 683538
rect 17880 683086 18000 683114
rect 17880 680406 17908 683086
rect 17868 680400 17920 680406
rect 17868 680342 17920 680348
rect 12900 680332 12952 680338
rect 12900 680274 12952 680280
rect 12912 676258 12940 680274
rect 12900 676252 12952 676258
rect 12900 676194 12952 676200
rect 10416 676184 10468 676190
rect 10416 676126 10468 676132
rect 10428 667962 10456 676126
rect 8024 667956 8076 667962
rect 8024 667898 8076 667904
rect 10416 667956 10468 667962
rect 10416 667898 10468 667904
rect 8036 665242 8064 667898
rect 4804 665236 4856 665242
rect 4804 665178 4856 665184
rect 8024 665236 8076 665242
rect 8024 665178 8076 665184
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 665178
rect 19996 658238 20024 684762
rect 359464 683596 359516 683602
rect 359464 683538 359516 683544
rect 21364 683528 21416 683534
rect 21364 683470 21416 683476
rect 19984 658232 20036 658238
rect 19984 658174 20036 658180
rect 21376 634814 21404 683470
rect 20916 634786 21404 634814
rect 20916 631378 20944 634786
rect 20904 631372 20956 631378
rect 20904 631314 20956 631320
rect 359476 601730 359504 683538
rect 361764 679040 361816 679046
rect 361762 679008 361764 679017
rect 364984 679040 365036 679046
rect 361816 679008 361818 679017
rect 364984 678982 365036 678988
rect 361762 678943 361818 678952
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 361764 667898 361816 667904
rect 361670 656976 361726 656985
rect 361670 656911 361726 656920
rect 361684 656198 361712 656911
rect 361672 656192 361724 656198
rect 361672 656134 361724 656140
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 361764 645866 361816 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 361578 612912 361634 612921
rect 361578 612847 361634 612856
rect 361592 612814 361620 612847
rect 361580 612808 361632 612814
rect 361580 612750 361632 612756
rect 361762 601896 361818 601905
rect 361762 601831 361818 601840
rect 361776 601730 361804 601831
rect 359464 601724 359516 601730
rect 359464 601666 359516 601672
rect 361764 601724 361816 601730
rect 361764 601666 361816 601672
rect 361762 590880 361818 590889
rect 361762 590815 361818 590824
rect 361776 590714 361804 590815
rect 361764 590708 361816 590714
rect 361764 590650 361816 590656
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 361762 568848 361818 568857
rect 361762 568783 361818 568792
rect 361776 568614 361804 568783
rect 361764 568608 361816 568614
rect 361764 568550 361816 568556
rect 361578 557832 361634 557841
rect 361578 557767 361580 557776
rect 361632 557767 361634 557776
rect 363604 557796 363656 557802
rect 361580 557738 361632 557744
rect 363604 557738 363656 557744
rect 361578 546816 361634 546825
rect 361578 546751 361634 546760
rect 361592 546650 361620 546751
rect 361580 546644 361632 546650
rect 361580 546586 361632 546592
rect 361578 535800 361634 535809
rect 361578 535735 361580 535744
rect 361632 535735 361634 535744
rect 361580 535706 361632 535712
rect 361762 524784 361818 524793
rect 361762 524719 361818 524728
rect 361776 524482 361804 524719
rect 361764 524476 361816 524482
rect 361764 524418 361816 524424
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 423600 3754 423609
rect 3698 423535 3754 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 361762 491736 361818 491745
rect 361762 491671 361818 491680
rect 361776 491366 361804 491671
rect 361764 491360 361816 491366
rect 361764 491302 361816 491308
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 362222 469704 362278 469713
rect 362222 469639 362278 469648
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 361762 436656 361818 436665
rect 361762 436591 361818 436600
rect 361776 436150 361804 436591
rect 361764 436144 361816 436150
rect 361764 436086 361816 436092
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 362236 413302 362264 469639
rect 362314 447672 362370 447681
rect 362314 447607 362370 447616
rect 362328 416090 362356 447607
rect 362406 425640 362462 425649
rect 362406 425575 362462 425584
rect 362420 418810 362448 425575
rect 362408 418804 362460 418810
rect 362408 418746 362460 418752
rect 362316 416084 362368 416090
rect 362316 416026 362368 416032
rect 362224 413296 362276 413302
rect 362224 413238 362276 413244
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3882 397488 3938 397497
rect 3882 397423 3938 397432
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 305046 3464 358391
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3528 301986 3556 345335
rect 3606 319288 3662 319297
rect 3606 319223 3662 319232
rect 3516 301980 3568 301986
rect 3516 301922 3568 301928
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3238 149832 3294 149841
rect 3238 149767 3294 149776
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3146 71632 3202 71641
rect 3146 71567 3202 71576
rect 3160 70446 3188 71567
rect 3148 70440 3200 70446
rect 3148 70382 3200 70388
rect 3146 58576 3202 58585
rect 3146 58511 3202 58520
rect 3160 58002 3188 58511
rect 3148 57996 3200 58002
rect 3148 57938 3200 57944
rect 3252 46850 3280 149767
rect 3240 46844 3292 46850
rect 3240 46786 3292 46792
rect 3344 46782 3372 162823
rect 3332 46776 3384 46782
rect 3332 46718 3384 46724
rect 3436 46374 3464 293111
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3528 46442 3556 267135
rect 3620 259418 3648 319223
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3608 259412 3660 259418
rect 3608 259354 3660 259360
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3620 46578 3648 254079
rect 3712 98666 3740 306167
rect 3896 241466 3924 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 363616 376650 363644 557738
rect 363696 546644 363748 546650
rect 363696 546586 363748 546592
rect 363708 376718 363736 546586
rect 363788 535764 363840 535770
rect 363788 535706 363840 535712
rect 363696 376712 363748 376718
rect 363696 376654 363748 376660
rect 363604 376644 363656 376650
rect 363604 376586 363656 376592
rect 363800 375358 363828 535706
rect 364996 385014 365024 678982
rect 381544 667956 381596 667962
rect 381544 667898 381596 667904
rect 378784 645924 378836 645930
rect 378784 645866 378836 645872
rect 376024 623824 376076 623830
rect 376024 623766 376076 623772
rect 374736 601724 374788 601730
rect 374736 601666 374788 601672
rect 366364 601656 366416 601662
rect 366364 601598 366416 601604
rect 366376 590646 366404 601598
rect 371884 590708 371936 590714
rect 371884 590650 371936 590656
rect 366364 590640 366416 590646
rect 366364 590582 366416 590588
rect 367560 590640 367612 590646
rect 367560 590582 367612 590588
rect 367572 586566 367600 590582
rect 367560 586560 367612 586566
rect 367560 586502 367612 586508
rect 370504 579692 370556 579698
rect 370504 579634 370556 579640
rect 367744 568608 367796 568614
rect 367744 568550 367796 568556
rect 364984 385008 365036 385014
rect 364984 384950 365036 384956
rect 367756 378146 367784 568550
rect 367744 378140 367796 378146
rect 367744 378082 367796 378088
rect 370516 378078 370544 579634
rect 371896 379506 371924 590650
rect 372528 586492 372580 586498
rect 372528 586434 372580 586440
rect 372540 580938 372568 586434
rect 372540 580910 372660 580938
rect 372632 577454 372660 580910
rect 372620 577448 372672 577454
rect 372620 577390 372672 577396
rect 374644 385076 374696 385082
rect 374644 385018 374696 385024
rect 371884 379500 371936 379506
rect 371884 379442 371936 379448
rect 370504 378072 370556 378078
rect 370504 378014 370556 378020
rect 363788 375352 363840 375358
rect 363788 375294 363840 375300
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3884 241460 3936 241466
rect 3884 241402 3936 241408
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3700 98660 3752 98666
rect 3700 98602 3752 98608
rect 3698 97608 3754 97617
rect 3698 97543 3754 97552
rect 3712 46918 3740 97543
rect 3700 46912 3752 46918
rect 3700 46854 3752 46860
rect 3608 46572 3660 46578
rect 3608 46514 3660 46520
rect 3804 46510 3832 241023
rect 3988 218074 4016 371311
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 362222 359544 362278 359553
rect 362222 359479 362278 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362236 347750 362264 359479
rect 362224 347744 362276 347750
rect 362224 347686 362276 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 336048 362276 336054
rect 362224 335990 362276 335996
rect 362236 326505 362264 335990
rect 364064 334008 364116 334014
rect 364064 333950 364116 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 363602 305824 363658 305833
rect 363602 305759 363658 305768
rect 360844 305720 360896 305726
rect 360844 305662 360896 305668
rect 4804 305040 4856 305046
rect 4804 304982 4856 304988
rect 3976 218068 4028 218074
rect 3976 218010 4028 218016
rect 3882 214976 3938 214985
rect 3882 214911 3938 214920
rect 3792 46504 3844 46510
rect 3792 46446 3844 46452
rect 3516 46436 3568 46442
rect 3516 46378 3568 46384
rect 3424 46368 3476 46374
rect 3424 46310 3476 46316
rect 3896 45558 3924 214911
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3988 46714 4016 201855
rect 4066 188864 4122 188873
rect 4066 188799 4122 188808
rect 3976 46708 4028 46714
rect 3976 46650 4028 46656
rect 4080 46646 4108 188799
rect 4816 57186 4844 304982
rect 4896 301980 4948 301986
rect 4896 301922 4948 301928
rect 4908 66230 4936 301922
rect 359464 276684 359516 276690
rect 359464 276626 359516 276632
rect 4988 259412 5040 259418
rect 4988 259354 5040 259360
rect 5000 69018 5028 259354
rect 5080 241460 5132 241466
rect 5080 241402 5132 241408
rect 4988 69012 5040 69018
rect 4988 68954 5040 68960
rect 4896 66224 4948 66230
rect 4896 66166 4948 66172
rect 5092 60722 5120 241402
rect 5172 218068 5224 218074
rect 5172 218010 5224 218016
rect 5080 60716 5132 60722
rect 5080 60658 5132 60664
rect 4804 57180 4856 57186
rect 4804 57122 4856 57128
rect 5184 54670 5212 218010
rect 20904 98660 20956 98666
rect 20904 98602 20956 98608
rect 20916 93854 20944 98602
rect 20916 93826 21404 93854
rect 20904 84244 20956 84250
rect 20904 84186 20956 84192
rect 20916 73681 20944 84186
rect 21376 77294 21404 93826
rect 21284 77266 21404 77294
rect 20902 73672 20958 73681
rect 20902 73607 20958 73616
rect 19984 70440 20036 70446
rect 19984 70382 20036 70388
rect 8208 69012 8260 69018
rect 8208 68954 8260 68960
rect 5540 66224 5592 66230
rect 5540 66166 5592 66172
rect 5552 64190 5580 66166
rect 8220 64874 8248 68954
rect 8220 64846 8340 64874
rect 5540 64184 5592 64190
rect 5540 64126 5592 64132
rect 8312 60926 8340 64846
rect 10968 64184 11020 64190
rect 10968 64126 11020 64132
rect 10980 63458 11008 64126
rect 10980 63430 11100 63458
rect 8300 60920 8352 60926
rect 8300 60862 8352 60868
rect 10324 60920 10376 60926
rect 10324 60862 10376 60868
rect 9496 60716 9548 60722
rect 9496 60658 9548 60664
rect 9508 59158 9536 60658
rect 9496 59152 9548 59158
rect 9496 59094 9548 59100
rect 7380 57180 7432 57186
rect 7380 57122 7432 57128
rect 7392 56166 7420 57122
rect 7380 56160 7432 56166
rect 7380 56102 7432 56108
rect 5172 54664 5224 54670
rect 5172 54606 5224 54612
rect 8208 54664 8260 54670
rect 8208 54606 8260 54612
rect 8220 51066 8248 54606
rect 8208 51060 8260 51066
rect 8208 51002 8260 51008
rect 10336 49774 10364 60862
rect 11072 59430 11100 63430
rect 11060 59424 11112 59430
rect 11060 59366 11112 59372
rect 13820 59356 13872 59362
rect 13820 59298 13872 59304
rect 11060 59152 11112 59158
rect 11060 59094 11112 59100
rect 11072 57934 11100 59094
rect 11060 57928 11112 57934
rect 11060 57870 11112 57876
rect 13728 57928 13780 57934
rect 13728 57870 13780 57876
rect 10508 56160 10560 56166
rect 10508 56102 10560 56108
rect 10520 53854 10548 56102
rect 13740 54398 13768 57870
rect 13832 56574 13860 59298
rect 13820 56568 13872 56574
rect 13820 56510 13872 56516
rect 16488 56568 16540 56574
rect 16488 56510 16540 56516
rect 13728 54392 13780 54398
rect 13728 54334 13780 54340
rect 15200 54392 15252 54398
rect 15200 54334 15252 54340
rect 10508 53848 10560 53854
rect 10508 53790 10560 53796
rect 11704 51060 11756 51066
rect 11704 51002 11756 51008
rect 10324 49768 10376 49774
rect 10324 49710 10376 49716
rect 11716 49026 11744 51002
rect 11704 49020 11756 49026
rect 11704 48962 11756 48968
rect 15212 48929 15240 54334
rect 16500 53514 16528 56510
rect 17500 53780 17552 53786
rect 17500 53722 17552 53728
rect 16488 53508 16540 53514
rect 16488 53450 16540 53456
rect 15292 49700 15344 49706
rect 15292 49642 15344 49648
rect 15198 48920 15254 48929
rect 15198 48855 15254 48864
rect 15304 47054 15332 49642
rect 17512 48346 17540 53722
rect 18880 53508 18932 53514
rect 18880 53450 18932 53456
rect 18892 49609 18920 53450
rect 18878 49600 18934 49609
rect 18878 49535 18934 49544
rect 17500 48340 17552 48346
rect 17500 48282 17552 48288
rect 15292 47048 15344 47054
rect 15292 46990 15344 46996
rect 4068 46640 4120 46646
rect 4068 46582 4120 46588
rect 19996 46306 20024 70382
rect 21284 67634 21312 77266
rect 21454 73672 21510 73681
rect 21454 73607 21510 73616
rect 21284 67606 21404 67634
rect 20076 57996 20128 58002
rect 20076 57938 20128 57944
rect 20088 46753 20116 57938
rect 20628 49020 20680 49026
rect 20628 48962 20680 48968
rect 20640 48362 20668 48962
rect 20640 48334 20852 48362
rect 20720 48272 20772 48278
rect 20720 48214 20772 48220
rect 20074 46744 20130 46753
rect 20074 46679 20130 46688
rect 19984 46300 20036 46306
rect 19984 46242 20036 46248
rect 3884 45552 3936 45558
rect 3422 45520 3478 45529
rect 3884 45494 3936 45500
rect 3422 45455 3424 45464
rect 3476 45455 3478 45464
rect 3424 45426 3476 45432
rect 20732 45354 20760 48214
rect 20824 46102 20852 48334
rect 21272 47048 21324 47054
rect 21272 46990 21324 46996
rect 21284 46170 21312 46990
rect 21272 46164 21324 46170
rect 21272 46106 21324 46112
rect 20812 46096 20864 46102
rect 20812 46038 20864 46044
rect 21376 45422 21404 67606
rect 21468 46238 21496 73607
rect 21456 46232 21508 46238
rect 21456 46174 21508 46180
rect 358268 45688 358320 45694
rect 358268 45630 358320 45636
rect 21364 45416 21416 45422
rect 21364 45358 21416 45364
rect 358280 45354 358308 45630
rect 20720 45348 20772 45354
rect 20720 45290 20772 45296
rect 358268 45348 358320 45354
rect 358268 45290 358320 45296
rect 69020 45280 69072 45286
rect 69020 45222 69072 45228
rect 64880 45212 64932 45218
rect 64880 45154 64932 45160
rect 60740 45144 60792 45150
rect 60740 45086 60792 45092
rect 57980 45076 58032 45082
rect 57980 45018 58032 45024
rect 53840 45008 53892 45014
rect 53840 44950 53892 44956
rect 51080 44940 51132 44946
rect 51080 44882 51132 44888
rect 46940 44872 46992 44878
rect 6918 44840 6974 44849
rect 46940 44814 46992 44820
rect 6918 44775 6974 44784
rect 2780 39364 2832 39370
rect 2780 39306 2832 39312
rect 2792 16574 2820 39306
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 6932 16574 6960 44775
rect 11060 42084 11112 42090
rect 11060 42026 11112 42032
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 2792 16546 3648 16574
rect 6932 16546 7696 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2884 480 2912 2042
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5262 4040 5318 4049
rect 5262 3975 5318 3984
rect 5276 480 5304 3975
rect 6458 3632 6514 3641
rect 6458 3567 6514 3576
rect 6472 480 6500 3567
rect 7668 480 7696 16546
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8772 480 8800 3703
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 33934
rect 11072 16574 11100 42026
rect 33140 39704 33192 39710
rect 33140 39646 33192 39652
rect 29000 39636 29052 39642
rect 29000 39578 29052 39584
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 20720 39500 20772 39506
rect 20720 39442 20772 39448
rect 17960 33788 18012 33794
rect 17960 33730 18012 33736
rect 13820 31068 13872 31074
rect 13820 31010 13872 31016
rect 13832 16574 13860 31010
rect 11072 16546 11928 16574
rect 13832 16546 14320 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13556 480 13584 3839
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 480 17080 3402
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 33730
rect 19340 28348 19392 28354
rect 19340 28290 19392 28296
rect 19352 16574 19380 28290
rect 20732 16574 20760 39442
rect 22100 33856 22152 33862
rect 22100 33798 22152 33804
rect 22112 16574 22140 33798
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19444 480 19472 16546
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 39510
rect 27620 28280 27672 28286
rect 27620 28222 27672 28228
rect 27632 16574 27660 28222
rect 29012 16574 29040 39578
rect 30380 33924 30432 33930
rect 30380 33866 30432 33872
rect 30392 16574 30420 33866
rect 31760 28416 31812 28422
rect 31760 28358 31812 28364
rect 31772 16574 31800 28358
rect 33152 16574 33180 39646
rect 40040 39432 40092 39438
rect 40040 39374 40092 39380
rect 34520 34060 34572 34066
rect 34520 34002 34572 34008
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27724 480 27752 3538
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 34002
rect 38660 28552 38712 28558
rect 38660 28494 38712 28500
rect 35900 28484 35952 28490
rect 35900 28426 35952 28432
rect 35912 16574 35940 28426
rect 38672 16574 38700 28494
rect 40052 16574 40080 39374
rect 44180 34196 44232 34202
rect 44180 34138 44232 34144
rect 41420 34128 41472 34134
rect 41420 34070 41472 34076
rect 41432 16574 41460 34070
rect 42800 28620 42852 28626
rect 42800 28562 42852 28568
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 36004 480 36032 16546
rect 38384 3664 38436 3670
rect 38384 3606 38436 3612
rect 37188 2168 37240 2174
rect 37188 2110 37240 2116
rect 37200 480 37228 2110
rect 38396 480 38424 3606
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 28562
rect 44192 16574 44220 34138
rect 46952 16574 46980 44814
rect 49700 34264 49752 34270
rect 49700 34206 49752 34212
rect 49712 16574 49740 34206
rect 44192 16546 45048 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44272 2236 44324 2242
rect 44272 2178 44324 2184
rect 44284 480 44312 2178
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 46676 480 46704 3674
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 3800 49016 3806
rect 48964 3742 49016 3748
rect 48976 480 49004 3742
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 44882
rect 52460 39772 52512 39778
rect 52460 39714 52512 39720
rect 52472 16574 52500 39714
rect 53852 16574 53880 44950
rect 55220 39840 55272 39846
rect 55220 39782 55272 39788
rect 55232 16574 55260 39782
rect 56600 34332 56652 34338
rect 56600 34274 56652 34280
rect 56612 16574 56640 34274
rect 57992 16574 58020 45018
rect 59360 39908 59412 39914
rect 59360 39850 59412 39856
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52564 480 52592 16546
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 53760 480 53788 3810
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 39850
rect 60752 3398 60780 45086
rect 62120 39976 62172 39982
rect 62120 39918 62172 39924
rect 60832 31204 60884 31210
rect 60832 31146 60884 31152
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 31146
rect 62132 16574 62160 39918
rect 63500 31136 63552 31142
rect 63500 31078 63552 31084
rect 63512 16574 63540 31078
rect 64892 16574 64920 45154
rect 66260 40044 66312 40050
rect 66260 39986 66312 39992
rect 66272 16574 66300 39986
rect 67640 31340 67692 31346
rect 67640 31282 67692 31288
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 31282
rect 69032 6914 69060 45222
rect 71780 44804 71832 44810
rect 71780 44746 71832 44752
rect 69112 36576 69164 36582
rect 69112 36518 69164 36524
rect 69124 16574 69152 36518
rect 70400 31272 70452 31278
rect 70400 31214 70452 31220
rect 70412 16574 70440 31214
rect 71792 16574 71820 44746
rect 75920 44736 75972 44742
rect 75920 44678 75972 44684
rect 73160 36644 73212 36650
rect 73160 36586 73212 36592
rect 73172 16574 73200 36586
rect 74540 31476 74592 31482
rect 74540 31418 74592 31424
rect 74552 16574 74580 31418
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 44678
rect 78680 44668 78732 44674
rect 78680 44610 78732 44616
rect 77300 31408 77352 31414
rect 77300 31350 77352 31356
rect 77312 16574 77340 31350
rect 78692 16574 78720 44610
rect 114560 42764 114612 42770
rect 114560 42706 114612 42712
rect 110420 42696 110472 42702
rect 110420 42638 110472 42644
rect 107660 42628 107712 42634
rect 107660 42570 107712 42576
rect 103520 42560 103572 42566
rect 103520 42502 103572 42508
rect 100760 42492 100812 42498
rect 100760 42434 100812 42440
rect 96620 42424 96672 42430
rect 96620 42366 96672 42372
rect 93860 42356 93912 42362
rect 93860 42298 93912 42304
rect 89720 42288 89772 42294
rect 89720 42230 89772 42236
rect 85580 42220 85632 42226
rect 85580 42162 85632 42168
rect 82820 42152 82872 42158
rect 82820 42094 82872 42100
rect 80060 36712 80112 36718
rect 80060 36654 80112 36660
rect 80072 16574 80100 36654
rect 82832 16574 82860 42094
rect 84200 36780 84252 36786
rect 84200 36722 84252 36728
rect 77312 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 82832 16546 83320 16574
rect 77392 3936 77444 3942
rect 77392 3878 77444 3884
rect 77404 480 77432 3878
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 82096 480 82124 3946
rect 83292 480 83320 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 36722
rect 85592 16574 85620 42162
rect 86960 36848 87012 36854
rect 86960 36790 87012 36796
rect 86972 16574 87000 36790
rect 88340 31544 88392 31550
rect 88340 31486 88392 31492
rect 88352 16574 88380 31486
rect 89732 16574 89760 42230
rect 91100 36916 91152 36922
rect 91100 36858 91152 36864
rect 91112 16574 91140 36858
rect 92480 29640 92532 29646
rect 92480 29582 92532 29588
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 85684 480 85712 4082
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 29582
rect 93872 6914 93900 42298
rect 93952 36984 94004 36990
rect 93952 36926 94004 36932
rect 93964 16574 93992 36926
rect 96632 16574 96660 42366
rect 98000 37052 98052 37058
rect 98000 36994 98052 37000
rect 98012 16574 98040 36994
rect 99380 31612 99432 31618
rect 99380 31554 99432 31560
rect 99392 16574 99420 31554
rect 93964 16546 94728 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96252 4072 96304 4078
rect 96252 4014 96304 4020
rect 96264 480 96292 4014
rect 97460 480 97488 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 42434
rect 102140 37120 102192 37126
rect 102140 37062 102192 37068
rect 102152 16574 102180 37062
rect 103532 16574 103560 42502
rect 104900 37188 104952 37194
rect 104900 37130 104952 37136
rect 104912 16574 104940 37130
rect 106280 31680 106332 31686
rect 106280 31622 106332 31628
rect 106292 16574 106320 31622
rect 107672 16574 107700 42570
rect 109040 37256 109092 37262
rect 109040 37198 109092 37204
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 37198
rect 110432 3330 110460 42638
rect 111800 36508 111852 36514
rect 111800 36450 111852 36456
rect 111812 16574 111840 36450
rect 113180 31748 113232 31754
rect 113180 31690 113232 31696
rect 113192 16574 113220 31690
rect 114572 16574 114600 42706
rect 118700 42016 118752 42022
rect 118700 41958 118752 41964
rect 115940 34400 115992 34406
rect 115940 34342 115992 34348
rect 115952 16574 115980 34342
rect 117320 28688 117372 28694
rect 117320 28630 117372 28636
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110420 3324 110472 3330
rect 110420 3266 110472 3272
rect 111616 3324 111668 3330
rect 111616 3266 111668 3272
rect 110512 3256 110564 3262
rect 110512 3198 110564 3204
rect 110524 480 110552 3198
rect 111628 480 111656 3266
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 28630
rect 118712 6914 118740 41958
rect 121460 39296 121512 39302
rect 121460 39238 121512 39244
rect 118792 34468 118844 34474
rect 118792 34410 118844 34416
rect 118804 16574 118832 34410
rect 121472 16574 121500 39238
rect 122840 33720 122892 33726
rect 122840 33662 122892 33668
rect 122852 16574 122880 33662
rect 124220 31000 124272 31006
rect 124220 30942 124272 30948
rect 124232 16574 124260 30942
rect 118804 16546 119936 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 121092 3256 121144 3262
rect 121092 3198 121144 3204
rect 121104 480 121132 3198
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 359476 4010 359504 276626
rect 359556 269816 359608 269822
rect 359556 269758 359608 269764
rect 359464 4004 359516 4010
rect 359464 3946 359516 3952
rect 359568 3874 359596 269758
rect 359648 163056 359700 163062
rect 359648 162998 359700 163004
rect 359660 46481 359688 162998
rect 359740 131164 359792 131170
rect 359740 131106 359792 131112
rect 359646 46472 359702 46481
rect 359646 46407 359702 46416
rect 359752 46102 359780 131106
rect 359832 119128 359884 119134
rect 359832 119070 359884 119076
rect 359844 46617 359872 119070
rect 359830 46608 359886 46617
rect 359830 46543 359886 46552
rect 359740 46096 359792 46102
rect 359740 46038 359792 46044
rect 359556 3868 359608 3874
rect 359556 3810 359608 3816
rect 360856 3330 360884 305662
rect 360936 305652 360988 305658
rect 360936 305594 360988 305600
rect 360948 4146 360976 305594
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 362224 304360 362276 304366
rect 362224 304302 362276 304308
rect 361028 304292 361080 304298
rect 361028 304234 361080 304240
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 360844 3324 360896 3330
rect 360844 3266 360896 3272
rect 361040 3262 361068 304234
rect 361120 302932 361172 302938
rect 361120 302874 361172 302880
rect 361132 3398 361160 302874
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361212 291848 361264 291854
rect 361212 291790 361264 291796
rect 361224 34134 361252 291790
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361672 216368 361724 216374
rect 361670 216336 361672 216345
rect 361724 216336 361726 216345
rect 361670 216271 361726 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361764 194540 361816 194546
rect 361764 194482 361816 194488
rect 361776 194313 361804 194482
rect 361762 194304 361818 194313
rect 361762 194239 361818 194248
rect 361764 183524 361816 183530
rect 361764 183466 361816 183472
rect 361776 183297 361804 183466
rect 361762 183288 361818 183297
rect 361762 183223 361818 183232
rect 361304 175976 361356 175982
rect 361304 175918 361356 175924
rect 361316 45694 361344 175918
rect 361762 172272 361818 172281
rect 361762 172207 361818 172216
rect 361776 171834 361804 172207
rect 361764 171828 361816 171834
rect 361764 171770 361816 171776
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361764 128308 361816 128314
rect 361764 128250 361816 128256
rect 361776 128217 361804 128250
rect 361762 128208 361818 128217
rect 361762 128143 361818 128152
rect 361396 127628 361448 127634
rect 361396 127570 361448 127576
rect 361408 46170 361436 127570
rect 361764 117292 361816 117298
rect 361764 117234 361816 117240
rect 361776 117201 361804 117234
rect 361762 117192 361818 117201
rect 361762 117127 361818 117136
rect 361764 106276 361816 106282
rect 361764 106218 361816 106224
rect 361776 106185 361804 106218
rect 361762 106176 361818 106185
rect 361762 106111 361818 106120
rect 361764 95192 361816 95198
rect 361762 95160 361764 95169
rect 361816 95160 361818 95169
rect 361762 95095 361818 95104
rect 361672 84176 361724 84182
rect 361670 84144 361672 84153
rect 361724 84144 361726 84153
rect 361670 84079 361726 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 51128 361816 51134
rect 361762 51096 361764 51105
rect 361816 51096 361818 51105
rect 361762 51031 361818 51040
rect 361396 46164 361448 46170
rect 361396 46106 361448 46112
rect 361304 45688 361356 45694
rect 361304 45630 361356 45636
rect 361212 34128 361264 34134
rect 361212 34070 361264 34076
rect 362236 4049 362264 304302
rect 362500 297764 362552 297770
rect 362500 297706 362552 297712
rect 362406 297664 362462 297673
rect 362406 297599 362462 297608
rect 362316 291916 362368 291922
rect 362316 291858 362368 291864
rect 362222 4040 362278 4049
rect 362222 3975 362278 3984
rect 362328 3670 362356 291858
rect 362420 39642 362448 297599
rect 362408 39636 362460 39642
rect 362408 39578 362460 39584
rect 362512 39574 362540 297706
rect 362592 291712 362644 291718
rect 362592 291654 362644 291660
rect 362604 271425 362632 291654
rect 362590 271416 362646 271425
rect 362590 271351 362646 271360
rect 362592 161492 362644 161498
rect 362592 161434 362644 161440
rect 362604 150249 362632 161434
rect 362590 150240 362646 150249
rect 362590 150175 362646 150184
rect 362592 142180 362644 142186
rect 362592 142122 362644 142128
rect 362604 131170 362632 142122
rect 362592 131164 362644 131170
rect 362592 131106 362644 131112
rect 362500 39568 362552 39574
rect 362500 39510 362552 39516
rect 363616 3738 363644 305759
rect 363696 297492 363748 297498
rect 363696 297434 363748 297440
rect 363708 39710 363736 297434
rect 363788 297424 363840 297430
rect 363788 297366 363840 297372
rect 363800 39778 363828 297366
rect 363972 289672 364024 289678
rect 363972 289614 364024 289620
rect 363880 289128 363932 289134
rect 363880 289070 363932 289076
rect 363788 39772 363840 39778
rect 363788 39714 363840 39720
rect 363696 39704 363748 39710
rect 363696 39646 363748 39652
rect 363892 34202 363920 289070
rect 363880 34196 363932 34202
rect 363880 34138 363932 34144
rect 363984 33998 364012 289614
rect 364076 216374 364104 333950
rect 370502 306912 370558 306921
rect 370502 306847 370558 306856
rect 367744 300484 367796 300490
rect 367744 300426 367796 300432
rect 365076 300280 365128 300286
rect 365076 300222 365128 300228
rect 364984 297696 365036 297702
rect 364984 297638 365036 297644
rect 364064 216368 364116 216374
rect 364064 216310 364116 216316
rect 364064 172576 364116 172582
rect 364064 172518 364116 172524
rect 364076 163062 364104 172518
rect 364064 163056 364116 163062
rect 364064 162998 364116 163004
rect 364064 158772 364116 158778
rect 364064 158714 364116 158720
rect 364076 84182 364104 158714
rect 364064 84176 364116 84182
rect 364064 84118 364116 84124
rect 363972 33992 364024 33998
rect 363972 33934 364024 33940
rect 364996 3806 365024 297638
rect 365088 42022 365116 300222
rect 366548 297628 366600 297634
rect 366548 297570 366600 297576
rect 365260 297560 365312 297566
rect 365166 297528 365222 297537
rect 365260 297502 365312 297508
rect 365166 297463 365222 297472
rect 365076 42016 365128 42022
rect 365076 41958 365128 41964
rect 365180 39506 365208 297463
rect 365168 39500 365220 39506
rect 365168 39442 365220 39448
rect 365272 39302 365300 297502
rect 365350 297392 365406 297401
rect 365350 297327 365406 297336
rect 365364 39370 365392 297327
rect 366456 294840 366508 294846
rect 366456 294782 366508 294788
rect 365444 294636 365496 294642
rect 365444 294578 365496 294584
rect 365456 40050 365484 294578
rect 366364 289536 366416 289542
rect 366364 289478 366416 289484
rect 365536 158024 365588 158030
rect 365536 157966 365588 157972
rect 365548 142186 365576 157966
rect 365536 142180 365588 142186
rect 365536 142122 365588 142128
rect 365536 126268 365588 126274
rect 365536 126210 365588 126216
rect 365548 119134 365576 126210
rect 365536 119128 365588 119134
rect 365536 119070 365588 119076
rect 365444 40044 365496 40050
rect 365444 39986 365496 39992
rect 365352 39364 365404 39370
rect 365352 39306 365404 39312
rect 365260 39296 365312 39302
rect 365260 39238 365312 39244
rect 366376 31618 366404 289478
rect 366468 36582 366496 294782
rect 366560 39846 366588 297570
rect 366732 295248 366784 295254
rect 366732 295190 366784 295196
rect 366640 289264 366692 289270
rect 366640 289206 366692 289212
rect 366548 39840 366600 39846
rect 366548 39782 366600 39788
rect 366456 36576 366508 36582
rect 366456 36518 366508 36524
rect 366652 34270 366680 289206
rect 366744 39982 366772 295190
rect 366824 185632 366876 185638
rect 366824 185574 366876 185580
rect 366836 172582 366864 185574
rect 366824 172576 366876 172582
rect 366824 172518 366876 172524
rect 367756 42566 367784 300426
rect 368020 300348 368072 300354
rect 368020 300290 368072 300296
rect 367928 300212 367980 300218
rect 367928 300154 367980 300160
rect 367836 300144 367888 300150
rect 367836 300086 367888 300092
rect 367848 42770 367876 300086
rect 367836 42764 367888 42770
rect 367836 42706 367888 42712
rect 367940 42702 367968 300154
rect 367928 42696 367980 42702
rect 367928 42638 367980 42644
rect 368032 42634 368060 300290
rect 368112 294908 368164 294914
rect 368112 294850 368164 294856
rect 368020 42628 368072 42634
rect 368020 42570 368072 42576
rect 367744 42560 367796 42566
rect 367744 42502 367796 42508
rect 366732 39976 366784 39982
rect 366732 39918 366784 39924
rect 368124 39914 368152 294850
rect 369308 294772 369360 294778
rect 369308 294714 369360 294720
rect 369216 294704 369268 294710
rect 369216 294646 369268 294652
rect 369124 289196 369176 289202
rect 369124 289138 369176 289144
rect 368204 273964 368256 273970
rect 368204 273906 368256 273912
rect 368216 45490 368244 273906
rect 368204 45484 368256 45490
rect 368204 45426 368256 45432
rect 368112 39908 368164 39914
rect 368112 39850 368164 39856
rect 366640 34264 366692 34270
rect 366640 34206 366692 34212
rect 369136 31686 369164 289138
rect 369228 36650 369256 294646
rect 369320 36718 369348 294714
rect 369400 289332 369452 289338
rect 369400 289274 369452 289280
rect 369308 36712 369360 36718
rect 369308 36654 369360 36660
rect 369216 36644 369268 36650
rect 369216 36586 369268 36592
rect 369412 34338 369440 289274
rect 369400 34332 369452 34338
rect 369400 34274 369452 34280
rect 369124 31680 369176 31686
rect 369124 31622 369176 31628
rect 366364 31612 366416 31618
rect 366364 31554 366416 31560
rect 364984 3800 365036 3806
rect 364984 3742 365036 3748
rect 363604 3732 363656 3738
rect 363604 3674 363656 3680
rect 362316 3664 362368 3670
rect 370516 3641 370544 306847
rect 373632 303000 373684 303006
rect 373632 302942 373684 302948
rect 371884 301504 371936 301510
rect 371884 301446 371936 301452
rect 370688 300756 370740 300762
rect 370688 300698 370740 300704
rect 370596 295180 370648 295186
rect 370596 295122 370648 295128
rect 370608 3942 370636 295122
rect 370700 42498 370728 300698
rect 370964 300688 371016 300694
rect 370964 300630 371016 300636
rect 370780 300552 370832 300558
rect 370780 300494 370832 300500
rect 370688 42492 370740 42498
rect 370688 42434 370740 42440
rect 370792 42294 370820 300494
rect 370872 300416 370924 300422
rect 370872 300358 370924 300364
rect 370884 42362 370912 300358
rect 370872 42356 370924 42362
rect 370872 42298 370924 42304
rect 370780 42288 370832 42294
rect 370780 42230 370832 42236
rect 370976 42226 371004 300630
rect 371056 300620 371108 300626
rect 371056 300562 371108 300568
rect 371068 42430 371096 300562
rect 371056 42424 371108 42430
rect 371056 42366 371108 42372
rect 370964 42220 371016 42226
rect 370964 42162 371016 42168
rect 371896 4078 371924 301446
rect 373448 300824 373500 300830
rect 373448 300766 373500 300772
rect 371974 297800 372030 297809
rect 371974 297735 372030 297744
rect 371884 4072 371936 4078
rect 371884 4014 371936 4020
rect 370596 3936 370648 3942
rect 370596 3878 370648 3884
rect 371988 3777 372016 297735
rect 373356 295044 373408 295050
rect 373356 294986 373408 294992
rect 372252 294976 372304 294982
rect 372252 294918 372304 294924
rect 372158 294536 372214 294545
rect 372158 294471 372214 294480
rect 372068 289604 372120 289610
rect 372068 289546 372120 289552
rect 372080 31210 372108 289546
rect 372068 31204 372120 31210
rect 372068 31146 372120 31152
rect 372172 3913 372200 294471
rect 372264 36854 372292 294918
rect 373264 286408 373316 286414
rect 373264 286350 373316 286356
rect 372344 286340 372396 286346
rect 372344 286282 372396 286288
rect 372252 36848 372304 36854
rect 372252 36790 372304 36796
rect 372356 31754 372384 286282
rect 372344 31748 372396 31754
rect 372344 31690 372396 31696
rect 373276 28626 373304 286350
rect 373368 36786 373396 294986
rect 373460 42158 373488 300766
rect 373538 300112 373594 300121
rect 373538 300047 373594 300056
rect 373448 42152 373500 42158
rect 373448 42094 373500 42100
rect 373552 42090 373580 300047
rect 373644 44674 373672 302942
rect 373632 44668 373684 44674
rect 373632 44610 373684 44616
rect 373540 42084 373592 42090
rect 373540 42026 373592 42032
rect 373356 36780 373408 36786
rect 373356 36722 373408 36728
rect 374656 28694 374684 385018
rect 374748 379438 374776 601666
rect 374828 577448 374880 577454
rect 374828 577390 374880 577396
rect 374840 572014 374868 577390
rect 374828 572008 374880 572014
rect 374828 571950 374880 571956
rect 376036 380866 376064 623766
rect 376208 572008 376260 572014
rect 376208 571950 376260 571956
rect 376220 568546 376248 571950
rect 376208 568540 376260 568546
rect 376208 568482 376260 568488
rect 377404 568540 377456 568546
rect 377404 568482 377456 568488
rect 377416 564126 377444 568482
rect 377404 564120 377456 564126
rect 377404 564062 377456 564068
rect 378796 382226 378824 645866
rect 380348 564120 380400 564126
rect 380348 564062 380400 564068
rect 380360 559230 380388 564062
rect 380348 559224 380400 559230
rect 380348 559166 380400 559172
rect 380256 386504 380308 386510
rect 380256 386446 380308 386452
rect 380164 386436 380216 386442
rect 380164 386378 380216 386384
rect 378784 382220 378836 382226
rect 378784 382162 378836 382168
rect 376024 380860 376076 380866
rect 376024 380802 376076 380808
rect 374736 379432 374788 379438
rect 374736 379374 374788 379380
rect 376022 306232 376078 306241
rect 376022 306167 376078 306176
rect 375932 300076 375984 300082
rect 375932 300018 375984 300024
rect 374736 295316 374788 295322
rect 374736 295258 374788 295264
rect 374748 36990 374776 295258
rect 375012 295112 375064 295118
rect 375012 295054 375064 295060
rect 374828 294568 374880 294574
rect 374828 294510 374880 294516
rect 374840 37058 374868 294510
rect 374920 289468 374972 289474
rect 374920 289410 374972 289416
rect 374828 37052 374880 37058
rect 374828 36994 374880 37000
rect 374736 36984 374788 36990
rect 374736 36926 374788 36932
rect 374932 31142 374960 289410
rect 375024 36922 375052 295054
rect 375104 291984 375156 291990
rect 375104 291926 375156 291932
rect 375116 37194 375144 291926
rect 375944 46374 375972 300018
rect 375932 46368 375984 46374
rect 375932 46310 375984 46316
rect 375104 37188 375156 37194
rect 375104 37130 375156 37136
rect 375012 36916 375064 36922
rect 375012 36858 375064 36864
rect 374920 31136 374972 31142
rect 374920 31078 374972 31084
rect 374644 28688 374696 28694
rect 374644 28630 374696 28636
rect 373264 28620 373316 28626
rect 373264 28562 373316 28568
rect 376036 6866 376064 306167
rect 379336 303544 379388 303550
rect 379336 303486 379388 303492
rect 376484 303476 376536 303482
rect 376484 303418 376536 303424
rect 376300 303408 376352 303414
rect 376300 303350 376352 303356
rect 376208 303068 376260 303074
rect 376208 303010 376260 303016
rect 376116 286476 376168 286482
rect 376116 286418 376168 286424
rect 376128 28558 376156 286418
rect 376220 44810 376248 303010
rect 376312 45286 376340 303350
rect 376392 303136 376444 303142
rect 376392 303078 376444 303084
rect 376300 45280 376352 45286
rect 376300 45222 376352 45228
rect 376404 45218 376432 303078
rect 376392 45212 376444 45218
rect 376392 45154 376444 45160
rect 376208 44804 376260 44810
rect 376208 44746 376260 44752
rect 376496 44742 376524 303418
rect 379152 303340 379204 303346
rect 379152 303282 379204 303288
rect 379060 303272 379112 303278
rect 379060 303214 379112 303220
rect 378968 303204 379020 303210
rect 378968 303146 379020 303152
rect 378692 302796 378744 302802
rect 378692 302738 378744 302744
rect 376668 299940 376720 299946
rect 376668 299882 376720 299888
rect 376576 292052 376628 292058
rect 376576 291994 376628 292000
rect 376484 44736 376536 44742
rect 376484 44678 376536 44684
rect 376588 37126 376616 291994
rect 376680 45422 376708 299882
rect 378600 292392 378652 292398
rect 378600 292334 378652 292340
rect 377680 292256 377732 292262
rect 377680 292198 377732 292204
rect 377588 292188 377640 292194
rect 377588 292130 377640 292136
rect 377496 289400 377548 289406
rect 377496 289342 377548 289348
rect 377404 286748 377456 286754
rect 377404 286690 377456 286696
rect 376668 45416 376720 45422
rect 376668 45358 376720 45364
rect 376576 37120 376628 37126
rect 376576 37062 376628 37068
rect 376116 28552 376168 28558
rect 376116 28494 376168 28500
rect 377416 28354 377444 286690
rect 377508 31346 377536 289342
rect 377600 34406 377628 292130
rect 377692 37262 377720 292198
rect 377680 37256 377732 37262
rect 377680 37198 377732 37204
rect 378612 36514 378640 292334
rect 378704 46442 378732 302738
rect 378784 302660 378836 302666
rect 378784 302602 378836 302608
rect 378692 46436 378744 46442
rect 378692 46378 378744 46384
rect 378600 36508 378652 36514
rect 378600 36450 378652 36456
rect 377588 34400 377640 34406
rect 377588 34342 377640 34348
rect 378796 33114 378824 302602
rect 378876 286544 378928 286550
rect 378876 286486 378928 286492
rect 378784 33108 378836 33114
rect 378784 33050 378836 33056
rect 377496 31340 377548 31346
rect 377496 31282 377548 31288
rect 378888 28490 378916 286486
rect 378980 45082 379008 303146
rect 378968 45076 379020 45082
rect 378968 45018 379020 45024
rect 379072 45014 379100 303214
rect 379164 45150 379192 303282
rect 379242 302832 379298 302841
rect 379242 302767 379298 302776
rect 379152 45144 379204 45150
rect 379152 45086 379204 45092
rect 379060 45008 379112 45014
rect 379060 44950 379112 44956
rect 379256 44946 379284 302767
rect 379348 46510 379376 303486
rect 379428 302864 379480 302870
rect 379428 302806 379480 302812
rect 379440 46578 379468 302806
rect 379428 46572 379480 46578
rect 379428 46514 379480 46520
rect 379336 46504 379388 46510
rect 379336 46446 379388 46452
rect 379244 44940 379296 44946
rect 379244 44882 379296 44888
rect 380176 31006 380204 386378
rect 380268 34474 380296 386446
rect 381556 383654 381584 667898
rect 406384 656192 406436 656198
rect 406384 656134 406436 656140
rect 384948 559224 385000 559230
rect 384948 559166 385000 559172
rect 384960 554826 384988 559166
rect 384960 554798 385080 554826
rect 385052 552022 385080 554798
rect 385040 552016 385092 552022
rect 385040 551958 385092 551964
rect 387064 552016 387116 552022
rect 387064 551958 387116 551964
rect 387076 540938 387104 551958
rect 387064 540932 387116 540938
rect 387064 540874 387116 540880
rect 388444 540932 388496 540938
rect 388444 540874 388496 540880
rect 388456 517546 388484 540874
rect 388444 517540 388496 517546
rect 388444 517482 388496 517488
rect 389456 517540 389508 517546
rect 389456 517482 389508 517488
rect 389468 512038 389496 517482
rect 389456 512032 389508 512038
rect 389456 511974 389508 511980
rect 393228 511964 393280 511970
rect 393228 511906 393280 511912
rect 393240 509130 393268 511906
rect 393240 509102 393360 509130
rect 393332 506802 393360 509102
rect 393320 506796 393372 506802
rect 393320 506738 393372 506744
rect 396724 506796 396776 506802
rect 396724 506738 396776 506744
rect 396736 476134 396764 506738
rect 396724 476128 396776 476134
rect 396724 476070 396776 476076
rect 400864 476060 400916 476066
rect 400864 476002 400916 476008
rect 400876 468246 400904 476002
rect 400864 468240 400916 468246
rect 400864 468182 400916 468188
rect 401968 468240 402020 468246
rect 401968 468182 402020 468188
rect 401980 465050 402008 468182
rect 401968 465044 402020 465050
rect 401968 464986 402020 464992
rect 403624 465044 403676 465050
rect 403624 464986 403676 464992
rect 383016 458244 383068 458250
rect 383016 458186 383068 458192
rect 382924 386572 382976 386578
rect 382924 386514 382976 386520
rect 381544 383648 381596 383654
rect 381544 383590 381596 383596
rect 380346 306776 380402 306785
rect 380346 306711 380402 306720
rect 380256 34468 380308 34474
rect 380256 34410 380308 34416
rect 380164 31000 380216 31006
rect 380164 30942 380216 30948
rect 378876 28484 378928 28490
rect 378876 28426 378928 28432
rect 377404 28348 377456 28354
rect 377404 28290 377456 28296
rect 376024 6860 376076 6866
rect 376024 6802 376076 6808
rect 372158 3904 372214 3913
rect 372158 3839 372214 3848
rect 371974 3768 372030 3777
rect 371974 3703 372030 3712
rect 362316 3606 362368 3612
rect 370502 3632 370558 3641
rect 370502 3567 370558 3576
rect 380360 3466 380388 306711
rect 381818 306096 381874 306105
rect 381728 306060 381780 306066
rect 381818 306031 381874 306040
rect 381728 306002 381780 306008
rect 381634 305960 381690 305969
rect 381634 305895 381690 305904
rect 381544 305856 381596 305862
rect 381544 305798 381596 305804
rect 381450 302968 381506 302977
rect 381450 302903 381506 302912
rect 380532 292460 380584 292466
rect 380532 292402 380584 292408
rect 380440 289808 380492 289814
rect 380440 289750 380492 289756
rect 380452 31278 380480 289750
rect 380544 33794 380572 292402
rect 381360 160132 381412 160138
rect 381360 160074 381412 160080
rect 381372 95198 381400 160074
rect 381360 95192 381412 95198
rect 381360 95134 381412 95140
rect 381464 44878 381492 302903
rect 381556 46646 381584 305798
rect 381544 46640 381596 46646
rect 381544 46582 381596 46588
rect 381452 44872 381504 44878
rect 381452 44814 381504 44820
rect 380532 33788 380584 33794
rect 380532 33730 380584 33736
rect 380440 31272 380492 31278
rect 380440 31214 380492 31220
rect 380348 3460 380400 3466
rect 380348 3402 380400 3408
rect 361120 3392 361172 3398
rect 361120 3334 361172 3340
rect 361028 3256 361080 3262
rect 361028 3198 361080 3204
rect 381648 2106 381676 305895
rect 381740 46714 381768 306002
rect 381728 46708 381780 46714
rect 381728 46650 381780 46656
rect 381832 3505 381860 306031
rect 382186 303104 382242 303113
rect 382186 303039 382242 303048
rect 382096 302728 382148 302734
rect 382096 302670 382148 302676
rect 382004 292120 382056 292126
rect 382004 292062 382056 292068
rect 381912 286612 381964 286618
rect 381912 286554 381964 286560
rect 381924 28422 381952 286554
rect 382016 34066 382044 292062
rect 382108 45558 382136 302670
rect 382096 45552 382148 45558
rect 382096 45494 382148 45500
rect 382200 44849 382228 303039
rect 382186 44840 382242 44849
rect 382186 44775 382242 44784
rect 382004 34060 382056 34066
rect 382004 34002 382056 34008
rect 382936 33726 382964 386514
rect 383028 371210 383056 458186
rect 403636 456822 403664 464986
rect 403624 456816 403676 456822
rect 403624 456758 403676 456764
rect 406396 383586 406424 656134
rect 407764 634840 407816 634846
rect 407764 634782 407816 634788
rect 406384 383580 406436 383586
rect 406384 383522 406436 383528
rect 407776 382158 407804 634782
rect 410524 612808 410576 612814
rect 410524 612750 410576 612756
rect 408408 456748 408460 456754
rect 408408 456690 408460 456696
rect 408420 455410 408448 456690
rect 408420 455382 408540 455410
rect 408512 452606 408540 455382
rect 408500 452600 408552 452606
rect 408500 452542 408552 452548
rect 410340 452600 410392 452606
rect 410340 452542 410392 452548
rect 410352 447098 410380 452542
rect 410340 447092 410392 447098
rect 410340 447034 410392 447040
rect 407764 382152 407816 382158
rect 407764 382094 407816 382100
rect 410536 380798 410564 612750
rect 411904 524476 411956 524482
rect 411904 524418 411956 524424
rect 410524 380792 410576 380798
rect 410524 380734 410576 380740
rect 411916 375290 411944 524418
rect 411904 375284 411956 375290
rect 411904 375226 411956 375232
rect 383016 371204 383068 371210
rect 383016 371146 383068 371152
rect 394700 351960 394752 351966
rect 394700 351902 394752 351908
rect 385776 338156 385828 338162
rect 385776 338098 385828 338104
rect 384304 306332 384356 306338
rect 384304 306274 384356 306280
rect 383014 300248 383070 300257
rect 383014 300183 383070 300192
rect 382924 33720 382976 33726
rect 382924 33662 382976 33668
rect 381912 28416 381964 28422
rect 381912 28358 381964 28364
rect 381818 3496 381874 3505
rect 381818 3431 381874 3440
rect 383028 2174 383056 300183
rect 383292 292528 383344 292534
rect 383292 292470 383344 292476
rect 383200 289740 383252 289746
rect 383200 289682 383252 289688
rect 383108 286816 383160 286822
rect 383108 286758 383160 286764
rect 383120 3534 383148 286758
rect 383212 31482 383240 289682
rect 383304 33862 383332 292470
rect 383384 275324 383436 275330
rect 383384 275266 383436 275272
rect 383292 33856 383344 33862
rect 383292 33798 383344 33804
rect 383200 31476 383252 31482
rect 383200 31418 383252 31424
rect 383396 20670 383424 275266
rect 383476 160472 383528 160478
rect 383476 160414 383528 160420
rect 383488 73166 383516 160414
rect 383476 73160 383528 73166
rect 383476 73102 383528 73108
rect 384316 46782 384344 306274
rect 384488 306196 384540 306202
rect 384488 306138 384540 306144
rect 384396 305584 384448 305590
rect 384396 305526 384448 305532
rect 384304 46776 384356 46782
rect 384304 46718 384356 46724
rect 384408 46306 384436 305526
rect 384500 46850 384528 306138
rect 384580 306128 384632 306134
rect 384580 306070 384632 306076
rect 384488 46844 384540 46850
rect 384488 46786 384540 46792
rect 384592 46753 384620 306070
rect 384948 305992 385000 305998
rect 384948 305934 385000 305940
rect 384672 305924 384724 305930
rect 384672 305866 384724 305872
rect 384578 46744 384634 46753
rect 384578 46679 384634 46688
rect 384396 46300 384448 46306
rect 384396 46242 384448 46248
rect 384684 46238 384712 305866
rect 384856 297832 384908 297838
rect 384856 297774 384908 297780
rect 384762 289096 384818 289105
rect 384762 289031 384818 289040
rect 384672 46232 384724 46238
rect 384672 46174 384724 46180
rect 384776 31074 384804 289031
rect 384868 39438 384896 297774
rect 384960 47025 384988 305934
rect 385684 297900 385736 297906
rect 385684 297842 385736 297848
rect 385592 160336 385644 160342
rect 385592 160278 385644 160284
rect 385604 62082 385632 160278
rect 385592 62076 385644 62082
rect 385592 62018 385644 62024
rect 385592 51128 385644 51134
rect 385592 51070 385644 51076
rect 384946 47016 385002 47025
rect 384946 46951 385002 46960
rect 384856 39432 384908 39438
rect 384856 39374 384908 39380
rect 385604 31754 385632 51070
rect 385592 31748 385644 31754
rect 385592 31690 385644 31696
rect 384764 31068 384816 31074
rect 384764 31010 384816 31016
rect 383384 20664 383436 20670
rect 383384 20606 383436 20612
rect 383108 3528 383160 3534
rect 383108 3470 383160 3476
rect 385696 2242 385724 297842
rect 385788 293962 385816 338098
rect 386052 306264 386104 306270
rect 386052 306206 386104 306212
rect 385960 305516 386012 305522
rect 385960 305458 386012 305464
rect 385868 304428 385920 304434
rect 385868 304370 385920 304376
rect 385776 293956 385828 293962
rect 385776 293898 385828 293904
rect 385776 291780 385828 291786
rect 385776 291722 385828 291728
rect 385788 3602 385816 291722
rect 385880 31550 385908 304370
rect 385972 46889 386000 305458
rect 386064 46918 386092 306206
rect 386328 292324 386380 292330
rect 386328 292266 386380 292272
rect 386236 289060 386288 289066
rect 386236 289002 386288 289008
rect 386144 286680 386196 286686
rect 386144 286622 386196 286628
rect 386052 46912 386104 46918
rect 385958 46880 386014 46889
rect 386052 46854 386104 46860
rect 385958 46815 386014 46824
rect 385868 31544 385920 31550
rect 385868 31486 385920 31492
rect 386156 28286 386184 286622
rect 386248 31414 386276 289002
rect 386340 33930 386368 292266
rect 388444 193860 388496 193866
rect 388444 193802 388496 193808
rect 388456 185638 388484 193802
rect 388444 185632 388496 185638
rect 388444 185574 388496 185580
rect 391112 181484 391164 181490
rect 391112 181426 391164 181432
rect 391124 175982 391152 181426
rect 391112 175976 391164 175982
rect 391112 175918 391164 175924
rect 393964 167068 394016 167074
rect 393964 167010 394016 167016
rect 393976 158030 394004 167010
rect 393964 158024 394016 158030
rect 393964 157966 394016 157972
rect 393964 150476 394016 150482
rect 393964 150418 394016 150424
rect 390192 149388 390244 149394
rect 390192 149330 390244 149336
rect 390204 143138 390232 149330
rect 387064 143132 387116 143138
rect 387064 143074 387116 143080
rect 390192 143132 390244 143138
rect 390192 143074 390244 143080
rect 387076 126274 387104 143074
rect 393976 129810 394004 150418
rect 390560 129804 390612 129810
rect 390560 129746 390612 129752
rect 393964 129804 394016 129810
rect 393964 129746 394016 129752
rect 390572 127634 390600 129746
rect 390560 127628 390612 127634
rect 390560 127570 390612 127576
rect 387064 126268 387116 126274
rect 387064 126210 387116 126216
rect 394712 113174 394740 351902
rect 405740 350600 405792 350606
rect 405740 350542 405792 350548
rect 402244 347812 402296 347818
rect 402244 347754 402296 347760
rect 402256 342922 402284 347754
rect 402244 342916 402296 342922
rect 402244 342858 402296 342864
rect 402980 342916 403032 342922
rect 402980 342858 403032 342864
rect 399484 339516 399536 339522
rect 399484 339458 399536 339464
rect 399496 315994 399524 339458
rect 402992 339454 403020 342858
rect 401600 339448 401652 339454
rect 401600 339390 401652 339396
rect 402980 339448 403032 339454
rect 402980 339390 403032 339396
rect 401612 334914 401640 339390
rect 401612 334886 402086 334914
rect 405752 334900 405780 350542
rect 412652 338774 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 416044 700664 416096 700670
rect 416044 700606 416096 700612
rect 414664 513392 414716 513398
rect 414664 513334 414716 513340
rect 413284 447092 413336 447098
rect 413284 447034 413336 447040
rect 413296 438326 413324 447034
rect 413284 438320 413336 438326
rect 413284 438262 413336 438268
rect 414676 373998 414704 513334
rect 414756 438320 414808 438326
rect 414756 438262 414808 438268
rect 414768 426426 414796 438262
rect 414756 426420 414808 426426
rect 414756 426362 414808 426368
rect 414664 373992 414716 373998
rect 414664 373934 414716 373940
rect 412640 338768 412692 338774
rect 412640 338710 412692 338716
rect 416056 336258 416084 700606
rect 429856 700330 429884 703520
rect 446496 700936 446548 700942
rect 446496 700878 446548 700884
rect 445024 700868 445076 700874
rect 445024 700810 445076 700816
rect 444288 700528 444340 700534
rect 444288 700470 444340 700476
rect 444104 700460 444156 700466
rect 444104 700402 444156 700408
rect 418804 700324 418856 700330
rect 418804 700266 418856 700272
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 416136 502376 416188 502382
rect 416136 502318 416188 502324
rect 416148 373930 416176 502318
rect 417424 491360 417476 491366
rect 417424 491302 417476 491308
rect 416136 373924 416188 373930
rect 416136 373866 416188 373872
rect 417436 372570 417464 491302
rect 417516 426420 417568 426426
rect 417516 426362 417568 426368
rect 417528 420510 417556 426362
rect 417516 420504 417568 420510
rect 417516 420446 417568 420452
rect 417424 372564 417476 372570
rect 417424 372506 417476 372512
rect 416780 336932 416832 336938
rect 416780 336874 416832 336880
rect 416044 336252 416096 336258
rect 416044 336194 416096 336200
rect 409420 335436 409472 335442
rect 409420 335378 409472 335384
rect 409432 334900 409460 335378
rect 413100 335368 413152 335374
rect 413100 335310 413152 335316
rect 413112 334900 413140 335310
rect 416792 334900 416820 336874
rect 418816 336122 418844 700266
rect 418988 685160 419040 685166
rect 418988 685102 419040 685108
rect 418896 684820 418948 684826
rect 418896 684762 418948 684768
rect 418908 336190 418936 684762
rect 419000 336326 419028 685102
rect 420184 684752 420236 684758
rect 420184 684694 420236 684700
rect 420092 682780 420144 682786
rect 420092 682722 420144 682728
rect 419080 480276 419132 480282
rect 419080 480218 419132 480224
rect 419092 372502 419120 480218
rect 419172 436144 419224 436150
rect 419172 436086 419224 436092
rect 419080 372496 419132 372502
rect 419080 372438 419132 372444
rect 419184 369850 419212 436086
rect 419172 369844 419224 369850
rect 419172 369786 419224 369792
rect 418988 336320 419040 336326
rect 418988 336262 419040 336268
rect 418896 336184 418948 336190
rect 418896 336126 418948 336132
rect 418804 336116 418856 336122
rect 418804 336058 418856 336064
rect 420104 334626 420132 682722
rect 420196 334694 420224 684694
rect 420276 684684 420328 684690
rect 420276 684626 420328 684632
rect 420288 334898 420316 684626
rect 420368 684616 420420 684622
rect 420368 684558 420420 684564
rect 420380 335102 420408 684558
rect 420552 683528 420604 683534
rect 420552 683470 420604 683476
rect 420460 336796 420512 336802
rect 420460 336738 420512 336744
rect 420368 335096 420420 335102
rect 420368 335038 420420 335044
rect 420276 334892 420328 334898
rect 420276 334834 420328 334840
rect 420184 334688 420236 334694
rect 420184 334630 420236 334636
rect 420472 334642 420500 336738
rect 420564 335102 420592 683470
rect 420644 683460 420696 683466
rect 420644 683402 420696 683408
rect 420552 335096 420604 335102
rect 420552 335038 420604 335044
rect 420656 335034 420684 683402
rect 420736 683392 420788 683398
rect 420736 683334 420788 683340
rect 420644 335028 420696 335034
rect 420644 334970 420696 334976
rect 420748 334762 420776 683334
rect 420826 682816 420882 682825
rect 420826 682751 420882 682760
rect 420840 334830 420868 682751
rect 436100 462460 436152 462466
rect 436100 462402 436152 462408
rect 431960 462392 432012 462398
rect 431960 462334 432012 462340
rect 423588 455456 423640 455462
rect 423588 455398 423640 455404
rect 423600 447574 423628 455398
rect 422484 447568 422536 447574
rect 422484 447510 422536 447516
rect 423588 447568 423640 447574
rect 423588 447510 423640 447516
rect 422496 444924 422524 447510
rect 423600 447166 423628 447510
rect 427452 447228 427504 447234
rect 427452 447170 427504 447176
rect 423588 447160 423640 447166
rect 423588 447102 423640 447108
rect 427464 444924 427492 447170
rect 431972 444530 432000 462334
rect 436112 445738 436140 462402
rect 443368 447160 443420 447166
rect 443368 447102 443420 447108
rect 436100 445732 436152 445738
rect 436100 445674 436152 445680
rect 437388 445732 437440 445738
rect 437388 445674 437440 445680
rect 437400 444938 437428 445674
rect 437308 444924 437428 444938
rect 437308 444910 437414 444924
rect 432696 444576 432748 444582
rect 431972 444524 432696 444530
rect 431972 444518 432748 444524
rect 431972 444502 432736 444518
rect 437308 444514 437336 444910
rect 437296 444508 437348 444514
rect 437296 444450 437348 444456
rect 442632 444440 442684 444446
rect 442382 444388 442632 444394
rect 442382 444382 442684 444388
rect 442382 444366 442672 444382
rect 443380 444378 443408 447102
rect 443368 444372 443420 444378
rect 443368 444314 443420 444320
rect 444116 421977 444144 700402
rect 444196 423428 444248 423434
rect 444196 423370 444248 423376
rect 444208 422226 444236 423370
rect 444300 422294 444328 700470
rect 444300 422266 444420 422294
rect 444208 422198 444328 422226
rect 444194 422104 444250 422113
rect 444194 422039 444250 422048
rect 444102 421968 444158 421977
rect 444102 421903 444158 421912
rect 424324 420504 424376 420510
rect 424324 420446 424376 420452
rect 421484 417790 421512 420036
rect 421472 417784 421524 417790
rect 421472 417726 421524 417732
rect 422128 417450 422156 420036
rect 422312 420022 422786 420050
rect 422864 420022 423430 420050
rect 422116 417444 422168 417450
rect 422116 417386 422168 417392
rect 422312 389842 422340 420022
rect 422864 412634 422892 420022
rect 424060 417586 424088 420036
rect 424048 417580 424100 417586
rect 424048 417522 424100 417528
rect 422404 412606 422892 412634
rect 422404 391270 422432 412606
rect 422392 391264 422444 391270
rect 422392 391206 422444 391212
rect 422300 389836 422352 389842
rect 422300 389778 422352 389784
rect 424336 352102 424364 420446
rect 424704 417518 424732 420036
rect 425348 417654 425376 420036
rect 425992 417722 426020 420036
rect 443644 418804 443696 418810
rect 443644 418746 443696 418752
rect 425980 417716 426032 417722
rect 425980 417658 426032 417664
rect 425336 417648 425388 417654
rect 425336 417590 425388 417596
rect 424692 417512 424744 417518
rect 424692 417454 424744 417460
rect 440884 416084 440936 416090
rect 440884 416026 440936 416032
rect 436744 413296 436796 413302
rect 436744 413238 436796 413244
rect 436756 371142 436784 413238
rect 439504 403028 439556 403034
rect 439504 402970 439556 402976
rect 436744 371136 436796 371142
rect 436744 371078 436796 371084
rect 439516 367062 439544 402970
rect 440896 369782 440924 416026
rect 442264 414044 442316 414050
rect 442264 413986 442316 413992
rect 440976 392012 441028 392018
rect 440976 391954 441028 391960
rect 440884 369776 440936 369782
rect 440884 369718 440936 369724
rect 439504 367056 439556 367062
rect 439504 366998 439556 367004
rect 440988 366994 441016 391954
rect 442276 368422 442304 413986
rect 442814 387152 442870 387161
rect 442814 387087 442870 387096
rect 442356 380928 442408 380934
rect 442356 380870 442408 380876
rect 442264 368416 442316 368422
rect 442264 368358 442316 368364
rect 440976 366988 441028 366994
rect 440976 366930 441028 366936
rect 442368 365634 442396 380870
rect 442356 365628 442408 365634
rect 442356 365570 442408 365576
rect 442264 363044 442316 363050
rect 442264 362986 442316 362992
rect 432604 362976 432656 362982
rect 432604 362918 432656 362924
rect 424324 352096 424376 352102
rect 424324 352038 424376 352044
rect 426900 352096 426952 352102
rect 426900 352038 426952 352044
rect 426912 347682 426940 352038
rect 426900 347676 426952 347682
rect 426900 347618 426952 347624
rect 430580 347676 430632 347682
rect 430580 347618 430632 347624
rect 430592 342242 430620 347618
rect 430580 342236 430632 342242
rect 430580 342178 430632 342184
rect 431408 336932 431460 336938
rect 431408 336874 431460 336880
rect 424140 336864 424192 336870
rect 424140 336806 424192 336812
rect 429936 336864 429988 336870
rect 429936 336806 429988 336812
rect 424152 334900 424180 336806
rect 420828 334824 420880 334830
rect 420828 334766 420880 334772
rect 420736 334756 420788 334762
rect 420736 334698 420788 334704
rect 420472 334628 420592 334642
rect 420092 334620 420144 334626
rect 420486 334614 420592 334628
rect 420092 334562 420144 334568
rect 420564 334506 420592 334614
rect 420734 334520 420790 334529
rect 420486 334478 420734 334506
rect 428094 334520 428150 334529
rect 427846 334478 428094 334506
rect 420734 334455 420790 334464
rect 428094 334455 428150 334464
rect 428108 334422 428136 334455
rect 428096 334416 428148 334422
rect 428096 334358 428148 334364
rect 429844 332648 429896 332654
rect 429844 332590 429896 332596
rect 399484 315988 399536 315994
rect 399484 315930 399536 315936
rect 426348 305788 426400 305794
rect 426348 305730 426400 305736
rect 407120 301572 407172 301578
rect 407120 301514 407172 301520
rect 406292 207664 406344 207670
rect 406292 207606 406344 207612
rect 406304 200802 406332 207606
rect 401600 200796 401652 200802
rect 401600 200738 401652 200744
rect 406292 200796 406344 200802
rect 406292 200738 406344 200744
rect 401612 193866 401640 200738
rect 406384 195288 406436 195294
rect 406384 195230 406436 195236
rect 401600 193860 401652 193866
rect 401600 193802 401652 193808
rect 406396 188426 406424 195230
rect 402244 188420 402296 188426
rect 402244 188362 402296 188368
rect 406384 188420 406436 188426
rect 406384 188362 406436 188368
rect 398840 188352 398892 188358
rect 398840 188294 398892 188300
rect 398852 181490 398880 188294
rect 398840 181484 398892 181490
rect 398840 181426 398892 181432
rect 396724 178696 396776 178702
rect 396724 178638 396776 178644
rect 396736 167074 396764 178638
rect 402256 178090 402284 188362
rect 398104 178084 398156 178090
rect 398104 178026 398156 178032
rect 402244 178084 402296 178090
rect 402244 178026 402296 178032
rect 396724 167068 396776 167074
rect 396724 167010 396776 167016
rect 398116 160206 398144 178026
rect 403624 161764 403676 161770
rect 403624 161706 403676 161712
rect 395344 160200 395396 160206
rect 395344 160142 395396 160148
rect 398104 160200 398156 160206
rect 398104 160142 398156 160148
rect 395356 149394 395384 160142
rect 398104 159384 398156 159390
rect 398104 159326 398156 159332
rect 398116 150482 398144 159326
rect 398104 150476 398156 150482
rect 398104 150418 398156 150424
rect 395344 149388 395396 149394
rect 395344 149330 395396 149336
rect 403636 117298 403664 161706
rect 406384 160200 406436 160206
rect 406384 160142 406436 160148
rect 403624 117292 403676 117298
rect 403624 117234 403676 117240
rect 394712 113146 395292 113174
rect 389824 107024 389876 107030
rect 389824 106966 389876 106972
rect 389836 104938 389864 106966
rect 389528 104910 389864 104938
rect 395264 104938 395292 113146
rect 406396 107030 406424 160142
rect 407132 113174 407160 301514
rect 424324 267028 424376 267034
rect 424324 266970 424376 266976
rect 424336 230518 424364 266970
rect 421564 230512 421616 230518
rect 421564 230454 421616 230460
rect 424324 230512 424376 230518
rect 424324 230454 424376 230460
rect 414664 220108 414716 220114
rect 414664 220050 414716 220056
rect 413284 218068 413336 218074
rect 413284 218010 413336 218016
rect 411260 206304 411312 206310
rect 411260 206246 411312 206252
rect 410524 186312 410576 186318
rect 410524 186254 410576 186260
rect 410536 178702 410564 186254
rect 410524 178696 410576 178702
rect 410524 178638 410576 178644
rect 411272 171134 411300 206246
rect 411352 191140 411404 191146
rect 411352 191082 411404 191088
rect 411364 188358 411392 191082
rect 411352 188352 411404 188358
rect 411352 188294 411404 188300
rect 413296 186318 413324 218010
rect 413284 186312 413336 186318
rect 413284 186254 413336 186260
rect 414676 171134 414704 220050
rect 421576 218074 421604 230454
rect 425704 220856 425756 220862
rect 425704 220798 425756 220804
rect 421564 218068 421616 218074
rect 421564 218010 421616 218016
rect 424324 209092 424376 209098
rect 424324 209034 424376 209040
rect 421564 200796 421616 200802
rect 421564 200738 421616 200744
rect 421576 179450 421604 200738
rect 424336 195294 424364 209034
rect 424324 195288 424376 195294
rect 424324 195230 424376 195236
rect 425716 194750 425744 220798
rect 425796 213240 425848 213246
rect 425796 213182 425848 213188
rect 425808 207670 425836 213182
rect 425796 207664 425848 207670
rect 425796 207606 425848 207612
rect 422852 194744 422904 194750
rect 422852 194686 422904 194692
rect 425704 194744 425756 194750
rect 425704 194686 425756 194692
rect 422864 191146 422892 194686
rect 422852 191140 422904 191146
rect 422852 191082 422904 191088
rect 416044 179444 416096 179450
rect 416044 179386 416096 179392
rect 421564 179444 421616 179450
rect 421564 179386 421616 179392
rect 411272 171106 411392 171134
rect 414676 171106 414796 171134
rect 410248 164892 410300 164898
rect 410248 164834 410300 164840
rect 410260 162314 410288 164834
rect 407764 162308 407816 162314
rect 407764 162250 407816 162256
rect 410248 162308 410300 162314
rect 410248 162250 410300 162256
rect 407776 159390 407804 162250
rect 407856 161560 407908 161566
rect 407856 161502 407908 161508
rect 407764 159384 407816 159390
rect 407764 159326 407816 159332
rect 407868 142154 407896 161502
rect 410616 160404 410668 160410
rect 410616 160346 410668 160352
rect 410524 160268 410576 160274
rect 410524 160210 410576 160216
rect 407776 142126 407896 142154
rect 407776 139398 407804 142126
rect 407764 139392 407816 139398
rect 407764 139334 407816 139340
rect 407132 113146 407620 113174
rect 406384 107024 406436 107030
rect 406384 106966 406436 106972
rect 402152 106956 402204 106962
rect 402152 106898 402204 106904
rect 402164 104938 402192 106898
rect 395264 104910 395692 104938
rect 401856 104910 402192 104938
rect 407592 104938 407620 113146
rect 410536 106282 410564 160210
rect 410628 128314 410656 160346
rect 411364 159882 411392 171106
rect 414768 160342 414796 171106
rect 416056 164898 416084 179386
rect 416044 164892 416096 164898
rect 416044 164834 416096 164840
rect 421562 162752 421618 162761
rect 421562 162687 421618 162696
rect 418712 162172 418764 162178
rect 418712 162114 418764 162120
rect 418160 160472 418212 160478
rect 418160 160414 418212 160420
rect 414756 160336 414808 160342
rect 414756 160278 414808 160284
rect 414768 159882 414796 160278
rect 418172 159882 418200 160414
rect 418724 159882 418752 162114
rect 421576 161634 421604 162687
rect 426360 161702 426388 305730
rect 429856 194546 429884 332590
rect 429948 326398 429976 336806
rect 431316 335436 431368 335442
rect 431316 335378 431368 335384
rect 431224 327140 431276 327146
rect 431224 327082 431276 327088
rect 429936 326392 429988 326398
rect 429936 326334 429988 326340
rect 429844 194540 429896 194546
rect 429844 194482 429896 194488
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 426348 161696 426400 161702
rect 426348 161638 426400 161644
rect 421564 161628 421616 161634
rect 421564 161570 421616 161576
rect 411364 159854 411792 159882
rect 414768 159854 415104 159882
rect 418172 159854 418752 159882
rect 421380 159384 421432 159390
rect 421576 159338 421604 161570
rect 426360 160138 426388 161638
rect 428660 160274 428688 162687
rect 431236 161770 431264 327082
rect 431328 323610 431356 335378
rect 431420 325650 431448 336874
rect 432616 332897 432644 362918
rect 435456 361616 435508 361622
rect 435456 361558 435508 361564
rect 432788 348424 432840 348430
rect 432788 348366 432840 348372
rect 432800 345014 432828 348366
rect 432800 344986 433012 345014
rect 432788 344344 432840 344350
rect 432788 344286 432840 344292
rect 432696 342236 432748 342242
rect 432696 342178 432748 342184
rect 432708 336734 432736 342178
rect 432696 336728 432748 336734
rect 432696 336670 432748 336676
rect 432800 336546 432828 344286
rect 432708 336518 432828 336546
rect 432602 332888 432658 332897
rect 432602 332823 432658 332832
rect 432604 330268 432656 330274
rect 432604 330210 432656 330216
rect 431408 325644 431460 325650
rect 431408 325586 431460 325592
rect 431316 323604 431368 323610
rect 431316 323546 431368 323552
rect 432144 318164 432196 318170
rect 432144 318106 432196 318112
rect 432156 314537 432184 318106
rect 432142 314528 432198 314537
rect 432142 314463 432198 314472
rect 432616 310865 432644 330210
rect 432708 325553 432736 336518
rect 432984 336410 433012 344986
rect 435364 338224 435416 338230
rect 435364 338166 435416 338172
rect 433984 336728 434036 336734
rect 433984 336670 434036 336676
rect 432800 336382 433012 336410
rect 432800 329225 432828 336382
rect 432880 331900 432932 331906
rect 432880 331842 432932 331848
rect 432786 329216 432842 329225
rect 432786 329151 432842 329160
rect 432694 325544 432750 325553
rect 432694 325479 432750 325488
rect 432892 318209 432920 331842
rect 432972 328704 433024 328710
rect 432972 328646 433024 328652
rect 432984 321881 433012 328646
rect 433996 328438 434024 336670
rect 433984 328432 434036 328438
rect 433984 328374 434036 328380
rect 432970 321872 433026 321881
rect 432970 321807 433026 321816
rect 432878 318200 432934 318209
rect 432878 318135 432934 318144
rect 432602 310856 432658 310865
rect 432602 310791 432658 310800
rect 432236 307760 432288 307766
rect 432236 307702 432288 307708
rect 432248 307193 432276 307702
rect 432234 307184 432290 307193
rect 432234 307119 432290 307128
rect 435376 282878 435404 338166
rect 435468 328710 435496 361558
rect 439596 360256 439648 360262
rect 439596 360198 439648 360204
rect 436836 358828 436888 358834
rect 436836 358770 436888 358776
rect 435548 335368 435600 335374
rect 435548 335310 435600 335316
rect 435456 328704 435508 328710
rect 435456 328646 435508 328652
rect 435560 325514 435588 335310
rect 436744 331356 436796 331362
rect 436744 331298 436796 331304
rect 436008 328500 436060 328506
rect 436008 328442 436060 328448
rect 435548 325508 435600 325514
rect 435548 325450 435600 325456
rect 435364 282872 435416 282878
rect 435364 282814 435416 282820
rect 433984 272536 434036 272542
rect 433984 272478 434036 272484
rect 433996 267034 434024 272478
rect 433984 267028 434036 267034
rect 433984 266970 434036 266976
rect 433984 260160 434036 260166
rect 433984 260102 434036 260108
rect 433708 255332 433760 255338
rect 433708 255274 433760 255280
rect 433720 248470 433748 255274
rect 431316 248464 431368 248470
rect 431316 248406 431368 248412
rect 433708 248464 433760 248470
rect 433708 248406 433760 248412
rect 431328 200802 431356 248406
rect 432604 221468 432656 221474
rect 432604 221410 432656 221416
rect 432616 209098 432644 221410
rect 433996 220862 434024 260102
rect 433984 220856 434036 220862
rect 433984 220798 434036 220804
rect 432604 209092 432656 209098
rect 432604 209034 432656 209040
rect 431316 200796 431368 200802
rect 431316 200738 431368 200744
rect 431224 161764 431276 161770
rect 431224 161706 431276 161712
rect 431236 161474 431264 161706
rect 431236 161446 431356 161474
rect 428004 160268 428056 160274
rect 428004 160210 428056 160216
rect 428648 160268 428700 160274
rect 428648 160210 428700 160216
rect 425014 160132 425066 160138
rect 425014 160074 425066 160080
rect 426348 160132 426400 160138
rect 426348 160074 426400 160080
rect 425026 159868 425054 160074
rect 428016 159882 428044 160210
rect 428660 159882 428688 160210
rect 428016 159854 428688 159882
rect 431328 159882 431356 161446
rect 436020 160342 436048 328442
rect 436756 183530 436784 331298
rect 436848 307766 436876 358770
rect 439504 335368 439556 335374
rect 439504 335310 439556 335316
rect 437020 334416 437072 334422
rect 437020 334358 437072 334364
rect 437032 328438 437060 334358
rect 438768 329112 438820 329118
rect 438768 329054 438820 329060
rect 436928 328432 436980 328438
rect 436928 328374 436980 328380
rect 437020 328432 437072 328438
rect 437020 328374 437072 328380
rect 436940 325038 436968 328374
rect 436928 325032 436980 325038
rect 436928 324974 436980 324980
rect 436836 307760 436888 307766
rect 436836 307702 436888 307708
rect 436744 183524 436796 183530
rect 436744 183466 436796 183472
rect 438780 161566 438808 329054
rect 439516 249762 439544 335310
rect 439608 318170 439636 360198
rect 441068 358896 441120 358902
rect 441068 358838 441120 358844
rect 439780 336796 439832 336802
rect 439780 336738 439832 336744
rect 440976 336796 441028 336802
rect 440976 336738 441028 336744
rect 439688 336252 439740 336258
rect 439688 336194 439740 336200
rect 439700 322046 439728 336194
rect 439792 327078 439820 336738
rect 440884 332716 440936 332722
rect 440884 332658 440936 332664
rect 440148 330608 440200 330614
rect 440148 330550 440200 330556
rect 439780 327072 439832 327078
rect 439780 327014 439832 327020
rect 439688 322040 439740 322046
rect 439688 321982 439740 321988
rect 439596 318164 439648 318170
rect 439596 318106 439648 318112
rect 439504 249756 439556 249762
rect 439504 249698 439556 249704
rect 438768 161560 438820 161566
rect 438768 161502 438820 161508
rect 438780 161474 438808 161502
rect 438596 161446 438808 161474
rect 435272 160336 435324 160342
rect 435272 160278 435324 160284
rect 436008 160336 436060 160342
rect 436008 160278 436060 160284
rect 431638 160132 431690 160138
rect 431638 160074 431690 160080
rect 431650 159882 431678 160074
rect 435284 159882 435312 160278
rect 438596 159882 438624 161446
rect 440160 161430 440188 330550
rect 440332 326392 440384 326398
rect 440332 326334 440384 326340
rect 440240 325032 440292 325038
rect 440240 324974 440292 324980
rect 440252 323678 440280 324974
rect 440240 323672 440292 323678
rect 440240 323614 440292 323620
rect 440344 316034 440372 326334
rect 440252 316006 440372 316034
rect 440252 305794 440280 316006
rect 440240 305788 440292 305794
rect 440240 305730 440292 305736
rect 440896 205630 440924 332658
rect 440988 260846 441016 336738
rect 441080 330274 441108 358838
rect 442276 348430 442304 362986
rect 442448 360324 442500 360330
rect 442448 360266 442500 360272
rect 442264 348424 442316 348430
rect 442264 348366 442316 348372
rect 442356 339584 442408 339590
rect 442356 339526 442408 339532
rect 442264 335504 442316 335510
rect 442264 335446 442316 335452
rect 442172 335096 442224 335102
rect 442172 335038 442224 335044
rect 441068 330268 441120 330274
rect 441068 330210 441120 330216
rect 442184 321842 442212 335038
rect 442172 321836 442224 321842
rect 442172 321778 442224 321784
rect 441068 288992 441120 288998
rect 441068 288934 441120 288940
rect 440976 260840 441028 260846
rect 440976 260782 441028 260788
rect 441080 255338 441108 288934
rect 441068 255332 441120 255338
rect 441068 255274 441120 255280
rect 442276 238746 442304 335446
rect 442368 304978 442396 339526
rect 442460 331906 442488 360266
rect 442540 336320 442592 336326
rect 442540 336262 442592 336268
rect 442448 331900 442500 331906
rect 442448 331842 442500 331848
rect 442552 320686 442580 336262
rect 442632 336184 442684 336190
rect 442632 336126 442684 336132
rect 442644 320754 442672 336126
rect 442724 336116 442776 336122
rect 442724 336058 442776 336064
rect 442736 321609 442764 336058
rect 442828 322454 442856 387087
rect 443656 368490 443684 418746
rect 444012 369912 444064 369918
rect 444012 369854 444064 369860
rect 443644 368484 443696 368490
rect 443644 368426 443696 368432
rect 444024 365702 444052 369854
rect 444012 365696 444064 365702
rect 444012 365638 444064 365644
rect 443644 361684 443696 361690
rect 443644 361626 443696 361632
rect 443656 344350 443684 361626
rect 443644 344344 443696 344350
rect 443644 344286 443696 344292
rect 444104 341012 444156 341018
rect 444104 340954 444156 340960
rect 443828 336864 443880 336870
rect 443828 336806 443880 336812
rect 443736 334076 443788 334082
rect 443736 334018 443788 334024
rect 443644 331288 443696 331294
rect 443644 331230 443696 331236
rect 442908 330132 442960 330138
rect 442908 330074 442960 330080
rect 442816 322448 442868 322454
rect 442816 322390 442868 322396
rect 442722 321600 442778 321609
rect 442722 321535 442778 321544
rect 442632 320748 442684 320754
rect 442632 320690 442684 320696
rect 442540 320680 442592 320686
rect 442540 320622 442592 320628
rect 442356 304972 442408 304978
rect 442356 304914 442408 304920
rect 442264 238740 442316 238746
rect 442264 238682 442316 238688
rect 440884 205624 440936 205630
rect 440884 205566 440936 205572
rect 442920 161498 442948 330074
rect 443656 171834 443684 331230
rect 443748 227730 443776 334018
rect 443840 291718 443868 336806
rect 444116 336054 444144 340954
rect 444104 336048 444156 336054
rect 444104 335990 444156 335996
rect 444208 319870 444236 422039
rect 444196 319864 444248 319870
rect 444196 319806 444248 319812
rect 444300 318782 444328 422198
rect 444392 421841 444420 422266
rect 444378 421832 444434 421841
rect 444378 421767 444434 421776
rect 444932 335028 444984 335034
rect 444932 334970 444984 334976
rect 444944 322114 444972 334970
rect 444932 322108 444984 322114
rect 444932 322050 444984 322056
rect 445036 321298 445064 700810
rect 445116 700732 445168 700738
rect 445116 700674 445168 700680
rect 445024 321292 445076 321298
rect 445024 321234 445076 321240
rect 445128 320958 445156 700674
rect 446404 700324 446456 700330
rect 446404 700266 446456 700272
rect 445208 686588 445260 686594
rect 445208 686530 445260 686536
rect 445116 320952 445168 320958
rect 445116 320894 445168 320900
rect 445220 319462 445248 686530
rect 445300 686520 445352 686526
rect 445300 686462 445352 686468
rect 445312 319598 445340 686462
rect 445392 684548 445444 684554
rect 445392 684490 445444 684496
rect 445300 319592 445352 319598
rect 445300 319534 445352 319540
rect 445404 319530 445432 684490
rect 445666 683360 445722 683369
rect 445484 683324 445536 683330
rect 445666 683295 445722 683304
rect 445484 683266 445536 683272
rect 445496 321366 445524 683266
rect 445576 683256 445628 683262
rect 445576 683198 445628 683204
rect 445484 321360 445536 321366
rect 445484 321302 445536 321308
rect 445588 321094 445616 683198
rect 445680 322182 445708 683295
rect 445760 444576 445812 444582
rect 445760 444518 445812 444524
rect 445772 329118 445800 444518
rect 445852 444508 445904 444514
rect 445852 444450 445904 444456
rect 445864 330138 445892 444450
rect 445944 444440 445996 444446
rect 445944 444382 445996 444388
rect 445956 331226 445984 444382
rect 445944 331220 445996 331226
rect 445944 331162 445996 331168
rect 445956 330614 445984 331162
rect 445944 330608 445996 330614
rect 445944 330550 445996 330556
rect 445852 330132 445904 330138
rect 445852 330074 445904 330080
rect 445760 329112 445812 329118
rect 445760 329054 445812 329060
rect 445668 322176 445720 322182
rect 445668 322118 445720 322124
rect 446416 321230 446444 700266
rect 446404 321224 446456 321230
rect 446404 321166 446456 321172
rect 445576 321088 445628 321094
rect 445576 321030 445628 321036
rect 446508 320822 446536 700878
rect 446588 700800 446640 700806
rect 446588 700742 446640 700748
rect 446600 322386 446628 700742
rect 450544 700596 450596 700602
rect 450544 700538 450596 700544
rect 447784 700324 447836 700330
rect 447784 700266 447836 700272
rect 446680 685228 446732 685234
rect 446680 685170 446732 685176
rect 446588 322380 446640 322386
rect 446588 322322 446640 322328
rect 446496 320816 446548 320822
rect 446496 320758 446548 320764
rect 446692 319734 446720 685170
rect 446772 683188 446824 683194
rect 446772 683130 446824 683136
rect 446784 321910 446812 683130
rect 446864 447228 446916 447234
rect 446864 447170 446916 447176
rect 446876 349110 446904 447170
rect 447796 423434 447824 700266
rect 450358 683224 450414 683233
rect 450358 683159 450414 683168
rect 448060 526448 448112 526454
rect 448060 526390 448112 526396
rect 447968 519580 448020 519586
rect 447968 519522 448020 519528
rect 447980 503713 448008 519522
rect 448072 514185 448100 526390
rect 448428 523728 448480 523734
rect 448428 523670 448480 523676
rect 448336 522300 448388 522306
rect 448336 522242 448388 522248
rect 448150 516760 448206 516769
rect 448150 516695 448206 516704
rect 448058 514176 448114 514185
rect 448058 514111 448114 514120
rect 448164 509234 448192 516695
rect 448348 512825 448376 522242
rect 448440 516225 448468 523670
rect 449716 520940 449768 520946
rect 449716 520882 449768 520888
rect 448426 516216 448482 516225
rect 448426 516151 448482 516160
rect 448428 516112 448480 516118
rect 448428 516054 448480 516060
rect 448334 512816 448390 512825
rect 448334 512751 448390 512760
rect 448242 510504 448298 510513
rect 448242 510439 448298 510448
rect 448072 509206 448192 509234
rect 448072 507793 448100 509206
rect 448058 507784 448114 507793
rect 448058 507719 448114 507728
rect 447966 503704 448022 503713
rect 447966 503639 448022 503648
rect 447876 444372 447928 444378
rect 447876 444314 447928 444320
rect 447784 423428 447836 423434
rect 447784 423370 447836 423376
rect 447888 386646 447916 444314
rect 447876 386640 447928 386646
rect 447876 386582 447928 386588
rect 447784 386028 447836 386034
rect 447784 385970 447836 385976
rect 447600 385416 447652 385422
rect 447600 385358 447652 385364
rect 447140 385008 447192 385014
rect 447140 384950 447192 384956
rect 447152 383897 447180 384950
rect 447138 383888 447194 383897
rect 447138 383823 447194 383832
rect 447140 383648 447192 383654
rect 447140 383590 447192 383596
rect 447152 383217 447180 383590
rect 447232 383580 447284 383586
rect 447232 383522 447284 383528
rect 447138 383208 447194 383217
rect 447138 383143 447194 383152
rect 447244 382537 447272 383522
rect 447230 382528 447286 382537
rect 447230 382463 447286 382472
rect 447140 382220 447192 382226
rect 447140 382162 447192 382168
rect 447152 381857 447180 382162
rect 447232 382152 447284 382158
rect 447232 382094 447284 382100
rect 447138 381848 447194 381857
rect 447138 381783 447194 381792
rect 447244 381177 447272 382094
rect 447230 381168 447286 381177
rect 447230 381103 447286 381112
rect 447140 380860 447192 380866
rect 447140 380802 447192 380808
rect 447152 380497 447180 380802
rect 447232 380792 447284 380798
rect 447232 380734 447284 380740
rect 447138 380488 447194 380497
rect 447138 380423 447194 380432
rect 447244 379817 447272 380734
rect 447230 379808 447286 379817
rect 447230 379743 447286 379752
rect 447232 379500 447284 379506
rect 447232 379442 447284 379448
rect 447140 379432 447192 379438
rect 447140 379374 447192 379380
rect 447152 379137 447180 379374
rect 447138 379128 447194 379137
rect 447138 379063 447194 379072
rect 447244 378457 447272 379442
rect 447230 378448 447286 378457
rect 447230 378383 447286 378392
rect 447232 378140 447284 378146
rect 447232 378082 447284 378088
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377777 447180 378014
rect 447138 377768 447194 377777
rect 447138 377703 447194 377712
rect 447244 377097 447272 378082
rect 447230 377088 447286 377097
rect 447230 377023 447286 377032
rect 447232 376712 447284 376718
rect 447232 376654 447284 376660
rect 447140 376644 447192 376650
rect 447140 376586 447192 376592
rect 447152 376417 447180 376586
rect 447138 376408 447194 376417
rect 447138 376343 447194 376352
rect 447244 375737 447272 376654
rect 447230 375728 447286 375737
rect 447230 375663 447286 375672
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 375057 447180 375294
rect 447232 375284 447284 375290
rect 447232 375226 447284 375232
rect 447138 375048 447194 375057
rect 447138 374983 447194 374992
rect 447244 374377 447272 375226
rect 447230 374368 447286 374377
rect 447230 374303 447286 374312
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373697 447180 373934
rect 447232 373924 447284 373930
rect 447232 373866 447284 373872
rect 447138 373688 447194 373697
rect 447138 373623 447194 373632
rect 447244 373017 447272 373866
rect 447230 373008 447286 373017
rect 447230 372943 447286 372952
rect 447140 372564 447192 372570
rect 447140 372506 447192 372512
rect 447152 372337 447180 372506
rect 447232 372496 447284 372502
rect 447232 372438 447284 372444
rect 447138 372328 447194 372337
rect 447138 372263 447194 372272
rect 447244 371657 447272 372438
rect 447230 371648 447286 371657
rect 447230 371583 447286 371592
rect 447232 371204 447284 371210
rect 447232 371146 447284 371152
rect 447140 371136 447192 371142
rect 447140 371078 447192 371084
rect 447152 370977 447180 371078
rect 447138 370968 447194 370977
rect 447138 370903 447194 370912
rect 447244 370297 447272 371146
rect 447230 370288 447286 370297
rect 447230 370223 447286 370232
rect 447232 369844 447284 369850
rect 447232 369786 447284 369792
rect 447140 369776 447192 369782
rect 447140 369718 447192 369724
rect 447152 369617 447180 369718
rect 447138 369608 447194 369617
rect 447138 369543 447194 369552
rect 447244 368937 447272 369786
rect 447230 368928 447286 368937
rect 447230 368863 447286 368872
rect 447140 368484 447192 368490
rect 447140 368426 447192 368432
rect 447152 368257 447180 368426
rect 447232 368416 447284 368422
rect 447232 368358 447284 368364
rect 447138 368248 447194 368257
rect 447138 368183 447194 368192
rect 447244 367577 447272 368358
rect 447230 367568 447286 367577
rect 447230 367503 447286 367512
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366897 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447138 366888 447194 366897
rect 447138 366823 447194 366832
rect 447244 366217 447272 366930
rect 447230 366208 447286 366217
rect 447230 366143 447286 366152
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364857 447180 365638
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447244 365537 447272 365570
rect 447230 365528 447286 365537
rect 447230 365463 447286 365472
rect 447138 364848 447194 364857
rect 447138 364783 447194 364792
rect 447138 364168 447194 364177
rect 447138 364103 447194 364112
rect 447152 362982 447180 364103
rect 447230 363488 447286 363497
rect 447230 363423 447286 363432
rect 447244 363050 447272 363423
rect 447232 363044 447284 363050
rect 447232 362986 447284 362992
rect 447140 362976 447192 362982
rect 447140 362918 447192 362924
rect 447230 362808 447286 362817
rect 447230 362743 447286 362752
rect 447138 362128 447194 362137
rect 447138 362063 447194 362072
rect 447152 361622 447180 362063
rect 447244 361690 447272 362743
rect 447232 361684 447284 361690
rect 447232 361626 447284 361632
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447230 361448 447286 361457
rect 447230 361383 447286 361392
rect 447138 360768 447194 360777
rect 447138 360703 447194 360712
rect 447152 360262 447180 360703
rect 447244 360330 447272 361383
rect 447232 360324 447284 360330
rect 447232 360266 447284 360272
rect 447140 360256 447192 360262
rect 447140 360198 447192 360204
rect 447230 360088 447286 360097
rect 447230 360023 447286 360032
rect 447138 359408 447194 359417
rect 447138 359343 447194 359352
rect 447152 358834 447180 359343
rect 447244 358902 447272 360023
rect 447232 358896 447284 358902
rect 447232 358838 447284 358844
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447612 352617 447640 385358
rect 447692 385144 447744 385150
rect 447692 385086 447744 385092
rect 447598 352608 447654 352617
rect 447598 352543 447654 352552
rect 447140 351960 447192 351966
rect 447138 351928 447140 351937
rect 447192 351928 447194 351937
rect 447138 351863 447194 351872
rect 447414 351248 447470 351257
rect 447414 351183 447470 351192
rect 447140 350600 447192 350606
rect 447138 350568 447140 350577
rect 447192 350568 447194 350577
rect 447138 350503 447194 350512
rect 446864 349104 446916 349110
rect 446864 349046 446916 349052
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347177 447180 347686
rect 447138 347168 447194 347177
rect 447138 347103 447194 347112
rect 447322 343768 447378 343777
rect 447322 343703 447378 343712
rect 447138 341728 447194 341737
rect 447138 341663 447194 341672
rect 447152 340950 447180 341663
rect 447230 341048 447286 341057
rect 447230 340983 447232 340992
rect 447284 340983 447286 340992
rect 447232 340954 447284 340960
rect 447140 340944 447192 340950
rect 447140 340886 447192 340892
rect 447138 340368 447194 340377
rect 447138 340303 447194 340312
rect 447152 339522 447180 340303
rect 447230 339688 447286 339697
rect 447230 339623 447286 339632
rect 447244 339590 447272 339623
rect 447232 339584 447284 339590
rect 447232 339526 447284 339532
rect 447140 339516 447192 339522
rect 447140 339458 447192 339464
rect 447230 339008 447286 339017
rect 447230 338943 447286 338952
rect 447138 338328 447194 338337
rect 447138 338263 447194 338272
rect 447152 338230 447180 338263
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 338943
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447230 337648 447286 337657
rect 447230 337583 447286 337592
rect 447138 336968 447194 336977
rect 447138 336903 447194 336912
rect 447152 336802 447180 336903
rect 447244 336870 447272 337583
rect 447232 336864 447284 336870
rect 447232 336806 447284 336812
rect 447140 336796 447192 336802
rect 447140 336738 447192 336744
rect 447336 336682 447364 343703
rect 447152 336654 447364 336682
rect 446956 334960 447008 334966
rect 446956 334902 447008 334908
rect 446864 334892 446916 334898
rect 446864 334834 446916 334840
rect 446772 321904 446824 321910
rect 446772 321846 446824 321852
rect 446876 320006 446904 334834
rect 446968 322318 446996 334902
rect 446956 322312 447008 322318
rect 446956 322254 447008 322260
rect 446864 320000 446916 320006
rect 446864 319942 446916 319948
rect 446680 319728 446732 319734
rect 446680 319670 446732 319676
rect 445392 319524 445444 319530
rect 445392 319466 445444 319472
rect 445208 319456 445260 319462
rect 445208 319398 445260 319404
rect 444288 318776 444340 318782
rect 444288 318718 444340 318724
rect 446404 308508 446456 308514
rect 446404 308450 446456 308456
rect 443828 291712 443880 291718
rect 443828 291654 443880 291660
rect 446416 288998 446444 308450
rect 446404 288992 446456 288998
rect 446404 288934 446456 288940
rect 445024 281920 445076 281926
rect 445024 281862 445076 281868
rect 443828 274712 443880 274718
rect 443828 274654 443880 274660
rect 443840 260166 443868 274654
rect 445036 272542 445064 281862
rect 445024 272536 445076 272542
rect 445024 272478 445076 272484
rect 445024 268524 445076 268530
rect 445024 268466 445076 268472
rect 443828 260160 443880 260166
rect 443828 260102 443880 260108
rect 443736 227724 443788 227730
rect 443736 227666 443788 227672
rect 445036 213246 445064 268466
rect 446404 249076 446456 249082
rect 446404 249018 446456 249024
rect 445024 213240 445076 213246
rect 445024 213182 445076 213188
rect 443644 171828 443696 171834
rect 443644 171770 443696 171776
rect 446416 163538 446444 249018
rect 445668 163532 445720 163538
rect 445668 163474 445720 163480
rect 446404 163532 446456 163538
rect 446404 163474 446456 163480
rect 441620 161492 441672 161498
rect 441620 161434 441672 161440
rect 442908 161492 442960 161498
rect 442908 161434 442960 161440
rect 440148 161424 440200 161430
rect 440148 161366 440200 161372
rect 440160 160750 440188 161366
rect 440148 160744 440200 160750
rect 440148 160686 440200 160692
rect 441632 160154 441660 161434
rect 445680 160206 445708 163474
rect 447152 161474 447180 336654
rect 447230 336288 447286 336297
rect 447230 336223 447286 336232
rect 447244 335374 447272 336223
rect 447322 335608 447378 335617
rect 447322 335543 447378 335552
rect 447336 335510 447364 335543
rect 447324 335504 447376 335510
rect 447324 335446 447376 335452
rect 447232 335368 447284 335374
rect 447232 335310 447284 335316
rect 447322 334928 447378 334937
rect 447322 334863 447378 334872
rect 447230 334248 447286 334257
rect 447230 334183 447286 334192
rect 447244 334014 447272 334183
rect 447336 334082 447364 334863
rect 447324 334076 447376 334082
rect 447324 334018 447376 334024
rect 447232 334008 447284 334014
rect 447232 333950 447284 333956
rect 447322 333568 447378 333577
rect 447322 333503 447378 333512
rect 447230 332888 447286 332897
rect 447230 332823 447286 332832
rect 447244 332654 447272 332823
rect 447336 332722 447364 333503
rect 447324 332716 447376 332722
rect 447324 332658 447376 332664
rect 447232 332648 447284 332654
rect 447232 332590 447284 332596
rect 447230 331528 447286 331537
rect 447230 331463 447286 331472
rect 447244 331294 447272 331463
rect 447232 331288 447284 331294
rect 447232 331230 447284 331236
rect 447324 331220 447376 331226
rect 447324 331162 447376 331168
rect 447336 330857 447364 331162
rect 447322 330848 447378 330857
rect 447322 330783 447378 330792
rect 447230 330168 447286 330177
rect 447230 330103 447232 330112
rect 447284 330103 447286 330112
rect 447232 330074 447284 330080
rect 447230 329488 447286 329497
rect 447230 329423 447286 329432
rect 447244 329118 447272 329423
rect 447232 329112 447284 329118
rect 447232 329054 447284 329060
rect 447230 328808 447286 328817
rect 447230 328743 447286 328752
rect 447244 328506 447272 328743
rect 447232 328500 447284 328506
rect 447232 328442 447284 328448
rect 447324 328432 447376 328438
rect 447324 328374 447376 328380
rect 447230 328128 447286 328137
rect 447230 328063 447286 328072
rect 447244 327146 447272 328063
rect 447336 327457 447364 328374
rect 447322 327448 447378 327457
rect 447322 327383 447378 327392
rect 447232 327140 447284 327146
rect 447232 327082 447284 327088
rect 447324 327072 447376 327078
rect 447324 327014 447376 327020
rect 447230 326768 447286 326777
rect 447230 326703 447286 326712
rect 447244 326398 447272 326703
rect 447232 326392 447284 326398
rect 447232 326334 447284 326340
rect 447336 326097 447364 327014
rect 447322 326088 447378 326097
rect 447322 326023 447378 326032
rect 447232 323672 447284 323678
rect 447232 323614 447284 323620
rect 447244 322250 447272 323614
rect 447232 322244 447284 322250
rect 447232 322186 447284 322192
rect 447428 163606 447456 351183
rect 447600 349104 447652 349110
rect 447600 349046 447652 349052
rect 447612 344457 447640 349046
rect 447704 347857 447732 385086
rect 447796 348537 447824 385970
rect 447782 348528 447838 348537
rect 447782 348463 447838 348472
rect 447690 347848 447746 347857
rect 447690 347783 447746 347792
rect 447598 344448 447654 344457
rect 447598 344383 447654 344392
rect 447888 343097 447916 386582
rect 447874 343088 447930 343097
rect 447874 343023 447930 343032
rect 447888 342922 447916 343023
rect 447876 342916 447928 342922
rect 447876 342858 447928 342864
rect 447506 332208 447562 332217
rect 447506 332143 447562 332152
rect 447520 331362 447548 332143
rect 447508 331356 447560 331362
rect 447508 331298 447560 331304
rect 447416 163600 447468 163606
rect 447416 163542 447468 163548
rect 447520 163538 447548 331298
rect 447980 325514 448008 503639
rect 448072 327078 448100 507719
rect 448150 505200 448206 505209
rect 448150 505135 448206 505144
rect 448060 327072 448112 327078
rect 448060 327014 448112 327020
rect 448164 325650 448192 505135
rect 448256 326777 448284 510439
rect 448348 498794 448376 512751
rect 448440 510513 448468 516054
rect 448426 510504 448482 510513
rect 448426 510439 448482 510448
rect 449728 505685 449756 520882
rect 449808 518220 449860 518226
rect 449808 518162 449860 518168
rect 449714 505676 449770 505685
rect 449714 505611 449770 505620
rect 449820 501333 449848 518162
rect 449806 501324 449862 501333
rect 449806 501259 449862 501268
rect 448518 500304 448574 500313
rect 448518 500239 448520 500248
rect 448572 500239 448574 500248
rect 448520 500210 448572 500216
rect 448520 498840 448572 498846
rect 448348 498788 448520 498794
rect 448348 498782 448572 498788
rect 448348 498766 448560 498782
rect 448348 328438 448376 498766
rect 448428 496120 448480 496126
rect 448426 496088 448428 496097
rect 448480 496088 448482 496097
rect 448426 496023 448482 496032
rect 449992 494760 450044 494766
rect 449992 494702 450044 494708
rect 449808 464364 449860 464370
rect 449808 464306 449860 464312
rect 449716 460216 449768 460222
rect 449716 460158 449768 460164
rect 449624 458856 449676 458862
rect 449624 458798 449676 458804
rect 449440 457496 449492 457502
rect 449440 457438 449492 457444
rect 449348 454708 449400 454714
rect 449348 454650 449400 454656
rect 449070 389872 449126 389881
rect 449070 389807 449126 389816
rect 448428 388476 448480 388482
rect 448428 388418 448480 388424
rect 448440 349217 448468 388418
rect 448978 387016 449034 387025
rect 448978 386951 449034 386960
rect 448992 353297 449020 386951
rect 449084 354657 449112 389807
rect 449164 387116 449216 387122
rect 449164 387058 449216 387064
rect 449070 354648 449126 354657
rect 449070 354583 449126 354592
rect 448978 353288 449034 353297
rect 448978 353223 449034 353232
rect 448426 349208 448482 349217
rect 448426 349143 448482 349152
rect 449176 342417 449204 387058
rect 449254 385656 449310 385665
rect 449254 385591 449310 385600
rect 449162 342408 449218 342417
rect 449162 342343 449218 342352
rect 449164 338768 449216 338774
rect 449164 338710 449216 338716
rect 449072 334688 449124 334694
rect 449072 334630 449124 334636
rect 448336 328432 448388 328438
rect 448336 328374 448388 328380
rect 448242 326768 448298 326777
rect 448242 326703 448298 326712
rect 448152 325644 448204 325650
rect 448152 325586 448204 325592
rect 447968 325508 448020 325514
rect 447968 325450 448020 325456
rect 447980 324737 448008 325450
rect 448164 325417 448192 325586
rect 448150 325408 448206 325417
rect 448150 325343 448206 325352
rect 448426 325408 448482 325417
rect 448426 325343 448482 325352
rect 447966 324728 448022 324737
rect 447966 324663 448022 324672
rect 447784 317008 447836 317014
rect 447784 316950 447836 316956
rect 447796 281926 447824 316950
rect 447784 281920 447836 281926
rect 447784 281862 447836 281868
rect 447980 220114 448008 324663
rect 448440 317082 448468 325343
rect 449084 319802 449112 334630
rect 449072 319796 449124 319802
rect 449072 319738 449124 319744
rect 449176 319258 449204 338710
rect 449268 324193 449296 385591
rect 449360 355337 449388 454650
rect 449452 356697 449480 457438
rect 449532 454776 449584 454782
rect 449532 454718 449584 454724
rect 449438 356688 449494 356697
rect 449438 356623 449494 356632
rect 449346 355328 449402 355337
rect 449346 355263 449402 355272
rect 449544 353977 449572 454718
rect 449636 357377 449664 458798
rect 449622 357368 449678 357377
rect 449622 357303 449678 357312
rect 449728 356017 449756 460158
rect 449714 356008 449770 356017
rect 449714 355943 449770 355952
rect 449530 353968 449586 353977
rect 449530 353903 449586 353912
rect 449714 349888 449770 349897
rect 449714 349823 449770 349832
rect 449622 343088 449678 343097
rect 449622 343023 449678 343032
rect 449440 334824 449492 334830
rect 449440 334766 449492 334772
rect 449348 334620 449400 334626
rect 449348 334562 449400 334568
rect 449254 324184 449310 324193
rect 449254 324119 449310 324128
rect 449268 323610 449296 324119
rect 449256 323604 449308 323610
rect 449256 323546 449308 323552
rect 449360 319326 449388 334562
rect 449452 319394 449480 334766
rect 449532 334756 449584 334762
rect 449532 334698 449584 334704
rect 449544 319666 449572 334698
rect 449532 319660 449584 319666
rect 449532 319602 449584 319608
rect 449440 319388 449492 319394
rect 449440 319330 449492 319336
rect 449348 319320 449400 319326
rect 449348 319262 449400 319268
rect 449164 319252 449216 319258
rect 449164 319194 449216 319200
rect 449636 318102 449664 343023
rect 449624 318096 449676 318102
rect 449624 318038 449676 318044
rect 448428 317076 448480 317082
rect 448428 317018 448480 317024
rect 449164 283620 449216 283626
rect 449164 283562 449216 283568
rect 449176 274718 449204 283562
rect 449164 274712 449216 274718
rect 449164 274654 449216 274660
rect 449728 263566 449756 349823
rect 449820 345817 449848 464306
rect 449900 460964 449952 460970
rect 449900 460906 449952 460912
rect 449912 346905 449940 460906
rect 450004 389298 450032 494702
rect 450084 391332 450136 391338
rect 450084 391274 450136 391280
rect 449992 389292 450044 389298
rect 449992 389234 450044 389240
rect 450096 358465 450124 391274
rect 450268 387184 450320 387190
rect 450268 387126 450320 387132
rect 450280 358873 450308 387126
rect 450266 358864 450322 358873
rect 450266 358799 450322 358808
rect 450082 358456 450138 358465
rect 450082 358391 450138 358400
rect 449898 346896 449954 346905
rect 449898 346831 449954 346840
rect 449806 345808 449862 345817
rect 449806 345743 449862 345752
rect 449806 345128 449862 345137
rect 449806 345063 449862 345072
rect 449820 276758 449848 345063
rect 449992 322448 450044 322454
rect 449992 322390 450044 322396
rect 450004 322250 450032 322390
rect 449900 322244 449952 322250
rect 449900 322186 449952 322192
rect 449992 322244 450044 322250
rect 449992 322186 450044 322192
rect 449912 320890 449940 322186
rect 449900 320884 449952 320890
rect 449900 320826 449952 320832
rect 450372 319977 450400 683159
rect 450452 682712 450504 682718
rect 450452 682654 450504 682660
rect 450358 319968 450414 319977
rect 450464 319938 450492 682654
rect 450556 321026 450584 700538
rect 450636 700392 450688 700398
rect 450636 700334 450688 700340
rect 450648 321978 450676 700334
rect 462332 669905 462360 703520
rect 478524 700330 478552 703520
rect 494808 700369 494836 703520
rect 494794 700360 494850 700369
rect 478512 700324 478564 700330
rect 494794 700295 494850 700304
rect 478512 700266 478564 700272
rect 527192 699825 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 462318 669896 462374 669905
rect 462318 669831 462374 669840
rect 458086 662552 458142 662561
rect 458086 662487 458142 662496
rect 457718 659968 457774 659977
rect 457718 659903 457774 659912
rect 457626 652896 457682 652905
rect 457626 652831 457682 652840
rect 457534 645960 457590 645969
rect 457534 645895 457590 645904
rect 457350 623928 457406 623937
rect 457350 623863 457406 623872
rect 457258 611416 457314 611425
rect 457258 611351 457314 611360
rect 457272 525094 457300 611351
rect 457364 600030 457392 623863
rect 457442 618352 457498 618361
rect 457442 618287 457498 618296
rect 457352 600024 457404 600030
rect 457352 599966 457404 599972
rect 457456 596222 457484 618287
rect 457548 600642 457576 645895
rect 457536 600636 457588 600642
rect 457536 600578 457588 600584
rect 457640 598262 457668 652831
rect 457732 598330 457760 659903
rect 457994 657520 458050 657529
rect 457994 657455 458050 657464
rect 457902 650176 457958 650185
rect 457902 650111 457958 650120
rect 457810 621072 457866 621081
rect 457810 621007 457866 621016
rect 457720 598324 457772 598330
rect 457720 598266 457772 598272
rect 457628 598256 457680 598262
rect 457628 598198 457680 598204
rect 457444 596216 457496 596222
rect 457444 596158 457496 596164
rect 457824 543046 457852 621007
rect 457916 599622 457944 650111
rect 457904 599616 457956 599622
rect 457904 599558 457956 599564
rect 457812 543040 457864 543046
rect 457812 542982 457864 542988
rect 457260 525088 457312 525094
rect 457260 525030 457312 525036
rect 458008 519654 458036 657455
rect 458100 521014 458128 662487
rect 459190 655752 459246 655761
rect 459190 655687 459246 655696
rect 459098 647728 459154 647737
rect 459098 647663 459154 647672
rect 459006 643240 459062 643249
rect 459006 643175 459062 643184
rect 458914 640384 458970 640393
rect 458914 640319 458970 640328
rect 458822 616040 458878 616049
rect 458822 615975 458878 615984
rect 458730 608696 458786 608705
rect 458730 608631 458786 608640
rect 458744 596970 458772 608631
rect 458836 599690 458864 615975
rect 458824 599684 458876 599690
rect 458824 599626 458876 599632
rect 458928 598233 458956 640319
rect 459020 599729 459048 643175
rect 459006 599720 459062 599729
rect 459006 599655 459062 599664
rect 459112 599593 459140 647663
rect 459098 599584 459154 599593
rect 459098 599519 459154 599528
rect 458914 598224 458970 598233
rect 458914 598159 458970 598168
rect 458732 596964 458784 596970
rect 458732 596906 458784 596912
rect 459204 595513 459232 655687
rect 459282 637936 459338 637945
rect 459282 637871 459338 637880
rect 459190 595504 459246 595513
rect 459190 595439 459246 595448
rect 459296 541657 459324 637871
rect 459374 635488 459430 635497
rect 459374 635423 459430 635432
rect 459282 541648 459338 541657
rect 459282 541583 459338 541592
rect 459388 522345 459416 635423
rect 459466 633448 459522 633457
rect 459466 633383 459522 633392
rect 459374 522336 459430 522345
rect 459374 522271 459430 522280
rect 458088 521008 458140 521014
rect 458088 520950 458140 520956
rect 457996 519648 458048 519654
rect 457996 519590 458048 519596
rect 459480 518129 459508 633383
rect 459742 628756 459798 628765
rect 459742 628691 459798 628700
rect 459558 626308 459614 626317
rect 459558 626243 459614 626252
rect 459572 541686 459600 626243
rect 459650 601896 459706 601905
rect 459650 601831 459706 601840
rect 459560 541680 459612 541686
rect 459560 541622 459612 541628
rect 459466 518120 459522 518129
rect 459466 518055 459522 518064
rect 459664 517546 459692 601831
rect 459756 596834 459784 628691
rect 459834 614136 459890 614145
rect 459834 614071 459890 614080
rect 459848 596902 459876 614071
rect 459926 606384 459982 606393
rect 459926 606319 459982 606328
rect 459940 598398 459968 606319
rect 460202 603664 460258 603673
rect 460202 603599 460258 603608
rect 460216 599826 460244 603599
rect 461584 600636 461636 600642
rect 461584 600578 461636 600584
rect 460204 599820 460256 599826
rect 460204 599762 460256 599768
rect 459928 598392 459980 598398
rect 459928 598334 459980 598340
rect 459836 596896 459888 596902
rect 459836 596838 459888 596844
rect 459744 596828 459796 596834
rect 459744 596770 459796 596776
rect 459652 517540 459704 517546
rect 459652 517482 459704 517488
rect 450740 494766 450768 500140
rect 451292 500126 452226 500154
rect 450728 494760 450780 494766
rect 450728 494702 450780 494708
rect 450728 389292 450780 389298
rect 450728 389234 450780 389240
rect 450740 385914 450768 389234
rect 451292 385914 451320 500126
rect 453304 497480 453356 497486
rect 453304 497422 453356 497428
rect 452844 496936 452896 496942
rect 452844 496878 452896 496884
rect 451372 496868 451424 496874
rect 451372 496810 451424 496816
rect 451384 402974 451412 496810
rect 451924 455524 451976 455530
rect 451924 455466 451976 455472
rect 451384 402946 451872 402974
rect 451844 385914 451872 402946
rect 451936 386034 451964 455466
rect 451924 386028 451976 386034
rect 451924 385970 451976 385976
rect 452856 385914 452884 496878
rect 450740 385886 450846 385914
rect 451292 385886 451582 385914
rect 451844 385886 452318 385914
rect 452856 385886 453054 385914
rect 453316 385422 453344 497422
rect 453684 496874 453712 500140
rect 454040 497072 454092 497078
rect 454040 497014 454092 497020
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 454052 389298 454080 497014
rect 454132 497004 454184 497010
rect 454132 496946 454184 496952
rect 454040 389292 454092 389298
rect 454040 389234 454092 389240
rect 453764 389156 453816 389162
rect 453764 389098 453816 389104
rect 453776 385900 453804 389098
rect 454144 385914 454172 496946
rect 455156 496942 455184 500140
rect 455144 496936 455196 496942
rect 455144 496878 455196 496884
rect 455420 496936 455472 496942
rect 455420 496878 455472 496884
rect 454684 496868 454736 496874
rect 454684 496810 454736 496816
rect 454696 389162 454724 496810
rect 455432 402974 455460 496878
rect 456628 496874 456656 500140
rect 458100 497010 458128 500140
rect 459572 497078 459600 500140
rect 459560 497072 459612 497078
rect 459560 497014 459612 497020
rect 458088 497004 458140 497010
rect 458088 496946 458140 496952
rect 461044 496942 461072 500140
rect 461032 496936 461084 496942
rect 461032 496878 461084 496884
rect 456616 496868 456668 496874
rect 456616 496810 456668 496816
rect 456892 430024 456944 430030
rect 456892 429966 456944 429972
rect 456904 402974 456932 429966
rect 458180 429956 458232 429962
rect 458180 429898 458232 429904
rect 457444 428460 457496 428466
rect 457444 428402 457496 428408
rect 455432 402946 455552 402974
rect 456904 402946 457024 402974
rect 454868 389292 454920 389298
rect 454868 389234 454920 389240
rect 454684 389156 454736 389162
rect 454684 389098 454736 389104
rect 454880 385914 454908 389234
rect 455524 385914 455552 402946
rect 456708 389156 456760 389162
rect 456708 389098 456760 389104
rect 454144 385886 454526 385914
rect 454880 385886 455262 385914
rect 455524 385886 455998 385914
rect 456720 385900 456748 389098
rect 456996 385914 457024 402946
rect 457456 389162 457484 428402
rect 457444 389156 457496 389162
rect 457444 389098 457496 389104
rect 456996 385886 457470 385914
rect 458192 385900 458220 429898
rect 458364 429888 458416 429894
rect 458364 429830 458416 429836
rect 458376 402974 458404 429830
rect 458376 402946 458496 402974
rect 458468 385914 458496 402946
rect 460940 395344 460992 395350
rect 460940 395286 460992 395292
rect 460388 389904 460440 389910
rect 460388 389846 460440 389852
rect 459652 388748 459704 388754
rect 459652 388690 459704 388696
rect 458468 385886 458942 385914
rect 459664 385900 459692 388690
rect 460400 385900 460428 389846
rect 460952 389298 460980 395286
rect 461032 393984 461084 393990
rect 461032 393926 461084 393932
rect 460940 389292 460992 389298
rect 460940 389234 460992 389240
rect 461044 385914 461072 393926
rect 461492 389292 461544 389298
rect 461492 389234 461544 389240
rect 461504 385914 461532 389234
rect 461596 388618 461624 600578
rect 462424 600086 463266 600114
rect 469232 600086 469614 600114
rect 474752 600086 475962 600114
rect 461676 596216 461728 596222
rect 461676 596158 461728 596164
rect 461688 388686 461716 596158
rect 462318 563000 462374 563009
rect 462318 562935 462374 562944
rect 461768 520464 461820 520470
rect 461768 520406 461820 520412
rect 461676 388680 461728 388686
rect 461676 388622 461728 388628
rect 461584 388612 461636 388618
rect 461584 388554 461636 388560
rect 461780 388482 461808 520406
rect 461768 388476 461820 388482
rect 461768 388418 461820 388424
rect 462332 385914 462360 562935
rect 462424 518226 462452 600086
rect 462964 600024 463016 600030
rect 462964 599966 463016 599972
rect 462412 518220 462464 518226
rect 462412 518162 462464 518168
rect 462504 517540 462556 517546
rect 462504 517482 462556 517488
rect 462516 402974 462544 517482
rect 462516 402946 462912 402974
rect 462884 385914 462912 402946
rect 462976 388210 463004 599966
rect 463700 599820 463752 599826
rect 463700 599762 463752 599768
rect 463608 392624 463660 392630
rect 463608 392566 463660 392572
rect 463620 388754 463648 392566
rect 463608 388748 463660 388754
rect 463608 388690 463660 388696
rect 462964 388204 463016 388210
rect 462964 388146 463016 388152
rect 463712 385914 463740 599762
rect 466460 599684 466512 599690
rect 466460 599626 466512 599632
rect 463792 598392 463844 598398
rect 463792 598334 463844 598340
rect 463804 402974 463832 598334
rect 464344 598324 464396 598330
rect 464344 598266 464396 598272
rect 463804 402946 464292 402974
rect 464264 386050 464292 402946
rect 464356 388482 464384 598266
rect 465080 596964 465132 596970
rect 465080 596906 465132 596912
rect 464344 388476 464396 388482
rect 464344 388418 464396 388424
rect 464264 386022 464384 386050
rect 464356 385914 464384 386022
rect 465092 385914 465120 596906
rect 465172 525088 465224 525094
rect 465172 525030 465224 525036
rect 465184 402974 465212 525030
rect 465724 521008 465776 521014
rect 465724 520950 465776 520956
rect 465184 402946 465672 402974
rect 465644 386050 465672 402946
rect 465736 388550 465764 520950
rect 465724 388544 465776 388550
rect 465724 388486 465776 388492
rect 466472 387802 466500 599626
rect 468484 598256 468536 598262
rect 469232 598210 469260 600086
rect 469864 599616 469916 599622
rect 469864 599558 469916 599564
rect 468484 598198 468536 598204
rect 466552 596896 466604 596902
rect 466552 596838 466604 596844
rect 466460 387796 466512 387802
rect 466460 387738 466512 387744
rect 465644 386022 465856 386050
rect 465828 385914 465856 386022
rect 466564 385914 466592 596838
rect 467840 520396 467892 520402
rect 467840 520338 467892 520344
rect 467852 519586 467880 520338
rect 467840 519580 467892 519586
rect 467840 519522 467892 519528
rect 468496 388822 468524 598198
rect 469140 598182 469260 598210
rect 468576 543040 468628 543046
rect 468576 542982 468628 542988
rect 468588 389162 468616 542982
rect 468666 523696 468722 523705
rect 468666 523631 468722 523640
rect 468576 389156 468628 389162
rect 468576 389098 468628 389104
rect 468484 388816 468536 388822
rect 468484 388758 468536 388764
rect 468680 388686 468708 523631
rect 469140 520402 469168 598182
rect 469128 520396 469180 520402
rect 469128 520338 469180 520344
rect 468760 519648 468812 519654
rect 468760 519590 468812 519596
rect 468772 388754 468800 519590
rect 469220 389156 469272 389162
rect 469220 389098 469272 389104
rect 468760 388748 468812 388754
rect 468760 388690 468812 388696
rect 468484 388680 468536 388686
rect 468484 388622 468536 388628
rect 468668 388680 468720 388686
rect 468668 388622 468720 388628
rect 467380 387796 467432 387802
rect 467380 387738 467432 387744
rect 467392 385914 467420 387738
rect 461044 385886 461150 385914
rect 461504 385886 461886 385914
rect 462332 385886 462622 385914
rect 462884 385886 463358 385914
rect 463712 385886 464094 385914
rect 464356 385886 464830 385914
rect 465092 385886 465566 385914
rect 465828 385886 466302 385914
rect 466564 385886 467038 385914
rect 467392 385886 467774 385914
rect 468496 385900 468524 388622
rect 469232 385900 469260 389098
rect 469876 388958 469904 599558
rect 470876 596828 470928 596834
rect 470876 596770 470928 596776
rect 470692 541680 470744 541686
rect 470692 541622 470744 541628
rect 469864 388952 469916 388958
rect 469864 388894 469916 388900
rect 469956 388204 470008 388210
rect 469956 388146 470008 388152
rect 469968 385900 469996 388146
rect 470704 385900 470732 541622
rect 470888 402974 470916 596770
rect 474752 521694 474780 600086
rect 482296 598262 482324 600100
rect 488644 598330 488672 600100
rect 488632 598324 488684 598330
rect 488632 598266 488684 598272
rect 494244 598324 494296 598330
rect 494244 598266 494296 598272
rect 482284 598256 482336 598262
rect 482284 598198 482336 598204
rect 494060 598256 494112 598262
rect 494060 598198 494112 598204
rect 493324 597916 493376 597922
rect 493324 597858 493376 597864
rect 493336 522306 493364 597858
rect 493324 522300 493376 522306
rect 493324 522242 493376 522248
rect 474740 521688 474792 521694
rect 474740 521630 474792 521636
rect 475200 521688 475252 521694
rect 475200 521630 475252 521636
rect 475212 520946 475240 521630
rect 475200 520940 475252 520946
rect 475200 520882 475252 520888
rect 482652 520940 482704 520946
rect 482652 520882 482704 520888
rect 482664 520334 482692 520882
rect 488632 520464 488684 520470
rect 488632 520406 488684 520412
rect 477408 520328 477460 520334
rect 477408 520270 477460 520276
rect 482652 520328 482704 520334
rect 482652 520270 482704 520276
rect 477420 461650 477448 520270
rect 482664 517970 482692 520270
rect 488644 517970 488672 520406
rect 482664 517942 483000 517970
rect 488644 517942 488980 517970
rect 494072 516769 494100 598198
rect 494256 586514 494284 598266
rect 494992 597922 495020 600100
rect 500972 600086 501354 600114
rect 506492 600086 507702 600114
rect 513392 600086 514050 600114
rect 520292 600086 520398 600114
rect 525812 600086 526746 600114
rect 494980 597916 495032 597922
rect 494980 597858 495032 597864
rect 494164 586486 494284 586514
rect 494058 516760 494114 516769
rect 494058 516695 494114 516704
rect 491850 516216 491906 516225
rect 491850 516151 491852 516160
rect 491904 516151 491906 516160
rect 491852 516122 491904 516128
rect 494058 515944 494114 515953
rect 494164 515930 494192 586486
rect 500972 526454 501000 600086
rect 500960 526448 501012 526454
rect 500960 526390 501012 526396
rect 506492 523734 506520 600086
rect 511264 576904 511316 576910
rect 511264 576846 511316 576852
rect 506480 523728 506532 523734
rect 506480 523670 506532 523676
rect 494336 521688 494388 521694
rect 494336 521630 494388 521636
rect 494244 520396 494296 520402
rect 494244 520338 494296 520344
rect 494114 515902 494192 515930
rect 494058 515879 494114 515888
rect 494072 515438 494100 515879
rect 494060 515432 494112 515438
rect 494060 515374 494112 515380
rect 494060 512644 494112 512650
rect 494060 512586 494112 512592
rect 494072 512553 494100 512586
rect 494058 512544 494114 512553
rect 494058 512479 494114 512488
rect 494256 505753 494284 520338
rect 494348 508881 494376 521630
rect 494426 516760 494482 516769
rect 494426 516695 494482 516704
rect 494440 512650 494468 516695
rect 494428 512644 494480 512650
rect 494428 512586 494480 512592
rect 494334 508872 494390 508881
rect 494334 508807 494390 508816
rect 494348 508570 494376 508807
rect 494336 508564 494388 508570
rect 494336 508506 494388 508512
rect 495072 505776 495124 505782
rect 494242 505744 494298 505753
rect 494242 505679 494298 505688
rect 495070 505744 495072 505753
rect 495124 505744 495126 505753
rect 495070 505679 495126 505688
rect 494058 501256 494114 501265
rect 494058 501191 494114 501200
rect 480272 500126 480608 500154
rect 480272 497486 480300 500126
rect 481790 499882 481818 500140
rect 482112 500126 483000 500154
rect 483860 500126 484196 500154
rect 484412 500126 485392 500154
rect 485792 500126 486588 500154
rect 487172 500126 487784 500154
rect 488552 500126 488980 500154
rect 490176 500126 491156 500154
rect 481790 499854 481864 499882
rect 480260 497480 480312 497486
rect 480260 497422 480312 497428
rect 481836 496913 481864 499854
rect 481822 496904 481878 496913
rect 481822 496839 481878 496848
rect 482112 489914 482140 500126
rect 483860 496913 483888 500126
rect 483846 496904 483902 496913
rect 483846 496839 483902 496848
rect 481652 489886 482140 489914
rect 477408 461644 477460 461650
rect 477408 461586 477460 461592
rect 477420 461514 477448 461586
rect 476028 461508 476080 461514
rect 476028 461450 476080 461456
rect 477408 461508 477460 461514
rect 477408 461450 477460 461456
rect 476040 456550 476068 461450
rect 473728 456544 473780 456550
rect 473728 456486 473780 456492
rect 476028 456544 476080 456550
rect 476028 456486 476080 456492
rect 473740 455462 473768 456486
rect 480996 455524 481048 455530
rect 480996 455466 481048 455472
rect 473728 455456 473780 455462
rect 473728 455398 473780 455404
rect 473740 453900 473768 455398
rect 481008 453900 481036 455466
rect 481652 454782 481680 489886
rect 481640 454776 481692 454782
rect 481640 454718 481692 454724
rect 484412 454714 484440 500126
rect 485792 460222 485820 500126
rect 485780 460216 485832 460222
rect 485780 460158 485832 460164
rect 487172 457502 487200 500126
rect 488264 463004 488316 463010
rect 488264 462946 488316 462952
rect 487160 457496 487212 457502
rect 487160 457438 487212 457444
rect 484400 454708 484452 454714
rect 484400 454650 484452 454656
rect 487986 453928 488042 453937
rect 488276 453914 488304 462946
rect 488552 458862 488580 500126
rect 488540 458856 488592 458862
rect 488540 458798 488592 458804
rect 488042 453900 488304 453914
rect 488042 453886 488290 453900
rect 487986 453863 488042 453872
rect 471624 428466 471652 432140
rect 474292 430030 474320 432140
rect 474280 430024 474332 430030
rect 474280 429966 474332 429972
rect 476960 429962 476988 432140
rect 479352 432126 479642 432154
rect 481652 432126 482310 432154
rect 476948 429956 477000 429962
rect 476948 429898 477000 429904
rect 479352 429894 479380 432126
rect 479340 429888 479392 429894
rect 479340 429830 479392 429836
rect 479524 429888 479576 429894
rect 479524 429830 479576 429836
rect 471612 428460 471664 428466
rect 471612 428402 471664 428408
rect 471978 410544 472034 410553
rect 471978 410479 472034 410488
rect 470888 402946 471008 402974
rect 470980 385914 471008 402946
rect 471992 385914 472020 410479
rect 479536 389910 479564 429830
rect 481652 392630 481680 432126
rect 484964 429894 484992 432140
rect 484952 429888 485004 429894
rect 484952 429830 485004 429836
rect 487632 429214 487660 432140
rect 490024 432126 490314 432154
rect 486424 429208 486476 429214
rect 486424 429150 486476 429156
rect 487620 429208 487672 429214
rect 487620 429150 487672 429156
rect 483020 423428 483072 423434
rect 483020 423370 483072 423376
rect 481640 392624 481692 392630
rect 481640 392566 481692 392572
rect 479524 389904 479576 389910
rect 479524 389846 479576 389852
rect 483032 389298 483060 423370
rect 485780 423360 485832 423366
rect 485780 423302 485832 423308
rect 483112 421592 483164 421598
rect 483112 421534 483164 421540
rect 483020 389292 483072 389298
rect 483020 389234 483072 389240
rect 472898 389056 472954 389065
rect 472898 388991 472954 389000
rect 474370 389056 474426 389065
rect 474370 388991 474426 389000
rect 475106 389056 475162 389065
rect 475106 388991 475162 389000
rect 477314 389056 477370 389065
rect 477314 388991 477370 389000
rect 479522 389056 479578 389065
rect 479522 388991 479578 389000
rect 470980 385886 471454 385914
rect 471992 385886 472190 385914
rect 472912 385900 472940 388991
rect 473634 388920 473690 388929
rect 473634 388855 473690 388864
rect 473648 385900 473676 388855
rect 474384 385900 474412 388991
rect 475120 385900 475148 388991
rect 475842 388920 475898 388929
rect 475842 388855 475898 388864
rect 475856 385900 475884 388855
rect 476580 388612 476632 388618
rect 476580 388554 476632 388560
rect 476592 385900 476620 388554
rect 477328 385900 477356 388991
rect 478052 388952 478104 388958
rect 478052 388894 478104 388900
rect 478064 385900 478092 388894
rect 478788 388816 478840 388822
rect 478788 388758 478840 388764
rect 478800 385900 478828 388758
rect 479536 385900 479564 388991
rect 480260 388748 480312 388754
rect 480260 388690 480312 388696
rect 480272 385900 480300 388690
rect 482468 388680 482520 388686
rect 482468 388622 482520 388628
rect 481732 388544 481784 388550
rect 481732 388486 481784 388492
rect 480996 388476 481048 388482
rect 480996 388418 481048 388424
rect 481008 385900 481036 388418
rect 481744 385900 481772 388486
rect 482480 385900 482508 388622
rect 483124 385914 483152 421534
rect 483572 389292 483624 389298
rect 483572 389234 483624 389240
rect 483584 385914 483612 389234
rect 484676 388952 484728 388958
rect 484676 388894 484728 388900
rect 483124 385886 483230 385914
rect 483584 385886 483966 385914
rect 484688 385900 484716 388894
rect 485412 388680 485464 388686
rect 485412 388622 485464 388628
rect 485424 385900 485452 388622
rect 485792 385914 485820 423302
rect 486436 393990 486464 429150
rect 487160 423292 487212 423298
rect 487160 423234 487212 423240
rect 486424 393984 486476 393990
rect 486424 393926 486476 393932
rect 486884 388612 486936 388618
rect 486884 388554 486936 388560
rect 485792 385886 486174 385914
rect 486896 385900 486924 388554
rect 487172 385914 487200 423234
rect 488540 423224 488592 423230
rect 488540 423166 488592 423172
rect 488552 402974 488580 423166
rect 488552 402946 488672 402974
rect 488356 388476 488408 388482
rect 488356 388418 488408 388424
rect 487172 385886 487646 385914
rect 488368 385900 488396 388418
rect 488644 385914 488672 402946
rect 490024 395350 490052 432126
rect 490012 395344 490064 395350
rect 490012 395286 490064 395292
rect 490564 392624 490616 392630
rect 490564 392566 490616 392572
rect 489828 388544 489880 388550
rect 489828 388486 489880 388492
rect 488644 385886 489118 385914
rect 489840 385900 489868 388486
rect 490576 385900 490604 392566
rect 491128 391338 491156 500126
rect 491312 500126 491372 500154
rect 491116 391332 491168 391338
rect 491116 391274 491168 391280
rect 491312 387190 491340 500126
rect 494072 463010 494100 501191
rect 494060 463004 494112 463010
rect 494060 462946 494112 462952
rect 502984 423564 503036 423570
rect 502984 423506 503036 423512
rect 496820 423156 496872 423162
rect 496820 423098 496872 423104
rect 494060 420232 494112 420238
rect 494060 420174 494112 420180
rect 492680 398132 492732 398138
rect 492680 398074 492732 398080
rect 491576 395344 491628 395350
rect 491576 395286 491628 395292
rect 491392 393984 491444 393990
rect 491392 393926 491444 393932
rect 491300 387184 491352 387190
rect 491300 387126 491352 387132
rect 491404 387002 491432 393926
rect 491312 386974 491432 387002
rect 491312 385900 491340 386974
rect 491588 385914 491616 395286
rect 492692 389298 492720 398074
rect 492772 396772 492824 396778
rect 492772 396714 492824 396720
rect 492680 389292 492732 389298
rect 492680 389234 492732 389240
rect 491588 385886 492062 385914
rect 492784 385900 492812 396714
rect 494072 389298 494100 420174
rect 494152 399492 494204 399498
rect 494152 399434 494204 399440
rect 493140 389292 493192 389298
rect 493140 389234 493192 389240
rect 494060 389292 494112 389298
rect 494060 389234 494112 389240
rect 493152 385914 493180 389234
rect 494164 385914 494192 399434
rect 496452 391332 496504 391338
rect 496452 391274 496504 391280
rect 495716 389904 495768 389910
rect 495716 389846 495768 389852
rect 494612 389292 494664 389298
rect 494612 389234 494664 389240
rect 494624 385914 494652 389234
rect 493152 385886 493534 385914
rect 494164 385886 494270 385914
rect 494624 385886 495006 385914
rect 495728 385900 495756 389846
rect 496464 385900 496492 391274
rect 496832 385914 496860 423098
rect 498200 423088 498252 423094
rect 498200 423030 498252 423036
rect 497464 400920 497516 400926
rect 497464 400862 497516 400868
rect 497476 385914 497504 400862
rect 498212 385914 498240 423030
rect 499580 423020 499632 423026
rect 499580 422962 499632 422968
rect 499592 402974 499620 422962
rect 501052 422952 501104 422958
rect 501052 422894 501104 422900
rect 501064 402974 501092 422894
rect 499592 402946 499712 402974
rect 501064 402946 501184 402974
rect 499396 388884 499448 388890
rect 499396 388826 499448 388832
rect 496832 385886 497214 385914
rect 497476 385886 497950 385914
rect 498212 385886 498686 385914
rect 499408 385900 499436 388826
rect 499684 385914 499712 402946
rect 500868 388816 500920 388822
rect 500868 388758 500920 388764
rect 499684 385886 500158 385914
rect 500880 385900 500908 388758
rect 501156 385914 501184 402946
rect 502616 402280 502668 402286
rect 502616 402222 502668 402228
rect 502340 388748 502392 388754
rect 502340 388690 502392 388696
rect 501156 385886 501630 385914
rect 502352 385900 502380 388690
rect 502628 385914 502656 402222
rect 502996 388958 503024 423506
rect 509884 418192 509936 418198
rect 509884 418134 509936 418140
rect 503720 417784 503772 417790
rect 503720 417726 503772 417732
rect 502984 388952 503036 388958
rect 502984 388894 503036 388900
rect 503732 385914 503760 417726
rect 507860 417716 507912 417722
rect 507860 417658 507912 417664
rect 506480 417580 506532 417586
rect 506480 417522 506532 417528
rect 503996 417444 504048 417450
rect 503996 417386 504048 417392
rect 504008 402974 504036 417386
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 506020 391264 506072 391270
rect 506020 391206 506072 391212
rect 505284 389836 505336 389842
rect 505284 389778 505336 389784
rect 502628 385886 503102 385914
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 389778
rect 506032 385900 506060 391206
rect 506492 385914 506520 417522
rect 506572 417512 506624 417518
rect 506572 417454 506624 417460
rect 506584 402974 506612 417454
rect 506584 402946 507072 402974
rect 507044 385914 507072 402946
rect 507872 389298 507900 417658
rect 507952 417648 508004 417654
rect 507952 417590 508004 417596
rect 507860 389292 507912 389298
rect 507860 389234 507912 389240
rect 507964 385914 507992 417590
rect 508596 389292 508648 389298
rect 508596 389234 508648 389240
rect 508608 385914 508636 389234
rect 506492 385886 506782 385914
rect 507044 385886 507518 385914
rect 507964 385886 508254 385914
rect 508608 385886 508990 385914
rect 453304 385416 453356 385422
rect 453304 385358 453356 385364
rect 509606 372464 509662 372473
rect 509606 372399 509662 372408
rect 509330 367024 509386 367033
rect 509330 366959 509386 366968
rect 450726 322960 450782 322969
rect 450726 322895 450782 322904
rect 450636 321972 450688 321978
rect 450636 321914 450688 321920
rect 450544 321020 450596 321026
rect 450544 320962 450596 320968
rect 450358 319903 450414 319912
rect 450452 319932 450504 319938
rect 450452 319874 450504 319880
rect 450544 316736 450596 316742
rect 450544 316678 450596 316684
rect 449808 276752 449860 276758
rect 449808 276694 449860 276700
rect 449716 263560 449768 263566
rect 449716 263502 449768 263508
rect 447968 220108 448020 220114
rect 447968 220050 448020 220056
rect 447508 163532 447560 163538
rect 447508 163474 447560 163480
rect 447152 161446 447824 161474
rect 431328 159868 431678 159882
rect 431328 159854 431664 159868
rect 434976 159854 435312 159882
rect 438288 159854 438624 159882
rect 441586 160126 441660 160154
rect 445208 160200 445260 160206
rect 445208 160142 445260 160148
rect 445668 160200 445720 160206
rect 445668 160142 445720 160148
rect 441586 159868 441614 160126
rect 445220 159882 445248 160142
rect 444912 159854 445248 159882
rect 447796 159882 447824 161446
rect 447796 159854 448224 159882
rect 421432 159332 421728 159338
rect 421380 159326 421728 159332
rect 421392 159310 421728 159326
rect 410616 128308 410668 128314
rect 410616 128250 410668 128256
rect 439136 107296 439188 107302
rect 439136 107238 439188 107244
rect 432972 107228 433024 107234
rect 432972 107170 433024 107176
rect 426808 107160 426860 107166
rect 426808 107102 426860 107108
rect 420644 107092 420696 107098
rect 420644 107034 420696 107040
rect 414480 107024 414532 107030
rect 414480 106966 414532 106972
rect 410524 106276 410576 106282
rect 410524 106218 410576 106224
rect 414492 104938 414520 106966
rect 420656 104938 420684 107034
rect 426820 104938 426848 107102
rect 432984 104938 433012 107170
rect 439148 104938 439176 107238
rect 450556 106554 450584 316678
rect 450740 316034 450768 322895
rect 507306 322688 507362 322697
rect 507306 322623 507362 322632
rect 507122 322552 507178 322561
rect 507122 322487 507178 322496
rect 470152 322386 470258 322402
rect 470140 322380 470258 322386
rect 470192 322374 470258 322380
rect 470140 322322 470192 322328
rect 483112 322312 483164 322318
rect 479812 322250 479918 322266
rect 483164 322260 483230 322266
rect 483112 322254 483230 322260
rect 479800 322244 479918 322250
rect 479852 322238 479918 322244
rect 483124 322238 483230 322254
rect 479800 322186 479852 322192
rect 471796 322176 471848 322182
rect 454328 322102 454526 322130
rect 454696 322102 454802 322130
rect 454972 322102 455078 322130
rect 455248 322102 455354 322130
rect 454040 319184 454092 319190
rect 454040 319126 454092 319132
rect 453304 316872 453356 316878
rect 453304 316814 453356 316820
rect 450740 316006 450952 316034
rect 450728 315376 450780 315382
rect 450728 315318 450780 315324
rect 450636 315308 450688 315314
rect 450636 315250 450688 315256
rect 450648 107302 450676 315250
rect 450636 107296 450688 107302
rect 450636 107238 450688 107244
rect 450740 107098 450768 315318
rect 450820 313948 450872 313954
rect 450820 313890 450872 313896
rect 450832 107166 450860 313890
rect 450924 206310 450952 316006
rect 451924 311296 451976 311302
rect 451924 311238 451976 311244
rect 450912 206304 450964 206310
rect 450912 206246 450964 206252
rect 450912 160336 450964 160342
rect 450912 160278 450964 160284
rect 450924 142866 450952 160278
rect 451556 158432 451608 158438
rect 451556 158374 451608 158380
rect 451568 158273 451596 158374
rect 451554 158264 451610 158273
rect 451554 158199 451610 158208
rect 451740 157344 451792 157350
rect 451740 157286 451792 157292
rect 451752 156913 451780 157286
rect 451738 156904 451794 156913
rect 451738 156839 451794 156848
rect 451740 154556 451792 154562
rect 451740 154498 451792 154504
rect 451752 154193 451780 154498
rect 451738 154184 451794 154193
rect 451738 154119 451794 154128
rect 451648 153196 451700 153202
rect 451648 153138 451700 153144
rect 451660 152833 451688 153138
rect 451646 152824 451702 152833
rect 451646 152759 451702 152768
rect 451464 151496 451516 151502
rect 451462 151464 451464 151473
rect 451516 151464 451518 151473
rect 451462 151399 451518 151408
rect 450912 142860 450964 142866
rect 450912 142802 450964 142808
rect 451556 139392 451608 139398
rect 451556 139334 451608 139340
rect 451568 139233 451596 139334
rect 451554 139224 451610 139233
rect 451554 139159 451610 139168
rect 451936 124273 451964 311238
rect 452016 309868 452068 309874
rect 452016 309810 452068 309816
rect 452028 128353 452056 309810
rect 452200 305448 452252 305454
rect 452200 305390 452252 305396
rect 452108 283688 452160 283694
rect 452108 283630 452160 283636
rect 452014 128344 452070 128353
rect 452014 128279 452070 128288
rect 452120 125633 452148 283630
rect 452212 148753 452240 305390
rect 452384 280900 452436 280906
rect 452384 280842 452436 280848
rect 452292 271176 452344 271182
rect 452292 271118 452344 271124
rect 452198 148744 452254 148753
rect 452198 148679 452254 148688
rect 452200 132456 452252 132462
rect 452198 132424 452200 132433
rect 452252 132424 452254 132433
rect 452198 132359 452254 132368
rect 452304 129713 452332 271118
rect 452396 150113 452424 280842
rect 452568 155576 452620 155582
rect 452566 155544 452568 155553
rect 452620 155544 452622 155553
rect 452566 155479 452622 155488
rect 452382 150104 452438 150113
rect 452382 150039 452438 150048
rect 452568 147552 452620 147558
rect 452568 147494 452620 147500
rect 452580 147393 452608 147494
rect 452566 147384 452622 147393
rect 452566 147319 452622 147328
rect 452568 146056 452620 146062
rect 452566 146024 452568 146033
rect 452620 146024 452622 146033
rect 452566 145959 452622 145968
rect 452568 144696 452620 144702
rect 452566 144664 452568 144673
rect 452620 144664 452622 144673
rect 452566 144599 452622 144608
rect 452568 143336 452620 143342
rect 452566 143304 452568 143313
rect 452620 143304 452622 143313
rect 452566 143239 452622 143248
rect 452568 141976 452620 141982
rect 452566 141944 452568 141953
rect 452620 141944 452622 141953
rect 452566 141879 452622 141888
rect 452568 140684 452620 140690
rect 452568 140626 452620 140632
rect 452580 140593 452608 140626
rect 452566 140584 452622 140593
rect 452566 140519 452622 140528
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452568 136536 452620 136542
rect 452566 136504 452568 136513
rect 452620 136504 452622 136513
rect 452566 136439 452622 136448
rect 452568 135176 452620 135182
rect 452566 135144 452568 135153
rect 452620 135144 452622 135153
rect 452566 135079 452622 135088
rect 452568 133816 452620 133822
rect 452566 133784 452568 133793
rect 452620 133784 452622 133793
rect 452566 133719 452622 133728
rect 453316 132462 453344 316814
rect 453396 308440 453448 308446
rect 453396 308382 453448 308388
rect 453304 132456 453356 132462
rect 453304 132398 453356 132404
rect 453408 131102 453436 308382
rect 454052 287706 454080 319126
rect 454224 319116 454276 319122
rect 454224 319058 454276 319064
rect 454132 319048 454184 319054
rect 454132 318990 454184 318996
rect 454144 294506 454172 318990
rect 454236 296002 454264 319058
rect 454328 297974 454356 322102
rect 454696 319122 454724 322102
rect 454684 319116 454736 319122
rect 454684 319058 454736 319064
rect 454972 319054 455000 322102
rect 455248 319190 455276 322102
rect 455236 319184 455288 319190
rect 455236 319126 455288 319132
rect 455512 319116 455564 319122
rect 455512 319058 455564 319064
rect 454960 319048 455012 319054
rect 454960 318990 455012 318996
rect 454684 316804 454736 316810
rect 454684 316746 454736 316752
rect 454316 297968 454368 297974
rect 454316 297910 454368 297916
rect 454224 295996 454276 296002
rect 454224 295938 454276 295944
rect 454132 294500 454184 294506
rect 454132 294442 454184 294448
rect 454132 288992 454184 288998
rect 454132 288934 454184 288940
rect 454040 287700 454092 287706
rect 454040 287642 454092 287648
rect 453488 285048 453540 285054
rect 453488 284990 453540 284996
rect 452384 131096 452436 131102
rect 452382 131064 452384 131073
rect 453396 131096 453448 131102
rect 452436 131064 452438 131073
rect 453396 131038 453448 131044
rect 452382 130999 452438 131008
rect 452290 129704 452346 129713
rect 452290 129639 452346 129648
rect 452382 126984 452438 126993
rect 453500 126954 453528 284990
rect 454144 283626 454172 288934
rect 454132 283620 454184 283626
rect 454132 283562 454184 283568
rect 453580 278044 453632 278050
rect 453580 277986 453632 277992
rect 453592 153202 453620 277986
rect 453672 272536 453724 272542
rect 453672 272478 453724 272484
rect 453580 153196 453632 153202
rect 453580 153138 453632 153144
rect 453684 151502 453712 272478
rect 453856 227792 453908 227798
rect 453856 227734 453908 227740
rect 453868 221474 453896 227734
rect 453856 221468 453908 221474
rect 453856 221410 453908 221416
rect 453672 151496 453724 151502
rect 453672 151438 453724 151444
rect 452382 126919 452384 126928
rect 452436 126919 452438 126928
rect 453488 126948 453540 126954
rect 452384 126890 452436 126896
rect 453488 126890 453540 126896
rect 452106 125624 452162 125633
rect 452106 125559 452162 125568
rect 451922 124264 451978 124273
rect 451922 124199 451978 124208
rect 451924 123412 451976 123418
rect 451924 123354 451976 123360
rect 451936 122913 451964 123354
rect 451922 122904 451978 122913
rect 451922 122839 451978 122848
rect 451924 122188 451976 122194
rect 451924 122130 451976 122136
rect 451936 121553 451964 122130
rect 451922 121544 451978 121553
rect 451922 121479 451978 121488
rect 451188 107432 451240 107438
rect 451188 107374 451240 107380
rect 450820 107160 450872 107166
rect 450820 107102 450872 107108
rect 450728 107092 450780 107098
rect 450728 107034 450780 107040
rect 445300 106548 445352 106554
rect 445300 106490 445352 106496
rect 450544 106548 450596 106554
rect 450544 106490 450596 106496
rect 445312 104938 445340 106490
rect 451200 104938 451228 107374
rect 454696 106962 454724 316746
rect 454776 298036 454828 298042
rect 454776 297978 454828 297984
rect 454788 107030 454816 297978
rect 455524 290494 455552 319058
rect 455616 311166 455644 322116
rect 455800 322102 455906 322130
rect 456076 322102 456182 322130
rect 455604 311160 455656 311166
rect 455604 311102 455656 311108
rect 455800 305794 455828 322102
rect 456076 319122 456104 322102
rect 456064 319116 456116 319122
rect 456064 319058 456116 319064
rect 456444 318170 456472 322116
rect 456720 321570 456748 322116
rect 456708 321564 456760 321570
rect 456708 321506 456760 321512
rect 456996 321502 457024 322116
rect 456984 321496 457036 321502
rect 456984 321438 457036 321444
rect 456800 320884 456852 320890
rect 456800 320826 456852 320832
rect 456812 320074 456840 320826
rect 457272 320142 457300 322116
rect 457548 321774 457576 322116
rect 457536 321768 457588 321774
rect 457536 321710 457588 321716
rect 457824 321638 457852 322116
rect 458100 321706 458128 322116
rect 458088 321700 458140 321706
rect 458088 321642 458140 321648
rect 457812 321632 457864 321638
rect 457812 321574 457864 321580
rect 458376 321434 458404 322116
rect 458652 321473 458680 322116
rect 458638 321464 458694 321473
rect 458364 321428 458416 321434
rect 458638 321399 458694 321408
rect 458364 321370 458416 321376
rect 457260 320136 457312 320142
rect 457260 320078 457312 320084
rect 456800 320068 456852 320074
rect 456800 320010 456852 320016
rect 458928 319870 458956 322116
rect 459204 321230 459232 322116
rect 459480 321298 459508 322116
rect 459468 321292 459520 321298
rect 459468 321234 459520 321240
rect 459192 321224 459244 321230
rect 459756 321201 459784 322116
rect 459192 321166 459244 321172
rect 459742 321192 459798 321201
rect 459742 321127 459798 321136
rect 460032 320958 460060 322116
rect 460308 321881 460336 322116
rect 460294 321872 460350 321881
rect 460294 321807 460350 321816
rect 460584 321065 460612 322116
rect 460768 322102 460874 322130
rect 460768 321978 460796 322102
rect 460756 321972 460808 321978
rect 460756 321914 460808 321920
rect 461136 321094 461164 322116
rect 461412 321366 461440 322116
rect 461400 321360 461452 321366
rect 461400 321302 461452 321308
rect 461124 321088 461176 321094
rect 460570 321056 460626 321065
rect 461124 321030 461176 321036
rect 460570 320991 460626 321000
rect 460020 320952 460072 320958
rect 460020 320894 460072 320900
rect 460204 320952 460256 320958
rect 460204 320894 460256 320900
rect 459560 320884 459612 320890
rect 459560 320826 459612 320832
rect 459572 320142 459600 320826
rect 459560 320136 459612 320142
rect 459560 320078 459612 320084
rect 458916 319864 458968 319870
rect 458916 319806 458968 319812
rect 456432 318164 456484 318170
rect 456432 318106 456484 318112
rect 458824 318164 458876 318170
rect 458824 318106 458876 318112
rect 456892 318096 456944 318102
rect 456892 318038 456944 318044
rect 456064 311228 456116 311234
rect 456064 311170 456116 311176
rect 455788 305788 455840 305794
rect 455788 305730 455840 305736
rect 455512 290488 455564 290494
rect 455512 290430 455564 290436
rect 454960 279472 455012 279478
rect 454960 279414 455012 279420
rect 454868 268388 454920 268394
rect 454868 268330 454920 268336
rect 454880 107438 454908 268330
rect 454972 123418 455000 279414
rect 455052 274032 455104 274038
rect 455052 273974 455104 273980
rect 455064 143342 455092 273974
rect 455144 269952 455196 269958
rect 455144 269894 455196 269900
rect 455156 158438 455184 269894
rect 455144 158432 455196 158438
rect 455144 158374 455196 158380
rect 455052 143336 455104 143342
rect 455052 143278 455104 143284
rect 454960 123412 455012 123418
rect 454960 123354 455012 123360
rect 454868 107432 454920 107438
rect 454868 107374 454920 107380
rect 456076 107234 456104 311170
rect 456340 276820 456392 276826
rect 456340 276762 456392 276768
rect 456248 271312 456300 271318
rect 456248 271254 456300 271260
rect 456156 271244 456208 271250
rect 456156 271186 456208 271192
rect 456168 136542 456196 271186
rect 456260 140690 456288 271254
rect 456352 147558 456380 276762
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 456904 258074 456932 318038
rect 457812 317076 457864 317082
rect 457812 317018 457864 317024
rect 457444 316940 457496 316946
rect 457444 316882 457496 316888
rect 457076 268456 457128 268462
rect 457076 268398 457128 268404
rect 457088 258074 457116 268398
rect 456812 258046 456932 258074
rect 456996 258046 457116 258074
rect 456812 249082 456840 258046
rect 456800 249076 456852 249082
rect 456800 249018 456852 249024
rect 456812 248849 456840 249018
rect 456798 248840 456854 248849
rect 456798 248775 456854 248784
rect 456798 207224 456854 207233
rect 456798 207159 456854 207168
rect 456812 206310 456840 207159
rect 456800 206304 456852 206310
rect 456800 206246 456852 206252
rect 456812 200802 456840 206246
rect 456800 200796 456852 200802
rect 456800 200738 456852 200744
rect 456340 147552 456392 147558
rect 456340 147494 456392 147500
rect 456248 140684 456300 140690
rect 456248 140626 456300 140632
rect 456156 136536 456208 136542
rect 456156 136478 456208 136484
rect 456064 107228 456116 107234
rect 456064 107170 456116 107176
rect 454776 107024 454828 107030
rect 454776 106966 454828 106972
rect 454684 106956 454736 106962
rect 454684 106898 454736 106904
rect 407592 104910 408020 104938
rect 414184 104910 414520 104938
rect 420348 104910 420684 104938
rect 426512 104910 426848 104938
rect 432676 104910 433012 104938
rect 438840 104910 439176 104938
rect 445004 104910 445340 104938
rect 451168 104910 451228 104938
rect 456996 104938 457024 258046
rect 457456 139398 457484 316882
rect 457536 291712 457588 291718
rect 457536 291654 457588 291660
rect 457444 139392 457496 139398
rect 457444 139334 457496 139340
rect 457548 135182 457576 291654
rect 457628 275460 457680 275466
rect 457628 275402 457680 275408
rect 457536 135176 457588 135182
rect 457536 135118 457588 135124
rect 457640 133822 457668 275402
rect 457720 275392 457772 275398
rect 457720 275334 457772 275340
rect 457732 144702 457760 275334
rect 457824 234977 457852 317018
rect 457810 234968 457866 234977
rect 457810 234903 457866 234912
rect 458086 234968 458142 234977
rect 458086 234903 458142 234912
rect 458100 162178 458128 234903
rect 458088 162172 458140 162178
rect 458088 162114 458140 162120
rect 457720 144696 457772 144702
rect 457720 144638 457772 144644
rect 457628 133816 457680 133822
rect 457628 133758 457680 133764
rect 458836 122194 458864 318106
rect 459100 318028 459152 318034
rect 459100 317970 459152 317976
rect 458916 315444 458968 315450
rect 458916 315386 458968 315392
rect 458928 141982 458956 315386
rect 459008 314016 459060 314022
rect 459008 313958 459060 313964
rect 459020 146062 459048 313958
rect 459112 154562 459140 317970
rect 459284 282260 459336 282266
rect 459284 282202 459336 282208
rect 459192 272604 459244 272610
rect 459192 272546 459244 272552
rect 459100 154556 459152 154562
rect 459100 154498 459152 154504
rect 459008 146056 459060 146062
rect 459008 145998 459060 146004
rect 458916 141976 458968 141982
rect 458916 141918 458968 141924
rect 459204 137902 459232 272546
rect 459296 155582 459324 282202
rect 459376 268592 459428 268598
rect 459376 268534 459428 268540
rect 459388 227798 459416 268534
rect 459376 227792 459428 227798
rect 459376 227734 459428 227740
rect 459466 221096 459522 221105
rect 459466 221031 459522 221040
rect 459480 220114 459508 221031
rect 459468 220108 459520 220114
rect 459468 220050 459520 220056
rect 459480 199442 459508 220050
rect 459468 199436 459520 199442
rect 459468 199378 459520 199384
rect 459284 155576 459336 155582
rect 459284 155518 459336 155524
rect 459192 137896 459244 137902
rect 459192 137838 459244 137844
rect 458824 122188 458876 122194
rect 458824 122130 458876 122136
rect 456996 104910 457332 104938
rect 386328 33924 386380 33930
rect 386328 33866 386380 33872
rect 386236 31408 386288 31414
rect 386236 31350 386288 31356
rect 460216 29646 460244 320894
rect 461688 319938 461716 322116
rect 461964 321910 461992 322116
rect 461952 321904 462004 321910
rect 461952 321846 462004 321852
rect 462240 320006 462268 322116
rect 462516 321842 462544 322116
rect 462504 321836 462556 321842
rect 462504 321778 462556 321784
rect 462228 320000 462280 320006
rect 462228 319942 462280 319948
rect 461676 319932 461728 319938
rect 461676 319874 461728 319880
rect 462688 319116 462740 319122
rect 462688 319058 462740 319064
rect 462412 319048 462464 319054
rect 462412 318990 462464 318996
rect 461584 318096 461636 318102
rect 461584 318038 461636 318044
rect 461596 299470 461624 318038
rect 462424 302802 462452 318990
rect 462412 302796 462464 302802
rect 462412 302738 462464 302744
rect 462700 302734 462728 319058
rect 462792 317014 462820 322116
rect 462976 322102 463082 322130
rect 463252 322102 463358 322130
rect 463528 322102 463634 322130
rect 463910 322102 464108 322130
rect 462780 317008 462832 317014
rect 462780 316950 462832 316956
rect 462976 308514 463004 322102
rect 463252 319054 463280 322102
rect 463528 319122 463556 322102
rect 463516 319116 463568 319122
rect 463516 319058 463568 319064
rect 463792 319116 463844 319122
rect 463792 319058 463844 319064
rect 463240 319048 463292 319054
rect 463240 318990 463292 318996
rect 462964 308508 463016 308514
rect 462964 308450 463016 308456
rect 463804 303618 463832 319058
rect 464080 306338 464108 322102
rect 464068 306332 464120 306338
rect 464068 306274 464120 306280
rect 464172 305522 464200 322116
rect 464356 322102 464462 322130
rect 464632 322102 464738 322130
rect 464908 322102 465014 322130
rect 464356 319274 464384 322102
rect 464264 319246 464384 319274
rect 464264 316062 464292 319246
rect 464632 319002 464660 322102
rect 464908 319122 464936 322102
rect 464896 319116 464948 319122
rect 464896 319058 464948 319064
rect 464356 318974 464660 319002
rect 465172 319048 465224 319054
rect 465172 318990 465224 318996
rect 464252 316056 464304 316062
rect 464252 315998 464304 316004
rect 464160 305516 464212 305522
rect 464160 305458 464212 305464
rect 463792 303612 463844 303618
rect 463792 303554 463844 303560
rect 462688 302728 462740 302734
rect 462688 302670 462740 302676
rect 464356 302666 464384 318974
rect 464436 316056 464488 316062
rect 464436 315998 464488 316004
rect 464448 305590 464476 315998
rect 464436 305584 464488 305590
rect 464436 305526 464488 305532
rect 464344 302660 464396 302666
rect 464344 302602 464396 302608
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 465184 280838 465212 318990
rect 465276 312594 465304 322116
rect 465448 319116 465500 319122
rect 465448 319058 465500 319064
rect 465264 312588 465316 312594
rect 465264 312530 465316 312536
rect 465356 291236 465408 291242
rect 465356 291178 465408 291184
rect 465368 288998 465396 291178
rect 465356 288992 465408 288998
rect 465356 288934 465408 288940
rect 465460 282198 465488 319058
rect 465552 300014 465580 322116
rect 465736 322102 465842 322130
rect 466012 322102 466118 322130
rect 466288 322102 466394 322130
rect 466564 322102 466670 322130
rect 466840 322102 466946 322130
rect 465540 300008 465592 300014
rect 465540 299950 465592 299956
rect 465736 283626 465764 322102
rect 466012 319122 466040 322102
rect 466000 319116 466052 319122
rect 466000 319058 466052 319064
rect 466288 319054 466316 322102
rect 466276 319048 466328 319054
rect 466276 318990 466328 318996
rect 465724 283620 465776 283626
rect 465724 283562 465776 283568
rect 465448 282192 465500 282198
rect 465448 282134 465500 282140
rect 465172 280832 465224 280838
rect 465172 280774 465224 280780
rect 465724 275528 465776 275534
rect 465724 275470 465776 275476
rect 460296 274100 460348 274106
rect 460296 274042 460348 274048
rect 460308 157350 460336 274042
rect 465736 268598 465764 275470
rect 466564 269890 466592 322102
rect 466840 313274 466868 322102
rect 467208 321298 467236 322116
rect 467498 322102 467696 322130
rect 467668 321978 467696 322102
rect 467656 321972 467708 321978
rect 467656 321914 467708 321920
rect 467760 321842 467788 322116
rect 467748 321836 467800 321842
rect 467748 321778 467800 321784
rect 467196 321292 467248 321298
rect 467196 321234 467248 321240
rect 468036 321094 468064 322116
rect 468312 321910 468340 322116
rect 468300 321904 468352 321910
rect 468300 321846 468352 321852
rect 468588 321366 468616 322116
rect 468576 321360 468628 321366
rect 468576 321302 468628 321308
rect 468024 321088 468076 321094
rect 468024 321030 468076 321036
rect 468864 319870 468892 322116
rect 469140 320006 469168 322116
rect 469128 320000 469180 320006
rect 469128 319942 469180 319948
rect 468852 319864 468904 319870
rect 468852 319806 468904 319812
rect 469416 318782 469444 322116
rect 469692 319258 469720 322116
rect 469968 319734 469996 322116
rect 469956 319728 470008 319734
rect 469956 319670 470008 319676
rect 470520 319462 470548 322116
rect 470704 322102 470810 322130
rect 477868 322176 477920 322182
rect 471848 322124 471914 322130
rect 471796 322118 471914 322124
rect 470704 322046 470732 322102
rect 470692 322040 470744 322046
rect 470692 321982 470744 321988
rect 471072 320113 471100 322116
rect 471058 320104 471114 320113
rect 471058 320039 471114 320048
rect 471348 319841 471376 322116
rect 471624 319977 471652 322116
rect 471808 322102 471914 322118
rect 471610 319968 471666 319977
rect 471610 319903 471666 319912
rect 471334 319832 471390 319841
rect 471334 319767 471390 319776
rect 470508 319456 470560 319462
rect 470508 319398 470560 319404
rect 472176 319326 472204 322116
rect 472452 319802 472480 322116
rect 472440 319796 472492 319802
rect 472440 319738 472492 319744
rect 472728 319666 472756 322116
rect 473004 320074 473032 322116
rect 473188 322102 473294 322130
rect 472992 320068 473044 320074
rect 472992 320010 473044 320016
rect 472716 319660 472768 319666
rect 472716 319602 472768 319608
rect 472164 319320 472216 319326
rect 472164 319262 472216 319268
rect 469680 319252 469732 319258
rect 469680 319194 469732 319200
rect 469404 318776 469456 318782
rect 469404 318718 469456 318724
rect 473188 316034 473216 322102
rect 473452 319252 473504 319258
rect 473452 319194 473504 319200
rect 472360 316006 473216 316034
rect 472360 314702 472388 316006
rect 469864 314696 469916 314702
rect 469864 314638 469916 314644
rect 472348 314696 472400 314702
rect 472348 314638 472400 314644
rect 466828 313268 466880 313274
rect 466828 313210 466880 313216
rect 469876 291242 469904 314638
rect 473464 302870 473492 319194
rect 473452 302864 473504 302870
rect 473452 302806 473504 302812
rect 473556 299946 473584 322116
rect 473740 322102 473846 322130
rect 474016 322102 474122 322130
rect 474292 322102 474398 322130
rect 474568 322102 474674 322130
rect 473740 319258 473768 322102
rect 473728 319252 473780 319258
rect 473728 319194 473780 319200
rect 474016 319138 474044 322102
rect 473740 319110 474044 319138
rect 473740 306066 473768 319110
rect 474292 319002 474320 322102
rect 474016 318974 474320 319002
rect 474016 306202 474044 318974
rect 474568 316034 474596 322102
rect 474832 319048 474884 319054
rect 474832 318990 474884 318996
rect 474292 316006 474596 316034
rect 474292 306270 474320 316006
rect 474280 306264 474332 306270
rect 474280 306206 474332 306212
rect 474004 306196 474056 306202
rect 474004 306138 474056 306144
rect 473728 306060 473780 306066
rect 473728 306002 473780 306008
rect 473544 299940 473596 299946
rect 473544 299882 473596 299888
rect 469864 291236 469916 291242
rect 469864 291178 469916 291184
rect 474844 288998 474872 318990
rect 474936 306134 474964 322116
rect 475108 319116 475160 319122
rect 475108 319058 475160 319064
rect 475120 307086 475148 319058
rect 475108 307080 475160 307086
rect 475108 307022 475160 307028
rect 474924 306128 474976 306134
rect 474924 306070 474976 306076
rect 474832 288992 474884 288998
rect 474832 288934 474884 288940
rect 475212 275330 475240 322116
rect 475396 322102 475502 322130
rect 475672 322102 475778 322130
rect 475948 322102 476054 322130
rect 475396 309806 475424 322102
rect 475672 319054 475700 322102
rect 475948 319122 475976 322102
rect 475936 319116 475988 319122
rect 475936 319058 475988 319064
rect 476212 319116 476264 319122
rect 476212 319058 476264 319064
rect 475660 319048 475712 319054
rect 475660 318990 475712 318996
rect 475384 309800 475436 309806
rect 475384 309742 475436 309748
rect 475384 285728 475436 285734
rect 475384 285670 475436 285676
rect 475200 275324 475252 275330
rect 475200 275266 475252 275272
rect 466552 269884 466604 269890
rect 466552 269826 466604 269832
rect 465724 268592 465776 268598
rect 465724 268534 465776 268540
rect 475396 268530 475424 285670
rect 476224 284986 476252 319058
rect 476316 301646 476344 322116
rect 476500 322102 476606 322130
rect 476776 322102 476882 322130
rect 477710 322124 477868 322130
rect 477710 322118 477920 322124
rect 476304 301640 476356 301646
rect 476304 301582 476356 301588
rect 476500 293282 476528 322102
rect 476776 319122 476804 322102
rect 476764 319116 476816 319122
rect 476764 319058 476816 319064
rect 477144 318374 477172 322116
rect 477420 319802 477448 322116
rect 477710 322102 477908 322118
rect 477972 321230 478000 322116
rect 478262 322102 478460 322130
rect 478432 322046 478460 322102
rect 478420 322040 478472 322046
rect 478420 321982 478472 321988
rect 477960 321224 478012 321230
rect 477960 321166 478012 321172
rect 478524 319938 478552 322116
rect 478800 320074 478828 322116
rect 479076 320142 479104 322116
rect 479352 321162 479380 322116
rect 479340 321156 479392 321162
rect 479340 321098 479392 321104
rect 479064 320136 479116 320142
rect 479628 320113 479656 322116
rect 480180 320822 480208 322116
rect 480456 321337 480484 322116
rect 480442 321328 480498 321337
rect 480442 321263 480498 321272
rect 480168 320816 480220 320822
rect 480168 320758 480220 320764
rect 480732 320686 480760 322116
rect 480720 320680 480772 320686
rect 480720 320622 480772 320628
rect 479064 320078 479116 320084
rect 479614 320104 479670 320113
rect 478788 320068 478840 320074
rect 479614 320039 479670 320048
rect 478788 320010 478840 320016
rect 478512 319932 478564 319938
rect 478512 319874 478564 319880
rect 477408 319796 477460 319802
rect 477408 319738 477460 319744
rect 481008 319598 481036 322116
rect 481284 321026 481312 322116
rect 481560 321745 481588 322116
rect 481546 321736 481602 321745
rect 481546 321671 481602 321680
rect 481836 321609 481864 322116
rect 481822 321600 481878 321609
rect 481822 321535 481878 321544
rect 481272 321020 481324 321026
rect 481272 320962 481324 320968
rect 482112 320754 482140 322116
rect 482100 320748 482152 320754
rect 482100 320690 482152 320696
rect 480996 319592 481048 319598
rect 480996 319534 481048 319540
rect 482388 319394 482416 322116
rect 482572 322114 482678 322130
rect 482560 322108 482678 322114
rect 482612 322102 482678 322108
rect 482560 322050 482612 322056
rect 482940 319530 482968 322116
rect 483400 322102 483506 322130
rect 482928 319524 482980 319530
rect 482928 319466 482980 319472
rect 482376 319388 482428 319394
rect 482376 319330 482428 319336
rect 483112 319116 483164 319122
rect 483112 319058 483164 319064
rect 480904 319048 480956 319054
rect 480904 318990 480956 318996
rect 477132 318368 477184 318374
rect 477132 318310 477184 318316
rect 479524 318368 479576 318374
rect 479524 318310 479576 318316
rect 478144 307828 478196 307834
rect 478144 307770 478196 307776
rect 476488 293276 476540 293282
rect 476488 293218 476540 293224
rect 478156 285734 478184 307770
rect 478236 291644 478288 291650
rect 478236 291586 478288 291592
rect 478144 285728 478196 285734
rect 478144 285670 478196 285676
rect 476212 284980 476264 284986
rect 476212 284922 476264 284928
rect 478248 275534 478276 291586
rect 478236 275528 478288 275534
rect 478236 275470 478288 275476
rect 479536 273222 479564 318310
rect 480916 307834 480944 318990
rect 480904 307828 480956 307834
rect 480904 307770 480956 307776
rect 483124 300082 483152 319058
rect 483112 300076 483164 300082
rect 483112 300018 483164 300024
rect 483400 291650 483428 322102
rect 483768 319054 483796 322116
rect 483952 322102 484058 322130
rect 484228 322102 484334 322130
rect 483952 319122 483980 322102
rect 483940 319116 483992 319122
rect 483940 319058 483992 319064
rect 483756 319048 483808 319054
rect 483756 318990 483808 318996
rect 484228 316034 484256 322102
rect 484492 319116 484544 319122
rect 484492 319058 484544 319064
rect 483676 316006 484256 316034
rect 483676 303550 483704 316006
rect 484504 306241 484532 319058
rect 484490 306232 484546 306241
rect 484490 306167 484546 306176
rect 484596 305862 484624 322116
rect 484780 322102 484886 322130
rect 484780 305998 484808 322102
rect 485044 318844 485096 318850
rect 485044 318786 485096 318792
rect 484768 305992 484820 305998
rect 484768 305934 484820 305940
rect 484584 305856 484636 305862
rect 484584 305798 484636 305804
rect 483664 303544 483716 303550
rect 483664 303486 483716 303492
rect 483388 291644 483440 291650
rect 483388 291586 483440 291592
rect 485056 273970 485084 318786
rect 485148 305930 485176 322116
rect 485332 322102 485438 322130
rect 485608 322102 485714 322130
rect 485332 318850 485360 322102
rect 485608 319122 485636 322102
rect 485596 319116 485648 319122
rect 485596 319058 485648 319064
rect 485320 318844 485372 318850
rect 485320 318786 485372 318792
rect 485872 316600 485924 316606
rect 485872 316542 485924 316548
rect 485136 305924 485188 305930
rect 485136 305866 485188 305872
rect 485884 286890 485912 316542
rect 485976 307154 486004 322116
rect 486148 316668 486200 316674
rect 486148 316610 486200 316616
rect 485964 307148 486016 307154
rect 485964 307090 486016 307096
rect 486160 303550 486188 316610
rect 486252 304502 486280 322116
rect 486436 322102 486542 322130
rect 486712 322102 486818 322130
rect 486988 322102 487094 322130
rect 486436 316606 486464 322102
rect 486712 316674 486740 322102
rect 486700 316668 486752 316674
rect 486700 316610 486752 316616
rect 486424 316600 486476 316606
rect 486424 316542 486476 316548
rect 486988 311894 487016 322102
rect 487356 318170 487384 322116
rect 487540 322102 487646 322130
rect 487344 318164 487396 318170
rect 487344 318106 487396 318112
rect 487252 312180 487304 312186
rect 487252 312122 487304 312128
rect 486436 311866 487016 311894
rect 486240 304496 486292 304502
rect 486240 304438 486292 304444
rect 486148 303544 486200 303550
rect 486148 303486 486200 303492
rect 485872 286884 485924 286890
rect 485872 286826 485924 286832
rect 485044 273964 485096 273970
rect 485044 273906 485096 273912
rect 479524 273216 479576 273222
rect 479524 273158 479576 273164
rect 486436 269958 486464 311866
rect 487264 283694 487292 312122
rect 487252 283688 487304 283694
rect 487252 283630 487304 283636
rect 487540 279478 487568 322102
rect 487804 316668 487856 316674
rect 487804 316610 487856 316616
rect 487816 285054 487844 316610
rect 487908 311302 487936 322116
rect 488092 322102 488198 322130
rect 488368 322102 488474 322130
rect 488092 312186 488120 322102
rect 488368 316674 488396 322102
rect 488736 321554 488764 322116
rect 488920 322102 489026 322130
rect 489196 322102 489302 322130
rect 488736 321526 488856 321554
rect 488356 316668 488408 316674
rect 488356 316610 488408 316616
rect 488632 316668 488684 316674
rect 488632 316610 488684 316616
rect 488080 312180 488132 312186
rect 488080 312122 488132 312128
rect 487896 311296 487948 311302
rect 487896 311238 487948 311244
rect 487804 285048 487856 285054
rect 487804 284990 487856 284996
rect 487528 279472 487580 279478
rect 487528 279414 487580 279420
rect 488644 275466 488672 316610
rect 488828 309874 488856 321526
rect 488816 309868 488868 309874
rect 488816 309810 488868 309816
rect 488632 275460 488684 275466
rect 488632 275402 488684 275408
rect 488920 271182 488948 322102
rect 489196 308446 489224 322102
rect 489564 316878 489592 322116
rect 489748 322102 489854 322130
rect 489552 316872 489604 316878
rect 489552 316814 489604 316820
rect 489748 316674 489776 322102
rect 490012 316872 490064 316878
rect 490012 316814 490064 316820
rect 489736 316668 489788 316674
rect 489736 316610 489788 316616
rect 489184 308440 489236 308446
rect 489184 308382 489236 308388
rect 490024 271250 490052 316814
rect 490116 311894 490144 322116
rect 490300 322102 490406 322130
rect 490576 322102 490682 322130
rect 490300 316878 490328 322102
rect 490288 316872 490340 316878
rect 490288 316814 490340 316820
rect 490288 316600 490340 316606
rect 490288 316542 490340 316548
rect 490116 311866 490236 311894
rect 490208 291718 490236 311866
rect 490196 291712 490248 291718
rect 490196 291654 490248 291660
rect 490300 271318 490328 316542
rect 490576 272610 490604 322102
rect 490944 316946 490972 322116
rect 491128 322102 491234 322130
rect 491404 322102 491510 322130
rect 491680 322102 491786 322130
rect 491956 322102 492062 322130
rect 490932 316940 490984 316946
rect 490932 316882 490984 316888
rect 491128 316606 491156 322102
rect 491116 316600 491168 316606
rect 491116 316542 491168 316548
rect 491404 315450 491432 322102
rect 491392 315444 491444 315450
rect 491392 315386 491444 315392
rect 491680 274038 491708 322102
rect 491956 275398 491984 322102
rect 492324 314022 492352 322116
rect 492508 322102 492614 322130
rect 492312 314016 492364 314022
rect 492312 313958 492364 313964
rect 492508 311894 492536 322102
rect 492876 321554 492904 322116
rect 492876 321526 492996 321554
rect 492772 316668 492824 316674
rect 492772 316610 492824 316616
rect 492232 311866 492536 311894
rect 492232 276826 492260 311866
rect 492784 278050 492812 316610
rect 492968 305454 492996 321526
rect 493152 316878 493180 322116
rect 493336 322102 493442 322130
rect 493612 322102 493718 322130
rect 493336 321554 493364 322102
rect 493244 321526 493364 321554
rect 493140 316872 493192 316878
rect 493140 316814 493192 316820
rect 493244 313970 493272 321526
rect 493324 316872 493376 316878
rect 493324 316814 493376 316820
rect 493060 313942 493272 313970
rect 492956 305448 493008 305454
rect 492956 305390 493008 305396
rect 492772 278044 492824 278050
rect 492772 277986 492824 277992
rect 492220 276820 492272 276826
rect 492220 276762 492272 276768
rect 491944 275392 491996 275398
rect 491944 275334 491996 275340
rect 491668 274032 491720 274038
rect 491668 273974 491720 273980
rect 490564 272604 490616 272610
rect 490564 272546 490616 272552
rect 493060 272542 493088 313942
rect 493336 309134 493364 316814
rect 493612 316674 493640 322102
rect 493980 318102 494008 322116
rect 493968 318096 494020 318102
rect 493968 318038 494020 318044
rect 493600 316668 493652 316674
rect 493600 316610 493652 316616
rect 494152 316668 494204 316674
rect 494152 316610 494204 316616
rect 493152 309106 493364 309134
rect 493152 280906 493180 309106
rect 493140 280900 493192 280906
rect 493140 280842 493192 280848
rect 493048 272536 493100 272542
rect 493048 272478 493100 272484
rect 490288 271312 490340 271318
rect 490288 271254 490340 271260
rect 490012 271244 490064 271250
rect 490012 271186 490064 271192
rect 488908 271176 488960 271182
rect 488908 271118 488960 271124
rect 494164 269958 494192 316610
rect 494256 282266 494284 322116
rect 494244 282260 494296 282266
rect 494244 282202 494296 282208
rect 494532 274106 494560 322116
rect 494808 318170 494836 322116
rect 494992 322102 495098 322130
rect 495268 322102 495374 322130
rect 494796 318164 494848 318170
rect 494796 318106 494848 318112
rect 494992 313993 495020 322102
rect 495268 316674 495296 322102
rect 495532 319116 495584 319122
rect 495532 319058 495584 319064
rect 495256 316668 495308 316674
rect 495256 316610 495308 316616
rect 494978 313984 495034 313993
rect 494978 313919 495034 313928
rect 494520 274100 494572 274106
rect 494520 274042 494572 274048
rect 486424 269952 486476 269958
rect 486424 269894 486476 269900
rect 494152 269952 494204 269958
rect 494152 269894 494204 269900
rect 495544 268530 495572 319058
rect 495636 318102 495664 322116
rect 495624 318096 495676 318102
rect 495624 318038 495676 318044
rect 495912 316878 495940 322116
rect 496096 322102 496202 322130
rect 496372 322102 496478 322130
rect 496648 322102 496754 322130
rect 495900 316872 495952 316878
rect 495900 316814 495952 316820
rect 496096 316690 496124 322102
rect 496372 319122 496400 322102
rect 496360 319116 496412 319122
rect 496360 319058 496412 319064
rect 495820 316662 496124 316690
rect 495820 314022 495848 316662
rect 496648 316034 496676 322102
rect 496912 319252 496964 319258
rect 496912 319194 496964 319200
rect 496096 316006 496676 316034
rect 496096 315450 496124 316006
rect 496084 315444 496136 315450
rect 496084 315386 496136 315392
rect 495808 314016 495860 314022
rect 495808 313958 495860 313964
rect 496924 271182 496952 319194
rect 497016 283694 497044 322116
rect 497292 319433 497320 322116
rect 497476 322102 497582 322130
rect 497752 322102 497858 322130
rect 498028 322102 498134 322130
rect 497278 319424 497334 319433
rect 497278 319359 497334 319368
rect 497476 319258 497504 322102
rect 497464 319252 497516 319258
rect 497464 319194 497516 319200
rect 497752 319104 497780 322102
rect 497200 319076 497780 319104
rect 497004 283688 497056 283694
rect 497004 283630 497056 283636
rect 497200 273970 497228 319076
rect 498028 316034 498056 322102
rect 498396 316946 498424 322116
rect 498580 322102 498686 322130
rect 498856 322102 498962 322130
rect 499132 322102 499238 322130
rect 499408 322102 499514 322130
rect 498580 319104 498608 322102
rect 498488 319076 498608 319104
rect 498384 316940 498436 316946
rect 498384 316882 498436 316888
rect 498488 316034 498516 319076
rect 498568 318980 498620 318986
rect 498568 318922 498620 318928
rect 497476 316006 498056 316034
rect 498304 316006 498516 316034
rect 497476 275330 497504 316006
rect 497464 275324 497516 275330
rect 497464 275266 497516 275272
rect 497188 273964 497240 273970
rect 497188 273906 497240 273912
rect 498304 271250 498332 316006
rect 498580 272542 498608 318922
rect 498856 276826 498884 322102
rect 499132 291718 499160 322102
rect 499408 318986 499436 322102
rect 499672 319116 499724 319122
rect 499672 319058 499724 319064
rect 499396 318980 499448 318986
rect 499396 318922 499448 318928
rect 499120 291712 499172 291718
rect 499120 291654 499172 291660
rect 498844 276820 498896 276826
rect 498844 276762 498896 276768
rect 498568 272536 498620 272542
rect 498568 272478 498620 272484
rect 498292 271244 498344 271250
rect 498292 271186 498344 271192
rect 496912 271176 496964 271182
rect 496912 271118 496964 271124
rect 499684 268598 499712 319058
rect 499776 315518 499804 322116
rect 500052 317014 500080 322116
rect 500328 319598 500356 322116
rect 500512 322102 500618 322130
rect 500788 322102 500894 322130
rect 500316 319592 500368 319598
rect 500316 319534 500368 319540
rect 500040 317008 500092 317014
rect 500040 316950 500092 316956
rect 500512 316034 500540 322102
rect 500788 319122 500816 322102
rect 501052 319252 501104 319258
rect 501052 319194 501104 319200
rect 500776 319116 500828 319122
rect 500776 319058 500828 319064
rect 499960 316006 500540 316034
rect 499764 315512 499816 315518
rect 499764 315454 499816 315460
rect 499960 278050 499988 316006
rect 501064 279478 501092 319194
rect 501156 311302 501184 322116
rect 501432 319734 501460 322116
rect 501616 322102 501722 322130
rect 501892 322102 501998 322130
rect 502168 322102 502274 322130
rect 501420 319728 501472 319734
rect 501420 319670 501472 319676
rect 501616 319258 501644 322102
rect 501604 319252 501656 319258
rect 501604 319194 501656 319200
rect 501892 319138 501920 322102
rect 501340 319110 501920 319138
rect 501144 311296 501196 311302
rect 501144 311238 501196 311244
rect 501340 285054 501368 319110
rect 502168 316034 502196 322102
rect 502536 319530 502564 322116
rect 502720 322102 502826 322130
rect 502996 322102 503102 322130
rect 503272 322102 503378 322130
rect 503548 322102 503654 322130
rect 502524 319524 502576 319530
rect 502524 319466 502576 319472
rect 502720 319410 502748 322102
rect 502352 319382 502748 319410
rect 502352 316810 502380 319382
rect 502996 319274 503024 322102
rect 502444 319246 503024 319274
rect 502340 316804 502392 316810
rect 502340 316746 502392 316752
rect 501616 316006 502196 316034
rect 501616 314090 501644 316006
rect 501604 314084 501656 314090
rect 501604 314026 501656 314032
rect 502444 301578 502472 319246
rect 503272 319138 503300 322102
rect 502720 319110 503300 319138
rect 502432 301572 502484 301578
rect 502432 301514 502484 301520
rect 502720 298042 502748 319110
rect 503548 316034 503576 322102
rect 502996 316006 503576 316034
rect 502996 315382 503024 316006
rect 502984 315376 503036 315382
rect 502984 315318 503036 315324
rect 503916 313954 503944 322116
rect 504088 322108 504140 322114
rect 504088 322050 504140 322056
rect 504100 321910 504128 322050
rect 504088 321904 504140 321910
rect 504088 321846 504140 321852
rect 504088 319116 504140 319122
rect 504088 319058 504140 319064
rect 503904 313948 503956 313954
rect 503904 313890 503956 313896
rect 502708 298036 502760 298042
rect 502708 297978 502760 297984
rect 501328 285048 501380 285054
rect 501328 284990 501380 284996
rect 501052 279472 501104 279478
rect 501052 279414 501104 279420
rect 499948 278044 500000 278050
rect 499948 277986 500000 277992
rect 499672 268592 499724 268598
rect 499672 268534 499724 268540
rect 475384 268524 475436 268530
rect 475384 268466 475436 268472
rect 495532 268524 495584 268530
rect 495532 268466 495584 268472
rect 504100 268394 504128 319058
rect 504192 311234 504220 322116
rect 504376 322102 504482 322130
rect 504376 315314 504404 322102
rect 504744 316742 504772 322116
rect 504928 322102 505034 322130
rect 505204 322102 505310 322130
rect 504928 319122 504956 322102
rect 504916 319116 504968 319122
rect 504916 319058 504968 319064
rect 504732 316736 504784 316742
rect 504732 316678 504784 316684
rect 504364 315308 504416 315314
rect 504364 315250 504416 315256
rect 504180 311228 504232 311234
rect 504180 311170 504232 311176
rect 505204 268462 505232 322102
rect 507032 321020 507084 321026
rect 507032 320962 507084 320968
rect 507044 304434 507072 320962
rect 507032 304428 507084 304434
rect 507032 304370 507084 304376
rect 507136 286822 507164 322487
rect 507216 322244 507268 322250
rect 507216 322186 507268 322192
rect 507124 286816 507176 286822
rect 507124 286758 507176 286764
rect 507228 286754 507256 322186
rect 507320 289678 507348 322623
rect 507492 322584 507544 322590
rect 507492 322526 507544 322532
rect 507400 321972 507452 321978
rect 507400 321914 507452 321920
rect 507412 291786 507440 321914
rect 507504 292398 507532 322526
rect 507584 320816 507636 320822
rect 507584 320758 507636 320764
rect 507674 320784 507730 320793
rect 507596 292534 507624 320758
rect 507674 320719 507730 320728
rect 507768 320748 507820 320754
rect 507584 292528 507636 292534
rect 507584 292470 507636 292476
rect 507688 292466 507716 320719
rect 507768 320690 507820 320696
rect 507780 297770 507808 320690
rect 509344 300762 509372 366959
rect 509422 358864 509478 358873
rect 509422 358799 509478 358808
rect 509436 300830 509464 358799
rect 509514 349480 509570 349489
rect 509514 349415 509570 349424
rect 509424 300824 509476 300830
rect 509424 300766 509476 300772
rect 509332 300756 509384 300762
rect 509332 300698 509384 300704
rect 507768 297764 507820 297770
rect 507768 297706 507820 297712
rect 509528 295254 509556 349415
rect 509620 322590 509648 372399
rect 509790 333160 509846 333169
rect 509790 333095 509846 333104
rect 509698 326088 509754 326097
rect 509698 326023 509754 326032
rect 509608 322584 509660 322590
rect 509608 322526 509660 322532
rect 509712 303113 509740 326023
rect 509804 321978 509832 333095
rect 509792 321972 509844 321978
rect 509792 321914 509844 321920
rect 509896 321910 509924 418134
rect 510710 368928 510766 368937
rect 510710 368863 510766 368872
rect 510618 366752 510674 366761
rect 510618 366687 510674 366696
rect 510066 333024 510122 333033
rect 510066 332959 510122 332968
rect 509884 321904 509936 321910
rect 509884 321846 509936 321852
rect 510080 320754 510108 332959
rect 510158 329216 510214 329225
rect 510158 329151 510214 329160
rect 510172 322969 510200 329151
rect 510250 328128 510306 328137
rect 510250 328063 510306 328072
rect 510158 322960 510214 322969
rect 510158 322895 510214 322904
rect 510068 320748 510120 320754
rect 510068 320690 510120 320696
rect 509698 303104 509754 303113
rect 509698 303039 509754 303048
rect 510264 300121 510292 328063
rect 510528 323604 510580 323610
rect 510528 323546 510580 323552
rect 510540 319870 510568 323546
rect 510528 319864 510580 319870
rect 510528 319806 510580 319812
rect 510250 300112 510306 300121
rect 510250 300047 510306 300056
rect 509516 295248 509568 295254
rect 509516 295190 509568 295196
rect 507676 292460 507728 292466
rect 507676 292402 507728 292408
rect 507492 292392 507544 292398
rect 507492 292334 507544 292340
rect 507400 291780 507452 291786
rect 507400 291722 507452 291728
rect 507308 289672 507360 289678
rect 507308 289614 507360 289620
rect 510632 289542 510660 366687
rect 510724 300490 510752 368863
rect 510802 360768 510858 360777
rect 510802 360703 510858 360712
rect 510816 300694 510844 360703
rect 510894 355872 510950 355881
rect 510894 355807 510950 355816
rect 510908 303482 510936 355807
rect 510986 352608 511042 352617
rect 510986 352543 511042 352552
rect 510896 303476 510948 303482
rect 510896 303418 510948 303424
rect 511000 303414 511028 352543
rect 511170 342816 511226 342825
rect 511170 342751 511226 342760
rect 510988 303408 511040 303414
rect 510988 303350 511040 303356
rect 511184 302977 511212 342751
rect 511276 322114 511304 576846
rect 511356 524476 511408 524482
rect 511356 524418 511408 524424
rect 511264 322108 511316 322114
rect 511264 322050 511316 322056
rect 511368 321094 511396 524418
rect 513392 387122 513420 600086
rect 519544 536852 519596 536858
rect 519544 536794 519596 536800
rect 518164 484424 518216 484430
rect 518164 484366 518216 484372
rect 516784 470620 516836 470626
rect 516784 470562 516836 470568
rect 515404 464432 515456 464438
rect 515404 464374 515456 464380
rect 513380 387116 513432 387122
rect 513380 387058 513432 387064
rect 512184 386572 512236 386578
rect 512184 386514 512236 386520
rect 512000 386436 512052 386442
rect 512000 386378 512052 386384
rect 512012 378185 512040 386378
rect 512092 385076 512144 385082
rect 512092 385018 512144 385024
rect 512104 380458 512132 385018
rect 512092 380452 512144 380458
rect 512092 380394 512144 380400
rect 512090 380352 512146 380361
rect 512090 380287 512146 380296
rect 512104 380186 512132 380287
rect 512092 380180 512144 380186
rect 512092 380122 512144 380128
rect 512196 378842 512224 386514
rect 512276 386504 512328 386510
rect 512276 386446 512328 386452
rect 512104 378814 512224 378842
rect 511998 378176 512054 378185
rect 511998 378111 512054 378120
rect 512104 377641 512132 378814
rect 512182 378720 512238 378729
rect 512182 378655 512238 378664
rect 512196 378350 512224 378655
rect 512184 378344 512236 378350
rect 512184 378286 512236 378292
rect 512090 377632 512146 377641
rect 512090 377567 512146 377576
rect 512182 376544 512238 376553
rect 512182 376479 512238 376488
rect 511998 371104 512054 371113
rect 511998 371039 512054 371048
rect 512012 370122 512040 371039
rect 512090 370560 512146 370569
rect 512090 370495 512146 370504
rect 512000 370116 512052 370122
rect 512000 370058 512052 370064
rect 512104 369986 512132 370495
rect 512092 369980 512144 369986
rect 512092 369922 512144 369928
rect 512090 364576 512146 364585
rect 512090 364511 512092 364520
rect 512144 364511 512146 364520
rect 512092 364482 512144 364488
rect 511998 364032 512054 364041
rect 511998 363967 512054 363976
rect 512012 363050 512040 363967
rect 512000 363044 512052 363050
rect 512000 362986 512052 362992
rect 511998 362400 512054 362409
rect 511998 362335 512054 362344
rect 512012 362234 512040 362335
rect 512000 362228 512052 362234
rect 512000 362170 512052 362176
rect 511998 358592 512054 358601
rect 511998 358527 512054 358536
rect 511538 343360 511594 343369
rect 511538 343295 511594 343304
rect 511356 321088 511408 321094
rect 511356 321030 511408 321036
rect 511170 302968 511226 302977
rect 511170 302903 511226 302912
rect 510804 300688 510856 300694
rect 510804 300630 510856 300636
rect 510712 300484 510764 300490
rect 510712 300426 510764 300432
rect 511552 297702 511580 343295
rect 511908 324352 511960 324358
rect 511908 324294 511960 324300
rect 511920 319802 511948 324294
rect 511908 319796 511960 319802
rect 511908 319738 511960 319744
rect 511540 297696 511592 297702
rect 511540 297638 511592 297644
rect 510620 289536 510672 289542
rect 510620 289478 510672 289484
rect 507216 286748 507268 286754
rect 507216 286690 507268 286696
rect 512012 276690 512040 358527
rect 512090 358048 512146 358057
rect 512090 357983 512146 357992
rect 512104 357678 512132 357983
rect 512092 357672 512144 357678
rect 512092 357614 512144 357620
rect 512090 357504 512146 357513
rect 512090 357439 512092 357448
rect 512144 357439 512146 357448
rect 512092 357410 512144 357416
rect 512090 356416 512146 356425
rect 512090 356351 512092 356360
rect 512144 356351 512146 356360
rect 512092 356322 512144 356328
rect 512090 354240 512146 354249
rect 512090 354175 512146 354184
rect 512104 353802 512132 354175
rect 512092 353796 512144 353802
rect 512092 353738 512144 353744
rect 512090 350976 512146 350985
rect 512090 350911 512146 350920
rect 512104 350810 512132 350911
rect 512092 350804 512144 350810
rect 512092 350746 512144 350752
rect 512090 349344 512146 349353
rect 512090 349279 512146 349288
rect 512104 349246 512132 349279
rect 512092 349240 512144 349246
rect 512092 349182 512144 349188
rect 512090 346080 512146 346089
rect 512090 346015 512146 346024
rect 512104 345982 512132 346015
rect 512092 345976 512144 345982
rect 512092 345918 512144 345924
rect 512090 345536 512146 345545
rect 512090 345471 512146 345480
rect 512000 276684 512052 276690
rect 512000 276626 512052 276632
rect 512104 269822 512132 345471
rect 512196 304298 512224 376479
rect 512288 376009 512316 386446
rect 512734 384704 512790 384713
rect 512734 384639 512790 384648
rect 512748 383790 512776 384639
rect 513286 384160 513342 384169
rect 513286 384095 513342 384104
rect 512736 383784 512788 383790
rect 512736 383726 512788 383732
rect 513300 383722 513328 384095
rect 513288 383716 513340 383722
rect 513288 383658 513340 383664
rect 512918 383616 512974 383625
rect 512918 383551 512974 383560
rect 512932 382294 512960 383551
rect 513286 383072 513342 383081
rect 513286 383007 513342 383016
rect 513194 382528 513250 382537
rect 513194 382463 513196 382472
rect 513248 382463 513250 382472
rect 513196 382434 513248 382440
rect 513300 382430 513328 383007
rect 513288 382424 513340 382430
rect 513288 382366 513340 382372
rect 512920 382288 512972 382294
rect 512920 382230 512972 382236
rect 512366 381984 512422 381993
rect 512366 381919 512422 381928
rect 512380 381138 512408 381919
rect 513286 381440 513342 381449
rect 513286 381375 513342 381384
rect 512368 381132 512420 381138
rect 512368 381074 512420 381080
rect 513300 380934 513328 381375
rect 513288 380928 513340 380934
rect 512366 380896 512422 380905
rect 513288 380870 513340 380876
rect 512366 380831 512422 380840
rect 512380 376038 512408 380831
rect 512460 380452 512512 380458
rect 512460 380394 512512 380400
rect 512368 376032 512420 376038
rect 512274 376000 512330 376009
rect 512368 375974 512420 375980
rect 512274 375935 512330 375944
rect 512472 374921 512500 380394
rect 514116 380180 514168 380186
rect 514116 380122 514168 380128
rect 512826 379808 512882 379817
rect 512826 379743 512882 379752
rect 512840 379574 512868 379743
rect 512828 379568 512880 379574
rect 512828 379510 512880 379516
rect 513286 379264 513342 379273
rect 513286 379199 513342 379208
rect 513300 378282 513328 379199
rect 513288 378276 513340 378282
rect 513288 378218 513340 378224
rect 514024 378208 514076 378214
rect 514024 378150 514076 378156
rect 513194 377088 513250 377097
rect 513194 377023 513250 377032
rect 513208 376922 513236 377023
rect 513196 376916 513248 376922
rect 513196 376858 513248 376864
rect 513286 375456 513342 375465
rect 513342 375414 513420 375442
rect 513286 375391 513342 375400
rect 512458 374912 512514 374921
rect 512458 374847 512514 374856
rect 512734 374368 512790 374377
rect 512734 374303 512790 374312
rect 512748 374202 512776 374303
rect 512736 374196 512788 374202
rect 512736 374138 512788 374144
rect 513392 373994 513420 375414
rect 513392 373966 513512 373994
rect 512826 373824 512882 373833
rect 512826 373759 512882 373768
rect 512840 372706 512868 373759
rect 513286 373280 513342 373289
rect 513286 373215 513342 373224
rect 512828 372700 512880 372706
rect 512828 372642 512880 372648
rect 513300 372638 513328 373215
rect 513288 372632 513340 372638
rect 513288 372574 513340 372580
rect 512550 372192 512606 372201
rect 512550 372127 512606 372136
rect 512274 371648 512330 371657
rect 512274 371583 512330 371592
rect 512288 305726 512316 371583
rect 512564 371278 512592 372127
rect 512552 371272 512604 371278
rect 512552 371214 512604 371220
rect 513288 370048 513340 370054
rect 513286 370016 513288 370025
rect 513340 370016 513342 370025
rect 513286 369951 513342 369960
rect 513010 369472 513066 369481
rect 513010 369407 513066 369416
rect 513024 368626 513052 369407
rect 513012 368620 513064 368626
rect 513012 368562 513064 368568
rect 512366 368384 512422 368393
rect 512366 368319 512422 368328
rect 512276 305720 512328 305726
rect 512276 305662 512328 305668
rect 512184 304292 512236 304298
rect 512184 304234 512236 304240
rect 512380 302938 512408 368319
rect 512642 367840 512698 367849
rect 512642 367775 512698 367784
rect 512656 367266 512684 367775
rect 512644 367260 512696 367266
rect 512644 367202 512696 367208
rect 512458 366208 512514 366217
rect 512458 366143 512514 366152
rect 512472 365906 512500 366143
rect 512460 365900 512512 365906
rect 512460 365842 512512 365848
rect 512458 365120 512514 365129
rect 512458 365055 512514 365064
rect 512368 302932 512420 302938
rect 512368 302874 512420 302880
rect 512472 301510 512500 365055
rect 513286 363488 513342 363497
rect 513286 363423 513342 363432
rect 513300 363118 513328 363423
rect 513288 363112 513340 363118
rect 513288 363054 513340 363060
rect 513286 362944 513342 362953
rect 513286 362879 513342 362888
rect 513300 362098 513328 362879
rect 513288 362092 513340 362098
rect 513288 362034 513340 362040
rect 513102 361856 513158 361865
rect 513102 361791 513104 361800
rect 513156 361791 513158 361800
rect 513104 361762 513156 361768
rect 513286 361312 513342 361321
rect 513286 361247 513342 361256
rect 513300 360330 513328 361247
rect 513288 360324 513340 360330
rect 513288 360266 513340 360272
rect 512550 360224 512606 360233
rect 512550 360159 512606 360168
rect 512564 305658 512592 360159
rect 513286 359680 513342 359689
rect 513286 359615 513342 359624
rect 513300 358902 513328 359615
rect 513288 358896 513340 358902
rect 513288 358838 513340 358844
rect 512734 356960 512790 356969
rect 512734 356895 512790 356904
rect 512748 356182 512776 356895
rect 512736 356176 512788 356182
rect 512736 356118 512788 356124
rect 513194 355328 513250 355337
rect 513194 355263 513250 355272
rect 513208 354754 513236 355263
rect 513288 354816 513340 354822
rect 513286 354784 513288 354793
rect 513340 354784 513342 354793
rect 513196 354748 513248 354754
rect 513286 354719 513342 354728
rect 513196 354690 513248 354696
rect 513286 353696 513342 353705
rect 513286 353631 513342 353640
rect 513300 353326 513328 353631
rect 513288 353320 513340 353326
rect 513288 353262 513340 353268
rect 512918 353152 512974 353161
rect 512918 353087 512974 353096
rect 512932 352170 512960 353087
rect 512920 352164 512972 352170
rect 512920 352106 512972 352112
rect 513286 352064 513342 352073
rect 513286 351999 513342 352008
rect 513300 351966 513328 351999
rect 513288 351960 513340 351966
rect 513288 351902 513340 351908
rect 512826 351520 512882 351529
rect 512826 351455 512828 351464
rect 512880 351455 512882 351464
rect 512828 351426 512880 351432
rect 513010 350432 513066 350441
rect 513010 350367 513066 350376
rect 513024 349314 513052 350367
rect 513012 349308 513064 349314
rect 513012 349250 513064 349256
rect 512826 348800 512882 348809
rect 512826 348735 512882 348744
rect 512840 347954 512868 348735
rect 512918 348256 512974 348265
rect 512918 348191 512974 348200
rect 512828 347948 512880 347954
rect 512828 347890 512880 347896
rect 512932 347818 512960 348191
rect 512920 347812 512972 347818
rect 512920 347754 512972 347760
rect 512642 347712 512698 347721
rect 512642 347647 512698 347656
rect 512656 346458 512684 347647
rect 513286 347168 513342 347177
rect 513286 347103 513342 347112
rect 513300 346730 513328 347103
rect 513288 346724 513340 346730
rect 513288 346666 513340 346672
rect 512826 346624 512882 346633
rect 512826 346559 512828 346568
rect 512880 346559 512882 346568
rect 512828 346530 512880 346536
rect 512644 346452 512696 346458
rect 512644 346394 512696 346400
rect 513286 344992 513342 345001
rect 513286 344927 513342 344936
rect 512642 344448 512698 344457
rect 512642 344383 512698 344392
rect 512656 344282 512684 344383
rect 512644 344276 512696 344282
rect 512644 344218 512696 344224
rect 513300 344010 513328 344927
rect 513288 344004 513340 344010
rect 513288 343946 513340 343952
rect 512826 343904 512882 343913
rect 512826 343839 512828 343848
rect 512880 343839 512882 343848
rect 512828 343810 512880 343816
rect 512642 342272 512698 342281
rect 512642 342207 512698 342216
rect 512656 305833 512684 342207
rect 513286 341728 513342 341737
rect 513286 341663 513342 341672
rect 513300 341290 513328 341663
rect 513288 341284 513340 341290
rect 513288 341226 513340 341232
rect 513010 341184 513066 341193
rect 513010 341119 513066 341128
rect 513024 341018 513052 341119
rect 513012 341012 513064 341018
rect 513012 340954 513064 340960
rect 513194 340640 513250 340649
rect 513194 340575 513250 340584
rect 513012 339584 513064 339590
rect 513010 339552 513012 339561
rect 513064 339552 513066 339561
rect 513208 339522 513236 340575
rect 513286 340096 513342 340105
rect 513286 340031 513342 340040
rect 513300 339930 513328 340031
rect 513288 339924 513340 339930
rect 513288 339866 513340 339872
rect 513010 339487 513066 339496
rect 513196 339516 513248 339522
rect 513196 339458 513248 339464
rect 513194 339008 513250 339017
rect 513194 338943 513250 338952
rect 513208 338162 513236 338943
rect 513286 338464 513342 338473
rect 513286 338399 513342 338408
rect 513300 338298 513328 338399
rect 513288 338292 513340 338298
rect 513288 338234 513340 338240
rect 513196 338156 513248 338162
rect 513196 338098 513248 338104
rect 513194 337920 513250 337929
rect 513194 337855 513250 337864
rect 513208 337482 513236 337855
rect 513196 337476 513248 337482
rect 513196 337418 513248 337424
rect 513194 337376 513250 337385
rect 513194 337311 513250 337320
rect 513208 336802 513236 337311
rect 513288 336864 513340 336870
rect 513286 336832 513288 336841
rect 513340 336832 513342 336841
rect 513196 336796 513248 336802
rect 513286 336767 513342 336776
rect 513196 336738 513248 336744
rect 513194 336288 513250 336297
rect 513194 336223 513250 336232
rect 513208 335850 513236 336223
rect 513196 335844 513248 335850
rect 513196 335786 513248 335792
rect 513286 335744 513342 335753
rect 513286 335679 513342 335688
rect 513300 335374 513328 335679
rect 513288 335368 513340 335374
rect 513288 335310 513340 335316
rect 513194 335200 513250 335209
rect 513194 335135 513250 335144
rect 513208 334354 513236 335135
rect 513196 334348 513248 334354
rect 513196 334290 513248 334296
rect 513286 334112 513342 334121
rect 513286 334047 513342 334056
rect 513300 334014 513328 334047
rect 513288 334008 513340 334014
rect 513288 333950 513340 333956
rect 513286 331936 513342 331945
rect 513342 331894 513420 331922
rect 513286 331871 513342 331880
rect 512734 330848 512790 330857
rect 512734 330783 512790 330792
rect 512748 330138 512776 330783
rect 512736 330132 512788 330138
rect 512736 330074 512788 330080
rect 512734 325408 512790 325417
rect 512734 325343 512790 325352
rect 512642 305824 512698 305833
rect 512642 305759 512698 305768
rect 512552 305652 512604 305658
rect 512552 305594 512604 305600
rect 512748 304366 512776 325343
rect 513392 320822 513420 331894
rect 513380 320816 513432 320822
rect 513380 320758 513432 320764
rect 512736 304360 512788 304366
rect 512736 304302 512788 304308
rect 512460 301504 512512 301510
rect 512460 301446 512512 301452
rect 513484 300286 513512 373966
rect 513562 365664 513618 365673
rect 513562 365599 513618 365608
rect 513576 300626 513604 365599
rect 513748 362228 513800 362234
rect 513748 362170 513800 362176
rect 513656 356380 513708 356386
rect 513656 356322 513708 356328
rect 513564 300620 513616 300626
rect 513564 300562 513616 300568
rect 513472 300280 513524 300286
rect 513472 300222 513524 300228
rect 513668 295186 513696 356322
rect 513760 300558 513788 362170
rect 513840 357468 513892 357474
rect 513840 357410 513892 357416
rect 513852 303006 513880 357410
rect 513932 349240 513984 349246
rect 513932 349182 513984 349188
rect 513944 303346 513972 349182
rect 514036 322182 514064 378150
rect 514128 358834 514156 380122
rect 514208 370116 514260 370122
rect 514208 370058 514260 370064
rect 514116 358828 514168 358834
rect 514116 358770 514168 358776
rect 514116 345976 514168 345982
rect 514116 345918 514168 345924
rect 514024 322176 514076 322182
rect 514024 322118 514076 322124
rect 513932 303340 513984 303346
rect 513932 303282 513984 303288
rect 514128 303278 514156 345918
rect 514116 303272 514168 303278
rect 514116 303214 514168 303220
rect 513840 303000 513892 303006
rect 513840 302942 513892 302948
rect 513748 300552 513800 300558
rect 513748 300494 513800 300500
rect 513656 295180 513708 295186
rect 513656 295122 513708 295128
rect 514220 292262 514248 370058
rect 514944 369980 514996 369986
rect 514944 369922 514996 369928
rect 514852 364540 514904 364546
rect 514852 364482 514904 364488
rect 514760 330132 514812 330138
rect 514760 330074 514812 330080
rect 514772 322250 514800 330074
rect 514760 322244 514812 322250
rect 514760 322186 514812 322192
rect 514864 295322 514892 364482
rect 514956 300354 514984 369922
rect 515036 363044 515088 363050
rect 515036 362986 515088 362992
rect 515048 300422 515076 362986
rect 515128 353796 515180 353802
rect 515128 353738 515180 353744
rect 515140 303074 515168 353738
rect 515220 350804 515272 350810
rect 515220 350746 515272 350752
rect 515232 303142 515260 350746
rect 515312 346452 515364 346458
rect 515312 346394 515364 346400
rect 515324 303210 515352 346394
rect 515416 320006 515444 464374
rect 515496 381132 515548 381138
rect 515496 381074 515548 381080
rect 515508 358494 515536 381074
rect 516140 374196 516192 374202
rect 516140 374138 516192 374144
rect 515588 365900 515640 365906
rect 515588 365842 515640 365848
rect 515496 358488 515548 358494
rect 515496 358430 515548 358436
rect 515496 344276 515548 344282
rect 515496 344218 515548 344224
rect 515404 320000 515456 320006
rect 515404 319942 515456 319948
rect 515312 303204 515364 303210
rect 515312 303146 515364 303152
rect 515220 303136 515272 303142
rect 515220 303078 515272 303084
rect 515128 303068 515180 303074
rect 515128 303010 515180 303016
rect 515508 302841 515536 344218
rect 515494 302832 515550 302841
rect 515494 302767 515550 302776
rect 515036 300416 515088 300422
rect 515036 300358 515088 300364
rect 514944 300348 514996 300354
rect 514944 300290 514996 300296
rect 514852 295316 514904 295322
rect 514852 295258 514904 295264
rect 515600 294574 515628 365842
rect 515588 294568 515640 294574
rect 515588 294510 515640 294516
rect 514208 292256 514260 292262
rect 514208 292198 514260 292204
rect 516152 292194 516180 374138
rect 516324 352164 516376 352170
rect 516324 352106 516376 352112
rect 516232 347948 516284 347954
rect 516232 347890 516284 347896
rect 516140 292188 516192 292194
rect 516140 292130 516192 292136
rect 516244 289610 516272 347890
rect 516336 294846 516364 352106
rect 516508 347812 516560 347818
rect 516508 347754 516560 347760
rect 516416 343868 516468 343874
rect 516416 343810 516468 343816
rect 516324 294840 516376 294846
rect 516324 294782 516376 294788
rect 516232 289604 516284 289610
rect 516232 289546 516284 289552
rect 516428 289270 516456 343810
rect 516520 294914 516548 347754
rect 516600 341012 516652 341018
rect 516600 340954 516652 340960
rect 516612 297906 516640 340954
rect 516692 339584 516744 339590
rect 516692 339526 516744 339532
rect 516600 297900 516652 297906
rect 516600 297842 516652 297848
rect 516704 297838 516732 339526
rect 516796 321842 516824 470562
rect 517520 376916 517572 376922
rect 517520 376858 517572 376864
rect 516876 361820 516928 361826
rect 516876 361762 516928 361768
rect 516784 321836 516836 321842
rect 516784 321778 516836 321784
rect 516888 321026 516916 361762
rect 516968 335844 517020 335850
rect 516968 335786 517020 335792
rect 516876 321020 516928 321026
rect 516876 320962 516928 320968
rect 516692 297832 516744 297838
rect 516692 297774 516744 297780
rect 516980 297498 517008 335786
rect 517532 297566 517560 376858
rect 517612 372700 517664 372706
rect 517612 372642 517664 372648
rect 517624 300150 517652 372642
rect 517704 371272 517756 371278
rect 517704 371214 517756 371220
rect 517716 300218 517744 371214
rect 517888 351484 517940 351490
rect 517888 351426 517940 351432
rect 517796 346724 517848 346730
rect 517796 346666 517848 346672
rect 517704 300212 517756 300218
rect 517704 300154 517756 300160
rect 517612 300144 517664 300150
rect 517612 300086 517664 300092
rect 517520 297560 517572 297566
rect 517520 297502 517572 297508
rect 516968 297492 517020 297498
rect 516968 297434 517020 297440
rect 516508 294908 516560 294914
rect 516508 294850 516560 294856
rect 517808 289338 517836 346666
rect 517900 294642 517928 351426
rect 517980 346588 518032 346594
rect 517980 346530 518032 346536
rect 517992 297634 518020 346530
rect 518072 344004 518124 344010
rect 518072 343946 518124 343952
rect 517980 297628 518032 297634
rect 517980 297570 518032 297576
rect 518084 297430 518112 343946
rect 518176 322046 518204 484366
rect 518348 382492 518400 382498
rect 518348 382434 518400 382440
rect 518256 363112 518308 363118
rect 518256 363054 518308 363060
rect 518164 322040 518216 322046
rect 518164 321982 518216 321988
rect 518268 320958 518296 363054
rect 518360 358630 518388 382434
rect 518900 368620 518952 368626
rect 518900 368562 518952 368568
rect 518348 358624 518400 358630
rect 518348 358566 518400 358572
rect 518348 337476 518400 337482
rect 518348 337418 518400 337424
rect 518256 320952 518308 320958
rect 518256 320894 518308 320900
rect 518360 300257 518388 337418
rect 518346 300248 518402 300257
rect 518346 300183 518402 300192
rect 518072 297424 518124 297430
rect 518072 297366 518124 297372
rect 517888 294636 517940 294642
rect 517888 294578 517940 294584
rect 518912 291990 518940 368562
rect 518992 362092 519044 362098
rect 518992 362034 519044 362040
rect 519004 295118 519032 362034
rect 519176 358896 519228 358902
rect 519176 358838 519228 358844
rect 519084 353320 519136 353326
rect 519084 353262 519136 353268
rect 518992 295112 519044 295118
rect 518992 295054 519044 295060
rect 518900 291984 518952 291990
rect 518900 291926 518952 291932
rect 519096 289814 519124 353262
rect 519188 295050 519216 358838
rect 519268 357672 519320 357678
rect 519268 357614 519320 357620
rect 519176 295044 519228 295050
rect 519176 294986 519228 294992
rect 519280 294778 519308 357614
rect 519452 354816 519504 354822
rect 519452 354758 519504 354764
rect 519360 349308 519412 349314
rect 519360 349250 519412 349256
rect 519268 294772 519320 294778
rect 519268 294714 519320 294720
rect 519084 289808 519136 289814
rect 519084 289750 519136 289756
rect 519372 289474 519400 349250
rect 519464 294710 519492 354758
rect 519556 319938 519584 536794
rect 520292 520946 520320 600086
rect 520280 520940 520332 520946
rect 520280 520882 520332 520888
rect 525812 464370 525840 600086
rect 538220 515432 538272 515438
rect 538220 515374 538272 515380
rect 535460 512644 535512 512650
rect 535460 512586 535512 512592
rect 532700 508564 532752 508570
rect 532700 508506 532752 508512
rect 529940 505776 529992 505782
rect 529940 505718 529992 505724
rect 529952 480254 529980 505718
rect 532712 480254 532740 508506
rect 535472 480254 535500 512586
rect 538232 480254 538260 515374
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 525800 464364 525852 464370
rect 525800 464306 525852 464312
rect 527640 463004 527692 463010
rect 527640 462946 527692 462952
rect 521752 461644 521804 461650
rect 521752 461586 521804 461592
rect 521764 460972 521792 461586
rect 524432 460970 524722 460986
rect 527652 460972 527680 462946
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542372 464438 542400 702406
rect 559668 699825 559696 703520
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 573364 696992 573416 696998
rect 573364 696934 573416 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 569224 670744 569276 670750
rect 569224 670686 569276 670692
rect 567844 510672 567896 510678
rect 567844 510614 567896 510620
rect 545120 500268 545172 500274
rect 545120 500210 545172 500216
rect 542452 498840 542504 498846
rect 542452 498782 542504 498788
rect 542360 464432 542412 464438
rect 542360 464374 542412 464380
rect 542464 460986 542492 498782
rect 524420 460964 524722 460970
rect 524472 460958 524722 460964
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542386 460958 542492 460986
rect 545132 460986 545160 500210
rect 547880 496120 547932 496126
rect 547880 496062 547932 496068
rect 547892 460986 547920 496062
rect 554136 462460 554188 462466
rect 554136 462402 554188 462408
rect 551192 462392 551244 462398
rect 551192 462334 551244 462340
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 551204 460972 551232 462334
rect 554148 460972 554176 462402
rect 524420 460906 524472 460912
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388890 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 522304 388884 522356 388890
rect 522304 388826 522356 388832
rect 523696 388822 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 527284 425054 527666 425082
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388816 523736 388822
rect 523684 388758 523736 388764
rect 524432 388686 524460 412606
rect 526456 388754 526484 423302
rect 527284 412634 527312 425054
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527192 412606 527312 412634
rect 526444 388748 526496 388754
rect 526444 388690 526496 388696
rect 524420 388680 524472 388686
rect 524420 388622 524472 388628
rect 527192 388618 527220 412606
rect 527180 388612 527232 388618
rect 527180 388554 527232 388560
rect 529216 388482 529244 423574
rect 530596 388550 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 534092 392630 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 393990 534212 412606
rect 535472 395350 535500 412606
rect 536852 396778 536880 412606
rect 538232 398138 538260 412606
rect 539612 399498 539640 412606
rect 539600 399492 539652 399498
rect 539600 399434 539652 399440
rect 538220 398132 538272 398138
rect 538220 398074 538272 398080
rect 536840 396772 536892 396778
rect 536840 396714 536892 396720
rect 535460 395344 535512 395350
rect 535460 395286 535512 395292
rect 534172 393984 534224 393990
rect 534172 393926 534224 393932
rect 534080 392624 534132 392630
rect 534080 392566 534132 392572
rect 542372 389910 542400 412606
rect 543752 391338 543780 412606
rect 546512 400926 546540 412606
rect 557552 402286 557580 442847
rect 557540 402280 557592 402286
rect 557540 402222 557592 402228
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 391332 543792 391338
rect 543740 391274 543792 391280
rect 542360 389904 542412 389910
rect 542360 389846 542412 389852
rect 530584 388544 530636 388550
rect 530584 388486 530636 388492
rect 529204 388476 529256 388482
rect 529204 388418 529256 388424
rect 553952 386640 554004 386646
rect 553952 386582 554004 386588
rect 534724 383784 534776 383790
rect 534724 383726 534776 383732
rect 519636 382424 519688 382430
rect 519636 382366 519688 382372
rect 519648 358698 519676 382366
rect 522304 382288 522356 382294
rect 522304 382230 522356 382236
rect 521660 372632 521712 372638
rect 521660 372574 521712 372580
rect 520280 367260 520332 367266
rect 520280 367202 520332 367208
rect 519636 358692 519688 358698
rect 519636 358634 519688 358640
rect 519636 341284 519688 341290
rect 519636 341226 519688 341232
rect 519544 319932 519596 319938
rect 519544 319874 519596 319880
rect 519452 294704 519504 294710
rect 519452 294646 519504 294652
rect 519360 289468 519412 289474
rect 519360 289410 519412 289416
rect 517796 289332 517848 289338
rect 517796 289274 517848 289280
rect 516416 289264 516468 289270
rect 516416 289206 516468 289212
rect 519648 289134 519676 341226
rect 519728 338292 519780 338298
rect 519728 338234 519780 338240
rect 519740 291922 519768 338234
rect 520292 292058 520320 367202
rect 520372 360324 520424 360330
rect 520372 360266 520424 360272
rect 520384 294982 520412 360266
rect 520556 339924 520608 339930
rect 520556 339866 520608 339872
rect 520464 338156 520516 338162
rect 520464 338098 520516 338104
rect 520372 294976 520424 294982
rect 520372 294918 520424 294924
rect 520280 292052 520332 292058
rect 520280 291994 520332 292000
rect 519728 291916 519780 291922
rect 519728 291858 519780 291864
rect 519636 289128 519688 289134
rect 519636 289070 519688 289076
rect 520476 286482 520504 338098
rect 520568 291854 520596 339866
rect 520648 336864 520700 336870
rect 520648 336806 520700 336812
rect 520660 292126 520688 336806
rect 520740 334348 520792 334354
rect 520740 334290 520792 334296
rect 520752 292330 520780 334290
rect 520740 292324 520792 292330
rect 520740 292266 520792 292272
rect 520648 292120 520700 292126
rect 520648 292062 520700 292068
rect 520556 291848 520608 291854
rect 520556 291790 520608 291796
rect 520464 286476 520516 286482
rect 520464 286418 520516 286424
rect 521672 286346 521700 372574
rect 521752 370048 521804 370054
rect 521752 369990 521804 369996
rect 521764 289202 521792 369990
rect 522316 358562 522344 382230
rect 523684 378344 523736 378350
rect 523684 378286 523736 378292
rect 523696 358970 523724 378286
rect 523684 358964 523736 358970
rect 523684 358906 523736 358912
rect 534736 358902 534764 383726
rect 548524 383716 548576 383722
rect 548524 383658 548576 383664
rect 544384 379568 544436 379574
rect 544384 379510 544436 379516
rect 544396 359106 544424 379510
rect 547144 378276 547196 378282
rect 547144 378218 547196 378224
rect 547156 359242 547184 378218
rect 547144 359236 547196 359242
rect 547144 359178 547196 359184
rect 544384 359100 544436 359106
rect 544384 359042 544436 359048
rect 548536 359038 548564 383658
rect 548616 380928 548668 380934
rect 548616 380870 548668 380876
rect 548628 359174 548656 380870
rect 553964 377890 553992 386582
rect 563428 385144 563480 385150
rect 563428 385086 563480 385092
rect 553964 377862 554438 377890
rect 563440 377876 563468 385086
rect 549904 376032 549956 376038
rect 549904 375974 549956 375980
rect 548616 359168 548668 359174
rect 548616 359110 548668 359116
rect 548524 359032 548576 359038
rect 548524 358974 548576 358980
rect 534724 358896 534776 358902
rect 534724 358838 534776 358844
rect 549916 358766 549944 375974
rect 550836 358970 550864 360060
rect 552308 359242 552336 360060
rect 552296 359236 552348 359242
rect 552296 359178 552348 359184
rect 553780 359106 553808 360060
rect 553768 359100 553820 359106
rect 553768 359042 553820 359048
rect 550824 358964 550876 358970
rect 550824 358906 550876 358912
rect 555252 358834 555280 360060
rect 555240 358828 555292 358834
rect 555240 358770 555292 358776
rect 556724 358766 556752 360060
rect 558196 359174 558224 360060
rect 558184 359168 558236 359174
rect 558184 359110 558236 359116
rect 549904 358760 549956 358766
rect 549904 358702 549956 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 522304 358556 522356 358562
rect 522304 358498 522356 358504
rect 559668 358494 559696 360060
rect 561140 358630 561168 360060
rect 562612 358698 562640 360060
rect 562600 358692 562652 358698
rect 562600 358634 562652 358640
rect 561128 358624 561180 358630
rect 561128 358566 561180 358572
rect 564084 358562 564112 360060
rect 565556 359038 565584 360060
rect 565544 359032 565596 359038
rect 565544 358974 565596 358980
rect 567028 358902 567056 360060
rect 567016 358896 567068 358902
rect 567016 358838 567068 358844
rect 564072 358556 564124 358562
rect 564072 358498 564124 358504
rect 559656 358488 559708 358494
rect 559656 358430 559708 358436
rect 521844 356176 521896 356182
rect 521844 356118 521896 356124
rect 521752 289196 521804 289202
rect 521752 289138 521804 289144
rect 521856 289066 521884 356118
rect 521936 354748 521988 354754
rect 521936 354690 521988 354696
rect 521948 289746 521976 354690
rect 522028 351960 522080 351966
rect 522028 351902 522080 351908
rect 521936 289740 521988 289746
rect 521936 289682 521988 289688
rect 522040 289406 522068 351902
rect 522120 339516 522172 339522
rect 522120 339458 522172 339464
rect 522028 289400 522080 289406
rect 522028 289342 522080 289348
rect 521844 289060 521896 289066
rect 521844 289002 521896 289008
rect 522132 286414 522160 339458
rect 522212 336796 522264 336802
rect 522212 336738 522264 336744
rect 522224 286550 522252 336738
rect 522304 335368 522356 335374
rect 522304 335310 522356 335316
rect 522316 286618 522344 335310
rect 522396 334008 522448 334014
rect 522396 333950 522448 333956
rect 522408 286686 522436 333950
rect 567856 321774 567884 510614
rect 567844 321768 567896 321774
rect 567844 321710 567896 321716
rect 569236 321434 569264 670686
rect 571984 590708 572036 590714
rect 571984 590650 572036 590656
rect 570604 364404 570656 364410
rect 570604 364346 570656 364352
rect 569224 321428 569276 321434
rect 569224 321370 569276 321376
rect 570616 321298 570644 364346
rect 570604 321292 570656 321298
rect 570604 321234 570656 321240
rect 571996 320074 572024 590650
rect 573376 321162 573404 696934
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 578882 644056 578938 644065
rect 578882 643991 578938 644000
rect 576124 630692 576176 630698
rect 576124 630634 576176 630640
rect 574744 430636 574796 430642
rect 574744 430578 574796 430584
rect 574756 321230 574784 430578
rect 576136 321366 576164 630634
rect 576124 321360 576176 321366
rect 576124 321302 576176 321308
rect 574744 321224 574796 321230
rect 574744 321166 574796 321172
rect 573364 321156 573416 321162
rect 573364 321098 573416 321104
rect 578896 320142 578924 643991
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 579632 470626 579660 471407
rect 579620 470620 579672 470626
rect 579620 470562 579672 470568
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579632 430642 579660 431559
rect 579620 430636 579672 430642
rect 579620 430578 579672 430584
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 579632 378214 579660 378383
rect 579620 378208 579672 378214
rect 579620 378150 579672 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580276 323610 580304 683839
rect 580354 617536 580410 617545
rect 580354 617471 580410 617480
rect 580264 323604 580316 323610
rect 580264 323546 580316 323552
rect 580368 321706 580396 617471
rect 580446 564360 580502 564369
rect 580446 564295 580502 564304
rect 580356 321700 580408 321706
rect 580356 321642 580408 321648
rect 580460 321638 580488 564295
rect 580538 458144 580594 458153
rect 580538 458079 580594 458088
rect 580448 321632 580500 321638
rect 580448 321574 580500 321580
rect 580552 320890 580580 458079
rect 580630 404968 580686 404977
rect 580630 404903 580686 404912
rect 580644 321502 580672 404903
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580736 321570 580764 351863
rect 580724 321564 580776 321570
rect 580724 321506 580776 321512
rect 580632 321496 580684 321502
rect 580632 321438 580684 321444
rect 580540 320884 580592 320890
rect 580540 320826 580592 320832
rect 578884 320136 578936 320142
rect 578884 320078 578936 320084
rect 571984 320068 572036 320074
rect 571984 320010 572036 320016
rect 534724 319592 534776 319598
rect 534724 319534 534776 319540
rect 533344 311160 533396 311166
rect 533344 311102 533396 311108
rect 529940 307148 529992 307154
rect 529940 307090 529992 307096
rect 528560 303544 528612 303550
rect 528560 303486 528612 303492
rect 528572 287054 528600 303486
rect 528572 287026 529336 287054
rect 522396 286680 522448 286686
rect 522396 286622 522448 286628
rect 522304 286612 522356 286618
rect 522304 286554 522356 286560
rect 522212 286544 522264 286550
rect 522212 286486 522264 286492
rect 522120 286408 522172 286414
rect 522120 286350 522172 286356
rect 521660 286340 521712 286346
rect 521660 286282 521712 286288
rect 512092 269816 512144 269822
rect 512092 269758 512144 269764
rect 505192 268456 505244 268462
rect 505192 268398 505244 268404
rect 504088 268388 504140 268394
rect 504088 268330 504140 268336
rect 529308 261633 529336 287026
rect 529294 261624 529350 261633
rect 529294 261559 529350 261568
rect 529952 209273 529980 307090
rect 530032 304496 530084 304502
rect 530032 304438 530084 304444
rect 530044 226250 530072 304438
rect 530124 286884 530176 286890
rect 530124 286826 530176 286832
rect 530136 243681 530164 286826
rect 530122 243672 530178 243681
rect 530122 243607 530178 243616
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 479524 200796 479576 200802
rect 479524 200738 479576 200744
rect 461584 163600 461636 163606
rect 461584 163542 461636 163548
rect 460296 157344 460348 157350
rect 460296 157286 460348 157292
rect 461596 41410 461624 163542
rect 461676 160268 461728 160274
rect 461676 160210 461728 160216
rect 461688 143002 461716 160210
rect 461676 142996 461728 143002
rect 461676 142938 461728 142944
rect 479536 142186 479564 200738
rect 485780 199436 485832 199442
rect 485780 199378 485832 199384
rect 483664 160200 483716 160206
rect 483664 160142 483716 160148
rect 483676 142934 483704 160142
rect 483664 142928 483716 142934
rect 483664 142870 483716 142876
rect 479524 142180 479576 142186
rect 479524 142122 479576 142128
rect 481916 142180 481968 142186
rect 481916 142122 481968 142128
rect 481928 140826 481956 142122
rect 462964 140820 463016 140826
rect 462964 140762 463016 140768
rect 481916 140820 481968 140826
rect 481916 140762 481968 140768
rect 462976 67561 463004 140762
rect 481928 139890 481956 140762
rect 485792 139890 485820 199378
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 489920 162172 489972 162178
rect 489920 162114 489972 162120
rect 489932 139890 489960 162114
rect 496820 161696 496872 161702
rect 496820 161638 496872 161644
rect 494060 161628 494112 161634
rect 494060 161570 494112 161576
rect 494072 139890 494100 161570
rect 496832 151814 496860 161638
rect 513380 161560 513432 161566
rect 513380 161502 513432 161508
rect 504364 160132 504416 160138
rect 504364 160074 504416 160080
rect 496832 151786 497688 151814
rect 497660 139890 497688 151786
rect 504376 143546 504404 160074
rect 513392 151814 513420 161502
rect 517520 161492 517572 161498
rect 517520 161434 517572 161440
rect 513392 151786 513512 151814
rect 504364 143540 504416 143546
rect 504364 143482 504416 143488
rect 505652 143540 505704 143546
rect 505652 143482 505704 143488
rect 501696 142996 501748 143002
rect 501696 142938 501748 142944
rect 501708 139890 501736 142938
rect 505664 139890 505692 143482
rect 509608 142860 509660 142866
rect 509608 142802 509660 142808
rect 509620 139890 509648 142802
rect 513484 139890 513512 151786
rect 517532 139890 517560 161434
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 533356 167006 533384 311102
rect 533344 167000 533396 167006
rect 533344 166942 533396 166948
rect 528560 163532 528612 163538
rect 528560 163474 528612 163480
rect 528572 151814 528600 163474
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 533988 142928 534040 142934
rect 533988 142870 534040 142876
rect 534000 142186 534028 142870
rect 533988 142180 534040 142186
rect 533988 142122 534040 142128
rect 534000 139890 534028 142122
rect 534736 140078 534764 319534
rect 538864 319524 538916 319530
rect 538864 319466 538916 319472
rect 537484 293276 537536 293282
rect 537484 293218 537536 293224
rect 536840 276752 536892 276758
rect 536840 276694 536892 276700
rect 536852 151814 536880 276694
rect 537496 193186 537524 293218
rect 537484 193180 537536 193186
rect 537484 193122 537536 193128
rect 536852 151786 537248 151814
rect 534724 140072 534776 140078
rect 534724 140014 534776 140020
rect 481928 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501708 139862 502044 139890
rect 505664 139862 506000 139890
rect 509620 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533692 139862 534028 139890
rect 537220 139890 537248 151786
rect 537220 139862 537648 139890
rect 538876 138582 538904 319466
rect 543740 319456 543792 319462
rect 543740 319398 543792 319404
rect 540980 318164 541032 318170
rect 540980 318106 541032 318112
rect 539692 315512 539744 315518
rect 539692 315454 539744 315460
rect 539600 315444 539652 315450
rect 539600 315386 539652 315392
rect 538956 314084 539008 314090
rect 538956 314026 539008 314032
rect 538864 138576 538916 138582
rect 538864 138518 538916 138524
rect 538968 138009 538996 314026
rect 539048 285048 539100 285054
rect 539048 284990 539100 284996
rect 539060 151814 539088 284990
rect 539060 151786 539364 151814
rect 538954 138000 539010 138009
rect 538954 137935 539010 137944
rect 539336 135697 539364 151786
rect 539322 135688 539378 135697
rect 539322 135623 539378 135632
rect 539612 97209 539640 315386
rect 539704 119649 539732 315454
rect 540336 311296 540388 311302
rect 540336 311238 540388 311244
rect 539784 283688 539836 283694
rect 539784 283630 539836 283636
rect 539690 119640 539746 119649
rect 539690 119575 539746 119584
rect 539796 99249 539824 283630
rect 540244 278044 540296 278050
rect 540244 277986 540296 277992
rect 539968 276820 540020 276826
rect 539968 276762 540020 276768
rect 539876 142180 539928 142186
rect 539876 142122 539928 142128
rect 539782 99240 539838 99249
rect 539782 99175 539838 99184
rect 539598 97200 539654 97209
rect 539598 97135 539654 97144
rect 462318 67552 462374 67561
rect 462318 67487 462374 67496
rect 462962 67552 463018 67561
rect 462962 67487 463018 67496
rect 461584 41404 461636 41410
rect 461584 41346 461636 41352
rect 462332 31754 462360 67487
rect 536840 41404 536892 41410
rect 536840 41346 536892 41352
rect 536852 41041 536880 41346
rect 536838 41032 536894 41041
rect 536838 40967 536894 40976
rect 539888 33697 539916 142122
rect 539980 112849 540008 276762
rect 540152 272536 540204 272542
rect 540152 272478 540204 272484
rect 540060 271244 540112 271250
rect 540060 271186 540112 271192
rect 539966 112840 540022 112849
rect 539966 112775 540022 112784
rect 540072 111489 540100 271186
rect 540164 117065 540192 272478
rect 540256 125225 540284 277986
rect 540348 129305 540376 311238
rect 540334 129296 540390 129305
rect 540334 129231 540390 129240
rect 540242 125216 540298 125225
rect 540242 125151 540298 125160
rect 540150 117056 540206 117065
rect 540150 116991 540206 117000
rect 540058 111480 540114 111489
rect 540058 111415 540114 111424
rect 540992 82385 541020 318106
rect 543280 318096 543332 318102
rect 543280 318038 543332 318044
rect 542636 317008 542688 317014
rect 542636 316950 542688 316956
rect 541072 316940 541124 316946
rect 541072 316882 541124 316888
rect 541084 108905 541112 316882
rect 542452 316872 542504 316878
rect 542452 316814 542504 316820
rect 541164 291712 541216 291718
rect 541164 291654 541216 291660
rect 541176 115025 541204 291654
rect 541532 279472 541584 279478
rect 541532 279414 541584 279420
rect 541440 275324 541492 275330
rect 541440 275266 541492 275272
rect 541256 273964 541308 273970
rect 541256 273906 541308 273912
rect 541162 115016 541218 115025
rect 541162 114951 541218 114960
rect 541070 108896 541126 108905
rect 541070 108831 541126 108840
rect 541268 104825 541296 273906
rect 541348 271176 541400 271182
rect 541348 271118 541400 271124
rect 541254 104816 541310 104825
rect 541254 104751 541310 104760
rect 541360 102785 541388 271118
rect 541452 106865 541480 275266
rect 541544 133385 541572 279414
rect 541530 133376 541586 133385
rect 541530 133311 541586 133320
rect 541438 106856 541494 106865
rect 541438 106791 541494 106800
rect 541346 102776 541402 102785
rect 541346 102711 541402 102720
rect 542464 90545 542492 316814
rect 542544 314016 542596 314022
rect 542544 313958 542596 313964
rect 542556 92585 542584 313958
rect 542648 121145 542676 316950
rect 542728 269952 542780 269958
rect 542728 269894 542780 269900
rect 542634 121136 542690 121145
rect 542634 121071 542690 121080
rect 542542 92576 542598 92585
rect 542542 92511 542598 92520
rect 542450 90536 542506 90545
rect 542450 90471 542506 90480
rect 542740 86465 542768 269894
rect 542912 268592 542964 268598
rect 542912 268534 542964 268540
rect 542820 268524 542872 268530
rect 542820 268466 542872 268472
rect 542832 94625 542860 268466
rect 542924 127265 542952 268534
rect 543188 140072 543240 140078
rect 543188 140014 543240 140020
rect 543096 138576 543148 138582
rect 543096 138518 543148 138524
rect 543002 136776 543058 136785
rect 543002 136711 543058 136720
rect 542910 127256 542966 127265
rect 542910 127191 542966 127200
rect 543016 100745 543044 136711
rect 543108 123185 543136 138518
rect 543200 131345 543228 140014
rect 543186 131336 543242 131345
rect 543186 131271 543242 131280
rect 543094 123176 543150 123185
rect 543094 123111 543150 123120
rect 543002 100736 543058 100745
rect 543002 100671 543058 100680
rect 542818 94616 542874 94625
rect 542818 94551 542874 94560
rect 543292 88505 543320 318038
rect 543278 88496 543334 88505
rect 543278 88431 543334 88440
rect 542726 86456 542782 86465
rect 542726 86391 542782 86400
rect 540978 82376 541034 82385
rect 540978 82311 541034 82320
rect 543752 51134 543780 319398
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 547144 312588 547196 312594
rect 547144 312530 547196 312536
rect 544384 288992 544436 288998
rect 544384 288934 544436 288940
rect 544396 73166 544424 288934
rect 544384 73160 544436 73166
rect 544384 73102 544436 73108
rect 547156 60722 547184 312530
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 565084 309800 565136 309806
rect 565084 309742 565136 309748
rect 562324 303612 562376 303618
rect 562324 303554 562376 303560
rect 548524 301640 548576 301646
rect 548524 301582 548576 301588
rect 548536 153202 548564 301582
rect 554044 283620 554096 283626
rect 554044 283562 554096 283568
rect 548524 153196 548576 153202
rect 548524 153138 548576 153144
rect 554056 139398 554084 283562
rect 555424 282192 555476 282198
rect 555424 282134 555476 282140
rect 555436 179382 555464 282134
rect 559564 280832 559616 280838
rect 559564 280774 559616 280780
rect 559576 219434 559604 280774
rect 559564 219428 559616 219434
rect 559564 219370 559616 219376
rect 555424 179376 555476 179382
rect 555424 179318 555476 179324
rect 554044 139392 554096 139398
rect 554044 139334 554096 139340
rect 547144 60716 547196 60722
rect 547144 60658 547196 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 539874 33688 539930 33697
rect 539874 33623 539930 33632
rect 462320 31748 462372 31754
rect 462320 31690 462372 31696
rect 460204 29640 460256 29646
rect 460204 29582 460256 29588
rect 386144 28280 386196 28286
rect 386144 28222 386196 28228
rect 562336 20670 562364 303554
rect 563704 297968 563756 297974
rect 563704 297910 563756 297916
rect 562324 20664 562376 20670
rect 562324 20606 562376 20612
rect 563716 6866 563744 297910
rect 565096 33114 565124 309742
rect 569224 307080 569276 307086
rect 569224 307022 569276 307028
rect 566464 300008 566516 300014
rect 566464 299950 566516 299956
rect 566476 100706 566504 299950
rect 569236 113150 569264 307022
rect 574744 305788 574796 305794
rect 574744 305730 574796 305736
rect 573364 295996 573416 296002
rect 573364 295938 573416 295944
rect 571984 290488 572036 290494
rect 571984 290430 572036 290436
rect 570604 284980 570656 284986
rect 570604 284922 570656 284928
rect 570616 233238 570644 284922
rect 571996 245614 572024 290430
rect 571984 245608 572036 245614
rect 571984 245550 572036 245556
rect 570604 233232 570656 233238
rect 570604 233174 570656 233180
rect 569224 113144 569276 113150
rect 569224 113086 569276 113092
rect 566464 100700 566516 100706
rect 566464 100642 566516 100648
rect 573376 46918 573404 295938
rect 574756 206990 574784 305730
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 578884 294500 578936 294506
rect 578884 294442 578936 294448
rect 576124 287700 576176 287706
rect 576124 287642 576176 287648
rect 574744 206984 574796 206990
rect 574744 206926 574796 206932
rect 576136 126954 576164 287642
rect 576124 126948 576176 126954
rect 576124 126890 576176 126896
rect 578896 86193 578924 294442
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580264 269884 580316 269890
rect 580264 269826 580316 269832
rect 580276 258913 580304 269826
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 578882 86184 578938 86193
rect 578882 86119 578938 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 573364 46912 573416 46918
rect 573364 46854 573416 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 565084 33108 565136 33114
rect 580170 33079 580172 33088
rect 565084 33050 565136 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 563704 6860 563756 6866
rect 563704 6802 563756 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 385776 3596 385828 3602
rect 385776 3538 385828 3544
rect 385684 2236 385736 2242
rect 385684 2178 385736 2184
rect 383016 2168 383068 2174
rect 383016 2110 383068 2116
rect 381636 2100 381688 2106
rect 381636 2042 381688 2048
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 23478 687792 23534 687848
rect 170310 700304 170366 700360
rect 332506 700576 332562 700632
rect 300122 700440 300178 700496
rect 88338 685072 88394 685128
rect 3422 684256 3478 684312
rect 3146 658180 3148 658200
rect 3148 658180 3200 658200
rect 3200 658180 3202 658200
rect 3146 658144 3202 658180
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3698 632032 3754 632088
rect 3606 475632 3662 475688
rect 3514 462576 3570 462632
rect 3422 449520 3478 449576
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 361762 678988 361764 679008
rect 361764 678988 361816 679008
rect 361816 678988 361818 679008
rect 361762 678952 361818 678988
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361670 656920 361726 656976
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612856 361634 612912
rect 361762 601840 361818 601896
rect 361762 590824 361818 590880
rect 361762 579808 361818 579864
rect 361762 568792 361818 568848
rect 361578 557796 361634 557832
rect 361578 557776 361580 557796
rect 361580 557776 361632 557796
rect 361632 557776 361634 557796
rect 361578 546760 361634 546816
rect 361578 535764 361634 535800
rect 361578 535744 361580 535764
rect 361580 535744 361632 535764
rect 361632 535744 361634 535764
rect 361762 524728 361818 524784
rect 3790 501744 3846 501800
rect 3698 423544 3754 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 361762 491680 361818 491736
rect 361762 480664 361818 480720
rect 362222 469648 362278 469704
rect 361762 458632 361818 458688
rect 361762 436600 361818 436656
rect 361578 414568 361634 414624
rect 362314 447616 362370 447672
rect 362406 425584 362462 425640
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3882 397432 3938 397488
rect 3422 358400 3478 358456
rect 3514 345344 3570 345400
rect 3606 319232 3662 319288
rect 3422 293120 3478 293176
rect 3330 162832 3386 162888
rect 3238 149776 3294 149832
rect 3146 84632 3202 84688
rect 3146 71576 3202 71632
rect 3146 58520 3202 58576
rect 3514 267144 3570 267200
rect 3698 306176 3754 306232
rect 3606 254088 3662 254144
rect 361578 392536 361634 392592
rect 361578 381520 361634 381576
rect 3974 371320 4030 371376
rect 3790 241032 3846 241088
rect 3698 97552 3754 97608
rect 361578 370504 361634 370560
rect 362222 359488 362278 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 361762 315424 361818 315480
rect 363602 305768 363658 305824
rect 3882 214920 3938 214976
rect 3974 201864 4030 201920
rect 4066 188808 4122 188864
rect 20902 73616 20958 73672
rect 15198 48864 15254 48920
rect 18878 49544 18934 49600
rect 21454 73616 21510 73672
rect 20074 46688 20130 46744
rect 3422 45484 3478 45520
rect 3422 45464 3424 45484
rect 3424 45464 3476 45484
rect 3476 45464 3478 45484
rect 6918 44784 6974 44840
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 5262 3984 5318 4040
rect 6458 3576 6514 3632
rect 8758 3712 8814 3768
rect 13542 3848 13598 3904
rect 359646 46416 359702 46472
rect 359830 46552 359886 46608
rect 361762 304408 361818 304464
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361670 216316 361672 216336
rect 361672 216316 361724 216336
rect 361724 216316 361726 216336
rect 361670 216280 361726 216316
rect 361762 205264 361818 205320
rect 361762 194248 361818 194304
rect 361762 183232 361818 183288
rect 361762 172216 361818 172272
rect 361762 161200 361818 161256
rect 361762 139168 361818 139224
rect 361762 128152 361818 128208
rect 361762 117136 361818 117192
rect 361762 106120 361818 106176
rect 361762 95140 361764 95160
rect 361764 95140 361816 95160
rect 361816 95140 361818 95160
rect 361762 95104 361818 95140
rect 361670 84124 361672 84144
rect 361672 84124 361724 84144
rect 361724 84124 361726 84144
rect 361670 84088 361726 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51076 361764 51096
rect 361764 51076 361816 51096
rect 361816 51076 361818 51096
rect 361762 51040 361818 51076
rect 362406 297608 362462 297664
rect 362222 3984 362278 4040
rect 362590 271360 362646 271416
rect 362590 150184 362646 150240
rect 370502 306856 370558 306912
rect 365166 297472 365222 297528
rect 365350 297336 365406 297392
rect 371974 297744 372030 297800
rect 372158 294480 372214 294536
rect 373538 300056 373594 300112
rect 376022 306176 376078 306232
rect 379242 302776 379298 302832
rect 380346 306720 380402 306776
rect 372158 3848 372214 3904
rect 371974 3712 372030 3768
rect 370502 3576 370558 3632
rect 381818 306040 381874 306096
rect 381634 305904 381690 305960
rect 381450 302912 381506 302968
rect 382186 303048 382242 303104
rect 382186 44784 382242 44840
rect 383014 300192 383070 300248
rect 381818 3440 381874 3496
rect 384578 46688 384634 46744
rect 384762 289040 384818 289096
rect 384946 46960 385002 47016
rect 385958 46824 386014 46880
rect 420826 682760 420882 682816
rect 444194 422048 444250 422104
rect 444102 421912 444158 421968
rect 442814 387096 442870 387152
rect 420734 334464 420790 334520
rect 428094 334464 428150 334520
rect 421562 162696 421618 162752
rect 428646 162696 428702 162752
rect 432602 332832 432658 332888
rect 432142 314472 432198 314528
rect 432786 329160 432842 329216
rect 432694 325488 432750 325544
rect 432970 321816 433026 321872
rect 432878 318144 432934 318200
rect 432602 310800 432658 310856
rect 432234 307128 432290 307184
rect 442722 321544 442778 321600
rect 444378 421776 444434 421832
rect 445666 683304 445722 683360
rect 450358 683168 450414 683224
rect 448150 516704 448206 516760
rect 448058 514120 448114 514176
rect 448426 516160 448482 516216
rect 448334 512760 448390 512816
rect 448242 510448 448298 510504
rect 448058 507728 448114 507784
rect 447966 503648 448022 503704
rect 447138 383832 447194 383888
rect 447138 383152 447194 383208
rect 447230 382472 447286 382528
rect 447138 381792 447194 381848
rect 447230 381112 447286 381168
rect 447138 380432 447194 380488
rect 447230 379752 447286 379808
rect 447138 379072 447194 379128
rect 447230 378392 447286 378448
rect 447138 377712 447194 377768
rect 447230 377032 447286 377088
rect 447138 376352 447194 376408
rect 447230 375672 447286 375728
rect 447138 374992 447194 375048
rect 447230 374312 447286 374368
rect 447138 373632 447194 373688
rect 447230 372952 447286 373008
rect 447138 372272 447194 372328
rect 447230 371592 447286 371648
rect 447138 370912 447194 370968
rect 447230 370232 447286 370288
rect 447138 369552 447194 369608
rect 447230 368872 447286 368928
rect 447138 368192 447194 368248
rect 447230 367512 447286 367568
rect 447138 366832 447194 366888
rect 447230 366152 447286 366208
rect 447230 365472 447286 365528
rect 447138 364792 447194 364848
rect 447138 364112 447194 364168
rect 447230 363432 447286 363488
rect 447230 362752 447286 362808
rect 447138 362072 447194 362128
rect 447230 361392 447286 361448
rect 447138 360712 447194 360768
rect 447230 360032 447286 360088
rect 447138 359352 447194 359408
rect 447598 352552 447654 352608
rect 447138 351908 447140 351928
rect 447140 351908 447192 351928
rect 447192 351908 447194 351928
rect 447138 351872 447194 351908
rect 447414 351192 447470 351248
rect 447138 350548 447140 350568
rect 447140 350548 447192 350568
rect 447192 350548 447194 350568
rect 447138 350512 447194 350548
rect 447138 347112 447194 347168
rect 447322 343712 447378 343768
rect 447138 341672 447194 341728
rect 447230 341012 447286 341048
rect 447230 340992 447232 341012
rect 447232 340992 447284 341012
rect 447284 340992 447286 341012
rect 447138 340312 447194 340368
rect 447230 339632 447286 339688
rect 447230 338952 447286 339008
rect 447138 338272 447194 338328
rect 447230 337592 447286 337648
rect 447138 336912 447194 336968
rect 447230 336232 447286 336288
rect 447322 335552 447378 335608
rect 447322 334872 447378 334928
rect 447230 334192 447286 334248
rect 447322 333512 447378 333568
rect 447230 332832 447286 332888
rect 447230 331472 447286 331528
rect 447322 330792 447378 330848
rect 447230 330132 447286 330168
rect 447230 330112 447232 330132
rect 447232 330112 447284 330132
rect 447284 330112 447286 330132
rect 447230 329432 447286 329488
rect 447230 328752 447286 328808
rect 447230 328072 447286 328128
rect 447322 327392 447378 327448
rect 447230 326712 447286 326768
rect 447322 326032 447378 326088
rect 447782 348472 447838 348528
rect 447690 347792 447746 347848
rect 447598 344392 447654 344448
rect 447874 343032 447930 343088
rect 447506 332152 447562 332208
rect 448150 505144 448206 505200
rect 448426 510448 448482 510504
rect 449714 505620 449770 505676
rect 449806 501268 449862 501324
rect 448518 500268 448574 500304
rect 448518 500248 448520 500268
rect 448520 500248 448572 500268
rect 448572 500248 448574 500268
rect 448426 496068 448428 496088
rect 448428 496068 448480 496088
rect 448480 496068 448482 496088
rect 448426 496032 448482 496068
rect 449070 389816 449126 389872
rect 448978 386960 449034 387016
rect 449070 354592 449126 354648
rect 448978 353232 449034 353288
rect 448426 349152 448482 349208
rect 449254 385600 449310 385656
rect 449162 342352 449218 342408
rect 448242 326712 448298 326768
rect 448150 325352 448206 325408
rect 448426 325352 448482 325408
rect 447966 324672 448022 324728
rect 449438 356632 449494 356688
rect 449346 355272 449402 355328
rect 449622 357312 449678 357368
rect 449714 355952 449770 356008
rect 449530 353912 449586 353968
rect 449714 349832 449770 349888
rect 449622 343032 449678 343088
rect 449254 324128 449310 324184
rect 450266 358808 450322 358864
rect 450082 358400 450138 358456
rect 449898 346840 449954 346896
rect 449806 345752 449862 345808
rect 449806 345072 449862 345128
rect 450358 319912 450414 319968
rect 494794 700304 494850 700360
rect 527178 699760 527234 699816
rect 462318 669840 462374 669896
rect 458086 662496 458142 662552
rect 457718 659912 457774 659968
rect 457626 652840 457682 652896
rect 457534 645904 457590 645960
rect 457350 623872 457406 623928
rect 457258 611360 457314 611416
rect 457442 618296 457498 618352
rect 457994 657464 458050 657520
rect 457902 650120 457958 650176
rect 457810 621016 457866 621072
rect 459190 655696 459246 655752
rect 459098 647672 459154 647728
rect 459006 643184 459062 643240
rect 458914 640328 458970 640384
rect 458822 615984 458878 616040
rect 458730 608640 458786 608696
rect 459006 599664 459062 599720
rect 459098 599528 459154 599584
rect 458914 598168 458970 598224
rect 459282 637880 459338 637936
rect 459190 595448 459246 595504
rect 459374 635432 459430 635488
rect 459282 541592 459338 541648
rect 459466 633392 459522 633448
rect 459374 522280 459430 522336
rect 459742 628700 459798 628756
rect 459558 626252 459614 626308
rect 459650 601840 459706 601896
rect 459466 518064 459522 518120
rect 459834 614080 459890 614136
rect 459926 606328 459982 606384
rect 460202 603608 460258 603664
rect 462318 562944 462374 563000
rect 468666 523640 468722 523696
rect 494058 516704 494114 516760
rect 491850 516180 491906 516216
rect 491850 516160 491852 516180
rect 491852 516160 491904 516180
rect 491904 516160 491906 516180
rect 494058 515888 494114 515944
rect 494058 512488 494114 512544
rect 494426 516704 494482 516760
rect 494334 508816 494390 508872
rect 494242 505688 494298 505744
rect 495070 505724 495072 505744
rect 495072 505724 495124 505744
rect 495124 505724 495126 505744
rect 495070 505688 495126 505724
rect 494058 501200 494114 501256
rect 481822 496848 481878 496904
rect 483846 496848 483902 496904
rect 487986 453872 488042 453928
rect 471978 410488 472034 410544
rect 472898 389000 472954 389056
rect 474370 389000 474426 389056
rect 475106 389000 475162 389056
rect 477314 389000 477370 389056
rect 479522 389000 479578 389056
rect 473634 388864 473690 388920
rect 475842 388864 475898 388920
rect 509606 372408 509662 372464
rect 509330 366968 509386 367024
rect 450726 322904 450782 322960
rect 507306 322632 507362 322688
rect 507122 322496 507178 322552
rect 451554 158208 451610 158264
rect 451738 156848 451794 156904
rect 451738 154128 451794 154184
rect 451646 152768 451702 152824
rect 451462 151444 451464 151464
rect 451464 151444 451516 151464
rect 451516 151444 451518 151464
rect 451462 151408 451518 151444
rect 451554 139168 451610 139224
rect 452014 128288 452070 128344
rect 452198 148688 452254 148744
rect 452198 132404 452200 132424
rect 452200 132404 452252 132424
rect 452252 132404 452254 132424
rect 452198 132368 452254 132404
rect 452566 155524 452568 155544
rect 452568 155524 452620 155544
rect 452620 155524 452622 155544
rect 452566 155488 452622 155524
rect 452382 150048 452438 150104
rect 452566 147328 452622 147384
rect 452566 146004 452568 146024
rect 452568 146004 452620 146024
rect 452620 146004 452622 146024
rect 452566 145968 452622 146004
rect 452566 144644 452568 144664
rect 452568 144644 452620 144664
rect 452620 144644 452622 144664
rect 452566 144608 452622 144644
rect 452566 143284 452568 143304
rect 452568 143284 452620 143304
rect 452620 143284 452622 143304
rect 452566 143248 452622 143284
rect 452566 141924 452568 141944
rect 452568 141924 452620 141944
rect 452620 141924 452622 141944
rect 452566 141888 452622 141924
rect 452566 140528 452622 140584
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452566 136484 452568 136504
rect 452568 136484 452620 136504
rect 452620 136484 452622 136504
rect 452566 136448 452622 136484
rect 452566 135124 452568 135144
rect 452568 135124 452620 135144
rect 452620 135124 452622 135144
rect 452566 135088 452622 135124
rect 452566 133764 452568 133784
rect 452568 133764 452620 133784
rect 452620 133764 452622 133784
rect 452566 133728 452622 133764
rect 452382 131044 452384 131064
rect 452384 131044 452436 131064
rect 452436 131044 452438 131064
rect 452382 131008 452438 131044
rect 452290 129648 452346 129704
rect 452382 126948 452438 126984
rect 452382 126928 452384 126948
rect 452384 126928 452436 126948
rect 452436 126928 452438 126948
rect 452106 125568 452162 125624
rect 451922 124208 451978 124264
rect 451922 122848 451978 122904
rect 451922 121488 451978 121544
rect 458638 321408 458694 321464
rect 459742 321136 459798 321192
rect 460294 321816 460350 321872
rect 460570 321000 460626 321056
rect 456798 262656 456854 262712
rect 456798 248784 456854 248840
rect 456798 207168 456854 207224
rect 457810 234912 457866 234968
rect 458086 234912 458142 234968
rect 459466 221040 459522 221096
rect 471058 320048 471114 320104
rect 471610 319912 471666 319968
rect 471334 319776 471390 319832
rect 480442 321272 480498 321328
rect 479614 320048 479670 320104
rect 481546 321680 481602 321736
rect 481822 321544 481878 321600
rect 484490 306176 484546 306232
rect 494978 313928 495034 313984
rect 497278 319368 497334 319424
rect 507674 320728 507730 320784
rect 509422 358808 509478 358864
rect 509514 349424 509570 349480
rect 509790 333104 509846 333160
rect 509698 326032 509754 326088
rect 510710 368872 510766 368928
rect 510618 366696 510674 366752
rect 510066 332968 510122 333024
rect 510158 329160 510214 329216
rect 510250 328072 510306 328128
rect 510158 322904 510214 322960
rect 509698 303048 509754 303104
rect 510250 300056 510306 300112
rect 510802 360712 510858 360768
rect 510894 355816 510950 355872
rect 510986 352552 511042 352608
rect 511170 342760 511226 342816
rect 512090 380296 512146 380352
rect 511998 378120 512054 378176
rect 512182 378664 512238 378720
rect 512090 377576 512146 377632
rect 512182 376488 512238 376544
rect 511998 371048 512054 371104
rect 512090 370504 512146 370560
rect 512090 364540 512146 364576
rect 512090 364520 512092 364540
rect 512092 364520 512144 364540
rect 512144 364520 512146 364540
rect 511998 363976 512054 364032
rect 511998 362344 512054 362400
rect 511998 358536 512054 358592
rect 511538 343304 511594 343360
rect 511170 302912 511226 302968
rect 512090 357992 512146 358048
rect 512090 357468 512146 357504
rect 512090 357448 512092 357468
rect 512092 357448 512144 357468
rect 512144 357448 512146 357468
rect 512090 356380 512146 356416
rect 512090 356360 512092 356380
rect 512092 356360 512144 356380
rect 512144 356360 512146 356380
rect 512090 354184 512146 354240
rect 512090 350920 512146 350976
rect 512090 349288 512146 349344
rect 512090 346024 512146 346080
rect 512090 345480 512146 345536
rect 512734 384648 512790 384704
rect 513286 384104 513342 384160
rect 512918 383560 512974 383616
rect 513286 383016 513342 383072
rect 513194 382492 513250 382528
rect 513194 382472 513196 382492
rect 513196 382472 513248 382492
rect 513248 382472 513250 382492
rect 512366 381928 512422 381984
rect 513286 381384 513342 381440
rect 512366 380840 512422 380896
rect 512274 375944 512330 376000
rect 512826 379752 512882 379808
rect 513286 379208 513342 379264
rect 513194 377032 513250 377088
rect 513286 375400 513342 375456
rect 512458 374856 512514 374912
rect 512734 374312 512790 374368
rect 512826 373768 512882 373824
rect 513286 373224 513342 373280
rect 512550 372136 512606 372192
rect 512274 371592 512330 371648
rect 513286 369996 513288 370016
rect 513288 369996 513340 370016
rect 513340 369996 513342 370016
rect 513286 369960 513342 369996
rect 513010 369416 513066 369472
rect 512366 368328 512422 368384
rect 512642 367784 512698 367840
rect 512458 366152 512514 366208
rect 512458 365064 512514 365120
rect 513286 363432 513342 363488
rect 513286 362888 513342 362944
rect 513102 361820 513158 361856
rect 513102 361800 513104 361820
rect 513104 361800 513156 361820
rect 513156 361800 513158 361820
rect 513286 361256 513342 361312
rect 512550 360168 512606 360224
rect 513286 359624 513342 359680
rect 512734 356904 512790 356960
rect 513194 355272 513250 355328
rect 513286 354764 513288 354784
rect 513288 354764 513340 354784
rect 513340 354764 513342 354784
rect 513286 354728 513342 354764
rect 513286 353640 513342 353696
rect 512918 353096 512974 353152
rect 513286 352008 513342 352064
rect 512826 351484 512882 351520
rect 512826 351464 512828 351484
rect 512828 351464 512880 351484
rect 512880 351464 512882 351484
rect 513010 350376 513066 350432
rect 512826 348744 512882 348800
rect 512918 348200 512974 348256
rect 512642 347656 512698 347712
rect 513286 347112 513342 347168
rect 512826 346588 512882 346624
rect 512826 346568 512828 346588
rect 512828 346568 512880 346588
rect 512880 346568 512882 346588
rect 513286 344936 513342 344992
rect 512642 344392 512698 344448
rect 512826 343868 512882 343904
rect 512826 343848 512828 343868
rect 512828 343848 512880 343868
rect 512880 343848 512882 343868
rect 512642 342216 512698 342272
rect 513286 341672 513342 341728
rect 513010 341128 513066 341184
rect 513194 340584 513250 340640
rect 513010 339532 513012 339552
rect 513012 339532 513064 339552
rect 513064 339532 513066 339552
rect 513010 339496 513066 339532
rect 513286 340040 513342 340096
rect 513194 338952 513250 339008
rect 513286 338408 513342 338464
rect 513194 337864 513250 337920
rect 513194 337320 513250 337376
rect 513286 336812 513288 336832
rect 513288 336812 513340 336832
rect 513340 336812 513342 336832
rect 513286 336776 513342 336812
rect 513194 336232 513250 336288
rect 513286 335688 513342 335744
rect 513194 335144 513250 335200
rect 513286 334056 513342 334112
rect 513286 331880 513342 331936
rect 512734 330792 512790 330848
rect 512734 325352 512790 325408
rect 512642 305768 512698 305824
rect 513562 365608 513618 365664
rect 515494 302776 515550 302832
rect 518346 300192 518402 300248
rect 559654 699760 559710 699816
rect 580170 697176 580226 697232
rect 557538 442856 557594 442912
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 578882 644000 578938 644056
rect 579986 630808 580042 630864
rect 579618 590960 579674 591016
rect 579618 577632 579674 577688
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579618 471416 579674 471472
rect 579618 431568 579674 431624
rect 579710 418240 579766 418296
rect 579618 378392 579674 378448
rect 580170 365064 580226 365120
rect 580170 325216 580226 325272
rect 580354 617480 580410 617536
rect 580446 564304 580502 564360
rect 580538 458088 580594 458144
rect 580630 404912 580686 404968
rect 580722 351872 580778 351928
rect 529294 261568 529350 261624
rect 530122 243616 530178 243672
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 538954 137944 539010 138000
rect 539322 135632 539378 135688
rect 539690 119584 539746 119640
rect 539782 99184 539838 99240
rect 539598 97144 539654 97200
rect 462318 67496 462374 67552
rect 462962 67496 463018 67552
rect 536838 40976 536894 41032
rect 539966 112784 540022 112840
rect 540334 129240 540390 129296
rect 540242 125160 540298 125216
rect 540150 117000 540206 117056
rect 540058 111424 540114 111480
rect 541162 114960 541218 115016
rect 541070 108840 541126 108896
rect 541254 104760 541310 104816
rect 541530 133320 541586 133376
rect 541438 106800 541494 106856
rect 541346 102720 541402 102776
rect 542634 121080 542690 121136
rect 542542 92520 542598 92576
rect 542450 90480 542506 90536
rect 543002 136720 543058 136776
rect 542910 127200 542966 127256
rect 543186 131280 543242 131336
rect 543094 123120 543150 123176
rect 543002 100680 543058 100736
rect 542818 94560 542874 94616
rect 543278 88440 543334 88496
rect 542726 86400 542782 86456
rect 540978 82320 541034 82376
rect 580170 312024 580226 312080
rect 540610 48864 540666 48920
rect 539874 33632 539930 33688
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 578882 86128 578938 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 332501 700634 332567 700637
rect 449566 700634 449572 700636
rect 332501 700632 449572 700634
rect 332501 700576 332506 700632
rect 332562 700576 449572 700632
rect 332501 700574 449572 700576
rect 332501 700571 332567 700574
rect 449566 700572 449572 700574
rect 449636 700572 449642 700636
rect 300117 700498 300183 700501
rect 444230 700498 444236 700500
rect 300117 700496 444236 700498
rect 300117 700440 300122 700496
rect 300178 700440 444236 700496
rect 300117 700438 444236 700440
rect 300117 700435 300183 700438
rect 444230 700436 444236 700438
rect 444300 700436 444306 700500
rect 170305 700362 170371 700365
rect 446254 700362 446260 700364
rect 170305 700360 446260 700362
rect 170305 700304 170310 700360
rect 170366 700304 446260 700360
rect 170305 700302 446260 700304
rect 170305 700299 170371 700302
rect 446254 700300 446260 700302
rect 446324 700300 446330 700364
rect 455086 700300 455092 700364
rect 455156 700362 455162 700364
rect 494789 700362 494855 700365
rect 455156 700360 494855 700362
rect 455156 700304 494794 700360
rect 494850 700304 494855 700360
rect 455156 700302 494855 700304
rect 455156 700300 455162 700302
rect 494789 700299 494855 700302
rect 527173 699818 527239 699821
rect 529974 699818 529980 699820
rect 527173 699816 529980 699818
rect 527173 699760 527178 699816
rect 527234 699760 529980 699816
rect 527173 699758 529980 699760
rect 527173 699755 527239 699758
rect 529974 699756 529980 699758
rect 530044 699756 530050 699820
rect 559414 699756 559420 699820
rect 559484 699818 559490 699820
rect 559649 699818 559715 699821
rect 559484 699816 559715 699818
rect 559484 699760 559654 699816
rect 559710 699760 559715 699816
rect 559484 699758 559715 699760
rect 559484 699756 559490 699758
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 23473 687850 23539 687853
rect 450486 687850 450492 687852
rect 23473 687848 450492 687850
rect 23473 687792 23478 687848
rect 23534 687792 450492 687848
rect 23473 687790 450492 687792
rect 23473 687787 23539 687790
rect 450486 687788 450492 687790
rect 450556 687788 450562 687852
rect 88333 685130 88399 685133
rect 446438 685130 446444 685132
rect 88333 685128 446444 685130
rect 88333 685072 88338 685128
rect 88394 685072 446444 685128
rect 88333 685070 446444 685072
rect 88333 685067 88399 685070
rect 446438 685068 446444 685070
rect 446508 685068 446514 685132
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect 3550 683300 3556 683364
rect 3620 683362 3626 683364
rect 445661 683362 445727 683365
rect 3620 683360 445727 683362
rect 3620 683304 445666 683360
rect 445722 683304 445727 683360
rect 3620 683302 445727 683304
rect 3620 683300 3626 683302
rect 445661 683299 445727 683302
rect 3734 683164 3740 683228
rect 3804 683226 3810 683228
rect 450353 683226 450419 683229
rect 3804 683224 450419 683226
rect 3804 683168 450358 683224
rect 450414 683168 450419 683224
rect 3804 683166 450419 683168
rect 3804 683164 3810 683166
rect 450353 683163 450419 683166
rect 3366 682756 3372 682820
rect 3436 682818 3442 682820
rect 420821 682818 420887 682821
rect 3436 682816 420887 682818
rect 3436 682760 420826 682816
rect 420882 682760 420887 682816
rect 3436 682758 420887 682760
rect 3436 682756 3442 682758
rect 420821 682755 420887 682758
rect 361757 679010 361823 679013
rect 359812 679008 361823 679010
rect 359812 678952 361762 679008
rect 361818 678952 361823 679008
rect 359812 678950 361823 678952
rect 361757 678947 361823 678950
rect -960 671258 480 671348
rect 3734 671258 3740 671260
rect -960 671198 3740 671258
rect -960 671108 480 671198
rect 3734 671196 3740 671198
rect 3804 671196 3810 671260
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 453246 669836 453252 669900
rect 453316 669898 453322 669900
rect 462313 669898 462379 669901
rect 453316 669896 462379 669898
rect 453316 669840 462318 669896
rect 462374 669840 462379 669896
rect 453316 669838 462379 669840
rect 453316 669836 453322 669838
rect 462313 669835 462379 669838
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 459502 667932 459508 667996
rect 459572 667994 459578 667996
rect 459572 667934 460092 667994
rect 459572 667932 459578 667934
rect 458030 665212 458036 665276
rect 458100 665274 458106 665276
rect 460062 665274 460122 665448
rect 458100 665214 460122 665274
rect 458100 665212 458106 665214
rect 458081 662554 458147 662557
rect 460062 662554 460122 663000
rect 458081 662552 460122 662554
rect 458081 662496 458086 662552
rect 458142 662496 460122 662552
rect 458081 662494 460122 662496
rect 458081 662491 458147 662494
rect 457713 659970 457779 659973
rect 460062 659970 460122 660552
rect 457713 659968 460122 659970
rect 457713 659912 457718 659968
rect 457774 659912 460122 659968
rect 457713 659910 460122 659912
rect 457713 659907 457779 659910
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 457989 657522 458055 657525
rect 460062 657522 460122 658104
rect 457989 657520 460122 657522
rect 457989 657464 457994 657520
rect 458050 657464 460122 657520
rect 457989 657462 460122 657464
rect 457989 657459 458055 657462
rect 583520 657236 584960 657476
rect 361665 656978 361731 656981
rect 359812 656976 361731 656978
rect 359812 656920 361670 656976
rect 361726 656920 361731 656976
rect 359812 656918 361731 656920
rect 361665 656915 361731 656918
rect 459185 655754 459251 655757
rect 459185 655752 460092 655754
rect 459185 655696 459190 655752
rect 459246 655696 460092 655752
rect 459185 655694 460092 655696
rect 459185 655691 459251 655694
rect 457621 652898 457687 652901
rect 460062 652898 460122 653208
rect 457621 652896 460122 652898
rect 457621 652840 457626 652896
rect 457682 652840 460122 652896
rect 457621 652838 460122 652840
rect 457621 652835 457687 652838
rect 457897 650178 457963 650181
rect 460062 650178 460122 650760
rect 457897 650176 460122 650178
rect 457897 650120 457902 650176
rect 457958 650120 460122 650176
rect 457897 650118 460122 650120
rect 457897 650115 457963 650118
rect 459093 647730 459159 647733
rect 460062 647730 460122 648312
rect 459093 647728 460122 647730
rect 459093 647672 459098 647728
rect 459154 647672 460122 647728
rect 459093 647670 460122 647672
rect 459093 647667 459159 647670
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 457529 645962 457595 645965
rect 457529 645960 460092 645962
rect 457529 645904 457534 645960
rect 457590 645904 460092 645960
rect 457529 645902 460092 645904
rect 457529 645899 457595 645902
rect -960 644996 480 645236
rect 578877 644058 578943 644061
rect 583520 644058 584960 644148
rect 578877 644056 584960 644058
rect 578877 644000 578882 644056
rect 578938 644000 584960 644056
rect 578877 643998 584960 644000
rect 578877 643995 578943 643998
rect 583520 643908 584960 643998
rect 459001 643242 459067 643245
rect 460062 643242 460122 643416
rect 459001 643240 460122 643242
rect 459001 643184 459006 643240
rect 459062 643184 460122 643240
rect 459001 643182 460122 643184
rect 459001 643179 459067 643182
rect 458909 640386 458975 640389
rect 460062 640386 460122 640968
rect 458909 640384 460122 640386
rect 458909 640328 458914 640384
rect 458970 640328 460122 640384
rect 458909 640326 460122 640328
rect 458909 640323 458975 640326
rect 459277 637938 459343 637941
rect 460062 637938 460122 638520
rect 459277 637936 460122 637938
rect 459277 637880 459282 637936
rect 459338 637880 460122 637936
rect 459277 637878 460122 637880
rect 459277 637875 459343 637878
rect 459369 635490 459435 635493
rect 460062 635490 460122 636072
rect 459369 635488 460122 635490
rect 459369 635432 459374 635488
rect 459430 635432 460122 635488
rect 459369 635430 460122 635432
rect 459369 635427 459435 635430
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459461 633450 459527 633453
rect 460062 633450 460122 633624
rect 459461 633448 460122 633450
rect 459461 633392 459466 633448
rect 459522 633392 460122 633448
rect 459461 633390 460122 633392
rect 459461 633387 459527 633390
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 459134 630668 459140 630732
rect 459204 630730 459210 630732
rect 460062 630730 460122 631176
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 459204 630670 460122 630730
rect 583520 630716 584960 630806
rect 459204 630668 459210 630670
rect 459737 628758 459803 628761
rect 459737 628756 460092 628758
rect 459737 628700 459742 628756
rect 459798 628700 460092 628756
rect 459737 628698 460092 628700
rect 459737 628695 459803 628698
rect 459553 626310 459619 626313
rect 459553 626308 460092 626310
rect 459553 626252 459558 626308
rect 459614 626252 460092 626308
rect 459553 626250 460092 626252
rect 459553 626247 459619 626250
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 457345 623930 457411 623933
rect 457345 623928 460092 623930
rect 457345 623872 457350 623928
rect 457406 623872 460092 623928
rect 457345 623870 460092 623872
rect 457345 623867 457411 623870
rect 457805 621074 457871 621077
rect 460062 621074 460122 621384
rect 457805 621072 460122 621074
rect 457805 621016 457810 621072
rect 457866 621016 460122 621072
rect 457805 621014 460122 621016
rect 457805 621011 457871 621014
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 457437 618354 457503 618357
rect 460062 618354 460122 618936
rect 457437 618352 460122 618354
rect 457437 618296 457442 618352
rect 457498 618296 460122 618352
rect 457437 618294 460122 618296
rect 457437 618291 457503 618294
rect 580349 617538 580415 617541
rect 583520 617538 584960 617628
rect 580349 617536 584960 617538
rect 580349 617480 580354 617536
rect 580410 617480 584960 617536
rect 580349 617478 584960 617480
rect 580349 617475 580415 617478
rect 583520 617388 584960 617478
rect 458817 616042 458883 616045
rect 460062 616042 460122 616488
rect 458817 616040 460122 616042
rect 458817 615984 458822 616040
rect 458878 615984 460122 616040
rect 458817 615982 460122 615984
rect 458817 615979 458883 615982
rect 459829 614138 459895 614141
rect 459829 614136 460092 614138
rect 459829 614080 459834 614136
rect 459890 614080 460092 614136
rect 459829 614078 460092 614080
rect 459829 614075 459895 614078
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 457253 611418 457319 611421
rect 460062 611418 460122 611592
rect 457253 611416 460122 611418
rect 457253 611360 457258 611416
rect 457314 611360 460122 611416
rect 457253 611358 460122 611360
rect 457253 611355 457319 611358
rect 458725 608698 458791 608701
rect 460062 608698 460122 609144
rect 458725 608696 460122 608698
rect 458725 608640 458730 608696
rect 458786 608640 460122 608696
rect 458725 608638 460122 608640
rect 458725 608635 458791 608638
rect 459921 606386 459987 606389
rect 460062 606386 460122 606696
rect 459921 606384 460122 606386
rect 459921 606328 459926 606384
rect 459982 606328 460122 606384
rect 459921 606326 460122 606328
rect 459921 606323 459987 606326
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 460062 603666 460122 604248
rect 583520 604060 584960 604300
rect 460197 603666 460263 603669
rect 460062 603664 460263 603666
rect 460062 603608 460202 603664
rect 460258 603608 460263 603664
rect 460062 603606 460263 603608
rect 460197 603603 460263 603606
rect 361757 601898 361823 601901
rect 359812 601896 361823 601898
rect 359812 601840 361762 601896
rect 361818 601840 361823 601896
rect 359812 601838 361823 601840
rect 361757 601835 361823 601838
rect 459645 601898 459711 601901
rect 459645 601896 460092 601898
rect 459645 601840 459650 601896
rect 459706 601840 460092 601896
rect 459645 601838 460092 601840
rect 459645 601835 459711 601838
rect 459001 599722 459067 599725
rect 474774 599722 474780 599724
rect 459001 599720 474780 599722
rect 459001 599664 459006 599720
rect 459062 599664 474780 599720
rect 459001 599662 474780 599664
rect 459001 599659 459067 599662
rect 474774 599660 474780 599662
rect 474844 599660 474850 599724
rect 459093 599586 459159 599589
rect 476430 599586 476436 599588
rect 459093 599584 476436 599586
rect 459093 599528 459098 599584
rect 459154 599528 476436 599584
rect 459093 599526 476436 599528
rect 459093 599523 459159 599526
rect 476430 599524 476436 599526
rect 476500 599524 476506 599588
rect 458909 598226 458975 598229
rect 474958 598226 474964 598228
rect 458909 598224 474964 598226
rect 458909 598168 458914 598224
rect 458970 598168 474964 598224
rect 458909 598166 474964 598168
rect 458909 598163 458975 598166
rect 474958 598164 474964 598166
rect 475028 598164 475034 598228
rect 459185 595506 459251 595509
rect 478822 595506 478828 595508
rect 459185 595504 478828 595506
rect 459185 595448 459190 595504
rect 459246 595448 478828 595504
rect 459185 595446 478828 595448
rect 459185 595443 459251 595446
rect 478822 595444 478828 595446
rect 478892 595444 478898 595508
rect -960 592908 480 593148
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 361757 590882 361823 590885
rect 359812 590880 361823 590882
rect 359812 590824 361762 590880
rect 361818 590824 361823 590880
rect 583520 590868 584960 590958
rect 359812 590822 361823 590824
rect 361757 590819 361823 590822
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect 361757 568850 361823 568853
rect 359812 568848 361823 568850
rect 359812 568792 361762 568848
rect 361818 568792 361823 568848
rect 359812 568790 361823 568792
rect 361757 568787 361823 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580441 564362 580507 564365
rect 583520 564362 584960 564452
rect 580441 564360 584960 564362
rect 580441 564304 580446 564360
rect 580502 564304 584960 564360
rect 580441 564302 584960 564304
rect 580441 564299 580507 564302
rect 583520 564212 584960 564302
rect 459502 562940 459508 563004
rect 459572 563002 459578 563004
rect 462313 563002 462379 563005
rect 459572 563000 462379 563002
rect 459572 562944 462318 563000
rect 462374 562944 462379 563000
rect 459572 562942 462379 562944
rect 459572 562940 459578 562942
rect 462313 562939 462379 562942
rect 361573 557834 361639 557837
rect 359812 557832 361639 557834
rect 359812 557776 361578 557832
rect 361634 557776 361639 557832
rect 359812 557774 361639 557776
rect 361573 557771 361639 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361573 546818 361639 546821
rect 359812 546816 361639 546818
rect 359812 546760 361578 546816
rect 361634 546760 361639 546816
rect 359812 546758 361639 546760
rect 361573 546755 361639 546758
rect 459277 541650 459343 541653
rect 474406 541650 474412 541652
rect 459277 541648 474412 541650
rect 459277 541592 459282 541648
rect 459338 541592 474412 541648
rect 459277 541590 474412 541592
rect 459277 541587 459343 541590
rect 474406 541588 474412 541590
rect 474476 541588 474482 541652
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 361573 535802 361639 535805
rect 359812 535800 361639 535802
rect 359812 535744 361578 535800
rect 361634 535744 361639 535800
rect 359812 535742 361639 535744
rect 361573 535739 361639 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361757 524786 361823 524789
rect 359812 524784 361823 524786
rect 359812 524728 361762 524784
rect 361818 524728 361823 524784
rect 359812 524726 361823 524728
rect 361757 524723 361823 524726
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 458030 523636 458036 523700
rect 458100 523698 458106 523700
rect 468661 523698 468727 523701
rect 458100 523696 468727 523698
rect 458100 523640 468666 523696
rect 468722 523640 468727 523696
rect 458100 523638 468727 523640
rect 458100 523636 458106 523638
rect 468661 523635 468727 523638
rect 459369 522338 459435 522341
rect 474590 522338 474596 522340
rect 459369 522336 474596 522338
rect 459369 522280 459374 522336
rect 459430 522280 474596 522336
rect 459369 522278 474596 522280
rect 459369 522275 459435 522278
rect 474590 522276 474596 522278
rect 474660 522276 474666 522340
rect 459461 518122 459527 518125
rect 472014 518122 472020 518124
rect 459461 518120 472020 518122
rect 459461 518064 459466 518120
rect 459522 518064 472020 518120
rect 459461 518062 472020 518064
rect 459461 518059 459527 518062
rect 472014 518060 472020 518062
rect 472084 518060 472090 518124
rect 448145 516762 448211 516765
rect 494053 516762 494119 516765
rect 494421 516762 494487 516765
rect 448145 516760 494487 516762
rect 448145 516704 448150 516760
rect 448206 516704 494058 516760
rect 494114 516704 494426 516760
rect 494482 516704 494487 516760
rect 448145 516702 494487 516704
rect 448145 516699 448211 516702
rect 494053 516699 494119 516702
rect 494421 516699 494487 516702
rect 448278 516156 448284 516220
rect 448348 516218 448354 516220
rect 448421 516218 448487 516221
rect 450126 516218 450186 516528
rect 448348 516216 450186 516218
rect 448348 516160 448426 516216
rect 448482 516160 450186 516216
rect 448348 516158 450186 516160
rect 491845 516218 491911 516221
rect 491845 516216 491954 516218
rect 491845 516160 491850 516216
rect 491906 516160 491954 516216
rect 448348 516156 448354 516158
rect 448421 516155 448487 516158
rect 491845 516155 491954 516160
rect 491894 515946 491954 516155
rect 494053 515946 494119 515949
rect 491894 515944 494119 515946
rect 491894 515888 494058 515944
rect 494114 515888 494119 515944
rect 491894 515886 494119 515888
rect 494053 515883 494119 515886
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 448053 514180 448119 514181
rect 448053 514178 448100 514180
rect 447972 514176 448100 514178
rect 448164 514178 448170 514180
rect 450126 514178 450186 514352
rect 447972 514120 448058 514176
rect 447972 514118 448100 514120
rect 448053 514116 448100 514118
rect 448164 514118 450186 514178
rect 448164 514116 448170 514118
rect 448053 514115 448119 514116
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 448329 512818 448395 512821
rect 448329 512816 450186 512818
rect 448329 512760 448334 512816
rect 448390 512760 450186 512816
rect 448329 512758 450186 512760
rect 448329 512755 448395 512758
rect 450126 512176 450186 512758
rect 494053 512546 494119 512549
rect 491894 512544 494119 512546
rect 491894 512488 494058 512544
rect 494114 512488 494119 512544
rect 491894 512486 494119 512488
rect 491894 512448 491954 512486
rect 494053 512483 494119 512486
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 448237 510506 448303 510509
rect 448421 510506 448487 510509
rect 448237 510504 450186 510506
rect 448237 510448 448242 510504
rect 448298 510448 448426 510504
rect 448482 510448 450186 510504
rect 448237 510446 450186 510448
rect 448237 510443 448303 510446
rect 448421 510443 448487 510446
rect 450126 510000 450186 510446
rect 491894 508874 491954 508912
rect 494329 508874 494395 508877
rect 491894 508872 494395 508874
rect 491894 508816 494334 508872
rect 494390 508816 494395 508872
rect 491894 508814 494395 508816
rect 494329 508811 494395 508814
rect 448053 507786 448119 507789
rect 450126 507786 450186 507824
rect 448053 507784 450186 507786
rect 448053 507728 448058 507784
rect 448114 507728 450186 507784
rect 448053 507726 450186 507728
rect 448053 507723 448119 507726
rect 494237 505746 494303 505749
rect 495065 505746 495131 505749
rect 491894 505744 495131 505746
rect 491894 505688 494242 505744
rect 494298 505688 495070 505744
rect 495126 505688 495131 505744
rect 491894 505686 495131 505688
rect 449709 505678 449775 505681
rect 449709 505676 450156 505678
rect 449709 505620 449714 505676
rect 449770 505648 450156 505676
rect 449770 505620 450186 505648
rect 449709 505618 450186 505620
rect 449709 505615 449775 505618
rect 448145 505202 448211 505205
rect 450126 505202 450186 505618
rect 491894 505376 491954 505686
rect 494237 505683 494303 505686
rect 495065 505683 495131 505686
rect 448145 505200 450186 505202
rect 448145 505144 448150 505200
rect 448206 505144 450186 505200
rect 448145 505142 450186 505144
rect 448145 505139 448211 505142
rect 447961 503706 448027 503709
rect 447961 503704 450186 503706
rect 447961 503648 447966 503704
rect 448022 503648 450186 503704
rect 447961 503646 450186 503648
rect 447961 503643 448027 503646
rect 450126 503472 450186 503646
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 449801 501326 449867 501329
rect 449801 501324 450156 501326
rect 449801 501268 449806 501324
rect 449862 501296 450156 501324
rect 449862 501268 450186 501296
rect 449801 501266 450186 501268
rect 449801 501263 449867 501266
rect 450126 500986 450186 501266
rect 491894 501258 491954 501840
rect 494053 501258 494119 501261
rect 489870 501256 494119 501258
rect 489870 501200 494058 501256
rect 494114 501200 494119 501256
rect 489870 501198 494119 501200
rect 489870 501122 489930 501198
rect 494053 501195 494119 501198
rect 470550 501062 489930 501122
rect 470550 500986 470610 501062
rect 450126 500926 470610 500986
rect 448094 500244 448100 500308
rect 448164 500306 448170 500308
rect 448513 500306 448579 500309
rect 448164 500304 448579 500306
rect 448164 500248 448518 500304
rect 448574 500248 448579 500304
rect 448164 500246 448579 500248
rect 448164 500244 448170 500246
rect 448513 500243 448579 500246
rect 583520 497844 584960 498084
rect 481817 496908 481883 496909
rect 481766 496906 481772 496908
rect 481726 496846 481772 496906
rect 481836 496904 481883 496908
rect 481878 496848 481883 496904
rect 481766 496844 481772 496846
rect 481836 496844 481883 496848
rect 483054 496844 483060 496908
rect 483124 496906 483130 496908
rect 483841 496906 483907 496909
rect 483124 496904 483907 496906
rect 483124 496848 483846 496904
rect 483902 496848 483907 496904
rect 483124 496846 483907 496848
rect 483124 496844 483130 496846
rect 481817 496843 481883 496844
rect 483841 496843 483907 496846
rect 448278 496028 448284 496092
rect 448348 496090 448354 496092
rect 448421 496090 448487 496093
rect 448348 496088 448487 496090
rect 448348 496032 448426 496088
rect 448482 496032 448487 496088
rect 448348 496030 448487 496032
rect 448348 496028 448354 496030
rect 448421 496027 448487 496030
rect 361757 491738 361823 491741
rect 359812 491736 361823 491738
rect 359812 491680 361762 491736
rect 361818 491680 361823 491736
rect 359812 491678 361823 491680
rect 361757 491675 361823 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 583520 471324 584960 471414
rect 362217 469706 362283 469709
rect 359812 469704 362283 469706
rect 359812 469648 362222 469704
rect 362278 469648 362283 469704
rect 359812 469646 362283 469648
rect 362217 469643 362283 469646
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 580533 458146 580599 458149
rect 583520 458146 584960 458236
rect 580533 458144 584960 458146
rect 580533 458088 580538 458144
rect 580594 458088 584960 458144
rect 580533 458086 584960 458088
rect 580533 458083 580599 458086
rect 583520 457996 584960 458086
rect 487102 453868 487108 453932
rect 487172 453930 487178 453932
rect 487981 453930 488047 453933
rect 487172 453928 488047 453930
rect 487172 453872 487986 453928
rect 488042 453872 488047 453928
rect 487172 453870 488047 453872
rect 487172 453868 487178 453870
rect 487981 453867 488047 453870
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 362309 447674 362375 447677
rect 359812 447672 362375 447674
rect 359812 447616 362314 447672
rect 362370 447616 362375 447672
rect 359812 447614 362375 447616
rect 362309 447611 362375 447614
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 361757 436658 361823 436661
rect 359812 436656 361823 436658
rect 359812 436600 361762 436656
rect 361818 436600 361823 436656
rect 359812 436598 361823 436600
rect 361757 436595 361823 436598
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect 362401 425642 362467 425645
rect 359812 425640 362467 425642
rect 359812 425584 362406 425640
rect 362462 425584 362467 425640
rect 359812 425582 362467 425584
rect 362401 425579 362467 425582
rect -960 423602 480 423692
rect 3693 423602 3759 423605
rect -960 423600 3759 423602
rect -960 423544 3698 423600
rect 3754 423544 3759 423600
rect -960 423542 3759 423544
rect -960 423452 480 423542
rect 3693 423539 3759 423542
rect 455086 422922 455092 422924
rect 444238 422862 455092 422922
rect 444238 422109 444298 422862
rect 455086 422860 455092 422862
rect 455156 422860 455162 422924
rect 444189 422104 444298 422109
rect 444189 422048 444194 422104
rect 444250 422048 444298 422104
rect 444189 422046 444298 422048
rect 444189 422043 444255 422046
rect 443494 421908 443500 421972
rect 443564 421970 443570 421972
rect 444097 421970 444163 421973
rect 443564 421968 444163 421970
rect 443564 421912 444102 421968
rect 444158 421912 444163 421968
rect 443564 421910 444163 421912
rect 443564 421908 443570 421910
rect 444097 421907 444163 421910
rect 444046 421772 444052 421836
rect 444116 421834 444122 421836
rect 444373 421834 444439 421837
rect 444116 421832 444439 421834
rect 444116 421776 444378 421832
rect 444434 421776 444439 421832
rect 444116 421774 444439 421776
rect 444116 421772 444122 421774
rect 444373 421771 444439 421774
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 459134 410484 459140 410548
rect 459204 410546 459210 410548
rect 471973 410546 472039 410549
rect 459204 410544 472039 410546
rect 459204 410488 471978 410544
rect 472034 410488 472039 410544
rect 459204 410486 472039 410488
rect 459204 410484 459210 410486
rect 471973 410483 472039 410486
rect 580625 404970 580691 404973
rect 583520 404970 584960 405060
rect 580625 404968 584960 404970
rect 580625 404912 580630 404968
rect 580686 404912 584960 404968
rect 580625 404910 584960 404912
rect 580625 404907 580691 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3877 397490 3943 397493
rect -960 397488 3943 397490
rect -960 397432 3882 397488
rect 3938 397432 3943 397488
rect -960 397430 3943 397432
rect -960 397340 480 397430
rect 3877 397427 3943 397430
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 583520 391628 584960 391868
rect 449065 389874 449131 389877
rect 483054 389874 483060 389876
rect 449065 389872 483060 389874
rect 449065 389816 449070 389872
rect 449126 389816 483060 389872
rect 449065 389814 483060 389816
rect 449065 389811 449131 389814
rect 483054 389812 483060 389814
rect 483124 389812 483130 389876
rect 472014 388996 472020 389060
rect 472084 389058 472090 389060
rect 472893 389058 472959 389061
rect 474365 389060 474431 389061
rect 474365 389058 474412 389060
rect 472084 389056 472959 389058
rect 472084 389000 472898 389056
rect 472954 389000 472959 389056
rect 472084 388998 472959 389000
rect 474320 389056 474412 389058
rect 474320 389000 474370 389056
rect 474320 388998 474412 389000
rect 472084 388996 472090 388998
rect 472893 388995 472959 388998
rect 474365 388996 474412 388998
rect 474476 388996 474482 389060
rect 474958 388996 474964 389060
rect 475028 389058 475034 389060
rect 475101 389058 475167 389061
rect 475028 389056 475167 389058
rect 475028 389000 475106 389056
rect 475162 389000 475167 389056
rect 475028 388998 475167 389000
rect 475028 388996 475034 388998
rect 474365 388995 474431 388996
rect 475101 388995 475167 388998
rect 476430 388996 476436 389060
rect 476500 389058 476506 389060
rect 477309 389058 477375 389061
rect 476500 389056 477375 389058
rect 476500 389000 477314 389056
rect 477370 389000 477375 389056
rect 476500 388998 477375 389000
rect 476500 388996 476506 388998
rect 477309 388995 477375 388998
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 479517 388995 479583 388998
rect 473629 388922 473695 388925
rect 474590 388922 474596 388924
rect 473629 388920 474596 388922
rect 473629 388864 473634 388920
rect 473690 388864 474596 388920
rect 473629 388862 474596 388864
rect 473629 388859 473695 388862
rect 474590 388860 474596 388862
rect 474660 388860 474666 388924
rect 474774 388860 474780 388924
rect 474844 388922 474850 388924
rect 475837 388922 475903 388925
rect 474844 388920 475903 388922
rect 474844 388864 475842 388920
rect 475898 388864 475903 388920
rect 474844 388862 475903 388864
rect 474844 388860 474850 388862
rect 475837 388859 475903 388862
rect 442809 387154 442875 387157
rect 453246 387154 453252 387156
rect 442809 387152 453252 387154
rect 442809 387096 442814 387152
rect 442870 387096 453252 387152
rect 442809 387094 453252 387096
rect 442809 387091 442875 387094
rect 453246 387092 453252 387094
rect 453316 387092 453322 387156
rect 448973 387018 449039 387021
rect 481766 387018 481772 387020
rect 448973 387016 481772 387018
rect 448973 386960 448978 387016
rect 449034 386960 481772 387016
rect 448973 386958 481772 386960
rect 448973 386955 449039 386958
rect 481766 386956 481772 386958
rect 481836 386956 481842 387020
rect 449249 385658 449315 385661
rect 487102 385658 487108 385660
rect 449249 385656 487108 385658
rect 449249 385600 449254 385656
rect 449310 385600 487108 385656
rect 449249 385598 487108 385600
rect 449249 385595 449315 385598
rect 487102 385596 487108 385598
rect 487172 385596 487178 385660
rect 512729 384706 512795 384709
rect 509956 384704 512795 384706
rect 509956 384648 512734 384704
rect 512790 384648 512795 384704
rect 509956 384646 512795 384648
rect 512729 384643 512795 384646
rect -960 384284 480 384524
rect 513281 384162 513347 384165
rect 509956 384160 513347 384162
rect 509956 384104 513286 384160
rect 513342 384104 513347 384160
rect 509956 384102 513347 384104
rect 513281 384099 513347 384102
rect 447133 383890 447199 383893
rect 447133 383888 450156 383890
rect 447133 383832 447138 383888
rect 447194 383832 450156 383888
rect 447133 383830 450156 383832
rect 447133 383827 447199 383830
rect 512913 383618 512979 383621
rect 509956 383616 512979 383618
rect 509956 383560 512918 383616
rect 512974 383560 512979 383616
rect 509956 383558 512979 383560
rect 512913 383555 512979 383558
rect 447133 383210 447199 383213
rect 447133 383208 450156 383210
rect 447133 383152 447138 383208
rect 447194 383152 450156 383208
rect 447133 383150 450156 383152
rect 447133 383147 447199 383150
rect 513281 383074 513347 383077
rect 509956 383072 513347 383074
rect 509956 383016 513286 383072
rect 513342 383016 513347 383072
rect 509956 383014 513347 383016
rect 513281 383011 513347 383014
rect 447225 382530 447291 382533
rect 513189 382530 513255 382533
rect 447225 382528 450156 382530
rect 447225 382472 447230 382528
rect 447286 382472 450156 382528
rect 447225 382470 450156 382472
rect 509956 382528 513255 382530
rect 509956 382472 513194 382528
rect 513250 382472 513255 382528
rect 509956 382470 513255 382472
rect 447225 382467 447291 382470
rect 513189 382467 513255 382470
rect 512361 381986 512427 381989
rect 509956 381984 512427 381986
rect 509956 381928 512366 381984
rect 512422 381928 512427 381984
rect 509956 381926 512427 381928
rect 512361 381923 512427 381926
rect 447133 381850 447199 381853
rect 447133 381848 450156 381850
rect 447133 381792 447138 381848
rect 447194 381792 450156 381848
rect 447133 381790 450156 381792
rect 447133 381787 447199 381790
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 513281 381442 513347 381445
rect 509956 381440 513347 381442
rect 509956 381384 513286 381440
rect 513342 381384 513347 381440
rect 509956 381382 513347 381384
rect 513281 381379 513347 381382
rect 447225 381170 447291 381173
rect 447225 381168 450156 381170
rect 447225 381112 447230 381168
rect 447286 381112 450156 381168
rect 447225 381110 450156 381112
rect 447225 381107 447291 381110
rect 512361 380898 512427 380901
rect 509956 380896 512427 380898
rect 509956 380840 512366 380896
rect 512422 380840 512427 380896
rect 509956 380838 512427 380840
rect 512361 380835 512427 380838
rect 447133 380490 447199 380493
rect 447133 380488 450156 380490
rect 447133 380432 447138 380488
rect 447194 380432 450156 380488
rect 447133 380430 450156 380432
rect 447133 380427 447199 380430
rect 512085 380354 512151 380357
rect 509956 380352 512151 380354
rect 509956 380296 512090 380352
rect 512146 380296 512151 380352
rect 509956 380294 512151 380296
rect 512085 380291 512151 380294
rect 447225 379810 447291 379813
rect 512821 379810 512887 379813
rect 447225 379808 450156 379810
rect 447225 379752 447230 379808
rect 447286 379752 450156 379808
rect 447225 379750 450156 379752
rect 509956 379808 512887 379810
rect 509956 379752 512826 379808
rect 512882 379752 512887 379808
rect 509956 379750 512887 379752
rect 447225 379747 447291 379750
rect 512821 379747 512887 379750
rect 513281 379266 513347 379269
rect 509956 379264 513347 379266
rect 509956 379208 513286 379264
rect 513342 379208 513347 379264
rect 509956 379206 513347 379208
rect 513281 379203 513347 379206
rect 447133 379130 447199 379133
rect 447133 379128 450156 379130
rect 447133 379072 447138 379128
rect 447194 379072 450156 379128
rect 447133 379070 450156 379072
rect 447133 379067 447199 379070
rect 512177 378722 512243 378725
rect 509956 378720 512243 378722
rect 509956 378664 512182 378720
rect 512238 378664 512243 378720
rect 509956 378662 512243 378664
rect 512177 378659 512243 378662
rect 447225 378450 447291 378453
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 447225 378448 450156 378450
rect 447225 378392 447230 378448
rect 447286 378392 450156 378448
rect 447225 378390 450156 378392
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 447225 378387 447291 378390
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect 511993 378178 512059 378181
rect 509956 378176 512059 378178
rect 509956 378120 511998 378176
rect 512054 378120 512059 378176
rect 509956 378118 512059 378120
rect 511993 378115 512059 378118
rect 447133 377770 447199 377773
rect 447133 377768 450156 377770
rect 447133 377712 447138 377768
rect 447194 377712 450156 377768
rect 447133 377710 450156 377712
rect 447133 377707 447199 377710
rect 512085 377634 512151 377637
rect 509956 377632 512151 377634
rect 509956 377576 512090 377632
rect 512146 377576 512151 377632
rect 509956 377574 512151 377576
rect 512085 377571 512151 377574
rect 447225 377090 447291 377093
rect 513189 377090 513255 377093
rect 447225 377088 450156 377090
rect 447225 377032 447230 377088
rect 447286 377032 450156 377088
rect 447225 377030 450156 377032
rect 509956 377088 513255 377090
rect 509956 377032 513194 377088
rect 513250 377032 513255 377088
rect 509956 377030 513255 377032
rect 447225 377027 447291 377030
rect 513189 377027 513255 377030
rect 512177 376546 512243 376549
rect 509956 376544 512243 376546
rect 509956 376488 512182 376544
rect 512238 376488 512243 376544
rect 509956 376486 512243 376488
rect 512177 376483 512243 376486
rect 447133 376410 447199 376413
rect 447133 376408 450156 376410
rect 447133 376352 447138 376408
rect 447194 376352 450156 376408
rect 447133 376350 450156 376352
rect 447133 376347 447199 376350
rect 512269 376002 512335 376005
rect 509956 376000 512335 376002
rect 509956 375944 512274 376000
rect 512330 375944 512335 376000
rect 509956 375942 512335 375944
rect 512269 375939 512335 375942
rect 447225 375730 447291 375733
rect 447225 375728 450156 375730
rect 447225 375672 447230 375728
rect 447286 375672 450156 375728
rect 447225 375670 450156 375672
rect 447225 375667 447291 375670
rect 513281 375458 513347 375461
rect 509956 375456 513347 375458
rect 509956 375400 513286 375456
rect 513342 375400 513347 375456
rect 509956 375398 513347 375400
rect 513281 375395 513347 375398
rect 447133 375050 447199 375053
rect 447133 375048 450156 375050
rect 447133 374992 447138 375048
rect 447194 374992 450156 375048
rect 447133 374990 450156 374992
rect 447133 374987 447199 374990
rect 512453 374914 512519 374917
rect 509956 374912 512519 374914
rect 509956 374856 512458 374912
rect 512514 374856 512519 374912
rect 509956 374854 512519 374856
rect 512453 374851 512519 374854
rect 447225 374370 447291 374373
rect 512729 374370 512795 374373
rect 447225 374368 450156 374370
rect 447225 374312 447230 374368
rect 447286 374312 450156 374368
rect 447225 374310 450156 374312
rect 509956 374368 512795 374370
rect 509956 374312 512734 374368
rect 512790 374312 512795 374368
rect 509956 374310 512795 374312
rect 447225 374307 447291 374310
rect 512729 374307 512795 374310
rect 512821 373826 512887 373829
rect 509956 373824 512887 373826
rect 509956 373768 512826 373824
rect 512882 373768 512887 373824
rect 509956 373766 512887 373768
rect 512821 373763 512887 373766
rect 447133 373690 447199 373693
rect 447133 373688 450156 373690
rect 447133 373632 447138 373688
rect 447194 373632 450156 373688
rect 447133 373630 450156 373632
rect 447133 373627 447199 373630
rect 513281 373282 513347 373285
rect 509956 373280 513347 373282
rect 509956 373224 513286 373280
rect 513342 373224 513347 373280
rect 509956 373222 513347 373224
rect 513281 373219 513347 373222
rect 447225 373010 447291 373013
rect 447225 373008 450156 373010
rect 447225 372952 447230 373008
rect 447286 372952 450156 373008
rect 447225 372950 450156 372952
rect 447225 372947 447291 372950
rect 509558 372469 509618 372708
rect 509558 372464 509667 372469
rect 509558 372408 509606 372464
rect 509662 372408 509667 372464
rect 509558 372406 509667 372408
rect 509601 372403 509667 372406
rect 447133 372330 447199 372333
rect 447133 372328 450156 372330
rect 447133 372272 447138 372328
rect 447194 372272 450156 372328
rect 447133 372270 450156 372272
rect 447133 372267 447199 372270
rect 512545 372194 512611 372197
rect 509956 372192 512611 372194
rect 509956 372136 512550 372192
rect 512606 372136 512611 372192
rect 509956 372134 512611 372136
rect 512545 372131 512611 372134
rect 447225 371650 447291 371653
rect 512269 371650 512335 371653
rect 447225 371648 450156 371650
rect 447225 371592 447230 371648
rect 447286 371592 450156 371648
rect 447225 371590 450156 371592
rect 509956 371648 512335 371650
rect 509956 371592 512274 371648
rect 512330 371592 512335 371648
rect 509956 371590 512335 371592
rect 447225 371587 447291 371590
rect 512269 371587 512335 371590
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 511993 371106 512059 371109
rect 509956 371104 512059 371106
rect 509956 371048 511998 371104
rect 512054 371048 512059 371104
rect 509956 371046 512059 371048
rect 511993 371043 512059 371046
rect 447133 370970 447199 370973
rect 447133 370968 450156 370970
rect 447133 370912 447138 370968
rect 447194 370912 450156 370968
rect 447133 370910 450156 370912
rect 447133 370907 447199 370910
rect 361573 370562 361639 370565
rect 512085 370562 512151 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 509956 370560 512151 370562
rect 509956 370504 512090 370560
rect 512146 370504 512151 370560
rect 509956 370502 512151 370504
rect 361573 370499 361639 370502
rect 512085 370499 512151 370502
rect 447225 370290 447291 370293
rect 447225 370288 450156 370290
rect 447225 370232 447230 370288
rect 447286 370232 450156 370288
rect 447225 370230 450156 370232
rect 447225 370227 447291 370230
rect 513281 370018 513347 370021
rect 509956 370016 513347 370018
rect 509956 369960 513286 370016
rect 513342 369960 513347 370016
rect 509956 369958 513347 369960
rect 513281 369955 513347 369958
rect 447133 369610 447199 369613
rect 447133 369608 450156 369610
rect 447133 369552 447138 369608
rect 447194 369552 450156 369608
rect 447133 369550 450156 369552
rect 447133 369547 447199 369550
rect 513005 369474 513071 369477
rect 509956 369472 513071 369474
rect 509956 369416 513010 369472
rect 513066 369416 513071 369472
rect 509956 369414 513071 369416
rect 513005 369411 513071 369414
rect 447225 368930 447291 368933
rect 510705 368930 510771 368933
rect 447225 368928 450156 368930
rect 447225 368872 447230 368928
rect 447286 368872 450156 368928
rect 447225 368870 450156 368872
rect 509956 368928 510771 368930
rect 509956 368872 510710 368928
rect 510766 368872 510771 368928
rect 509956 368870 510771 368872
rect 447225 368867 447291 368870
rect 510705 368867 510771 368870
rect 512361 368386 512427 368389
rect 509956 368384 512427 368386
rect 509956 368328 512366 368384
rect 512422 368328 512427 368384
rect 509956 368326 512427 368328
rect 512361 368323 512427 368326
rect 447133 368250 447199 368253
rect 447133 368248 450156 368250
rect 447133 368192 447138 368248
rect 447194 368192 450156 368248
rect 447133 368190 450156 368192
rect 447133 368187 447199 368190
rect 512637 367842 512703 367845
rect 509956 367840 512703 367842
rect 509956 367784 512642 367840
rect 512698 367784 512703 367840
rect 509956 367782 512703 367784
rect 512637 367779 512703 367782
rect 447225 367570 447291 367573
rect 447225 367568 450156 367570
rect 447225 367512 447230 367568
rect 447286 367512 450156 367568
rect 447225 367510 450156 367512
rect 447225 367507 447291 367510
rect 509374 367029 509434 367268
rect 509325 367024 509434 367029
rect 509325 366968 509330 367024
rect 509386 366968 509434 367024
rect 509325 366966 509434 366968
rect 509325 366963 509391 366966
rect 447133 366890 447199 366893
rect 447133 366888 450156 366890
rect 447133 366832 447138 366888
rect 447194 366832 450156 366888
rect 447133 366830 450156 366832
rect 447133 366827 447199 366830
rect 510613 366754 510679 366757
rect 509956 366752 510679 366754
rect 509956 366696 510618 366752
rect 510674 366696 510679 366752
rect 509956 366694 510679 366696
rect 510613 366691 510679 366694
rect 447225 366210 447291 366213
rect 512453 366210 512519 366213
rect 447225 366208 450156 366210
rect 447225 366152 447230 366208
rect 447286 366152 450156 366208
rect 447225 366150 450156 366152
rect 509956 366208 512519 366210
rect 509956 366152 512458 366208
rect 512514 366152 512519 366208
rect 509956 366150 512519 366152
rect 447225 366147 447291 366150
rect 512453 366147 512519 366150
rect 513557 365666 513623 365669
rect 509956 365664 513623 365666
rect 509956 365608 513562 365664
rect 513618 365608 513623 365664
rect 509956 365606 513623 365608
rect 513557 365603 513623 365606
rect 447225 365530 447291 365533
rect 447225 365528 450156 365530
rect 447225 365472 447230 365528
rect 447286 365472 450156 365528
rect 447225 365470 450156 365472
rect 447225 365467 447291 365470
rect 512453 365122 512519 365125
rect 509956 365120 512519 365122
rect 509956 365064 512458 365120
rect 512514 365064 512519 365120
rect 509956 365062 512519 365064
rect 512453 365059 512519 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364850 447199 364853
rect 447133 364848 450156 364850
rect 447133 364792 447138 364848
rect 447194 364792 450156 364848
rect 447133 364790 450156 364792
rect 447133 364787 447199 364790
rect 512085 364578 512151 364581
rect 509956 364576 512151 364578
rect 509956 364520 512090 364576
rect 512146 364520 512151 364576
rect 509956 364518 512151 364520
rect 512085 364515 512151 364518
rect 447133 364170 447199 364173
rect 447133 364168 450156 364170
rect 447133 364112 447138 364168
rect 447194 364112 450156 364168
rect 447133 364110 450156 364112
rect 447133 364107 447199 364110
rect 511993 364034 512059 364037
rect 509956 364032 512059 364034
rect 509956 363976 511998 364032
rect 512054 363976 512059 364032
rect 509956 363974 512059 363976
rect 511993 363971 512059 363974
rect 447225 363490 447291 363493
rect 513281 363490 513347 363493
rect 447225 363488 450156 363490
rect 447225 363432 447230 363488
rect 447286 363432 450156 363488
rect 447225 363430 450156 363432
rect 509956 363488 513347 363490
rect 509956 363432 513286 363488
rect 513342 363432 513347 363488
rect 509956 363430 513347 363432
rect 447225 363427 447291 363430
rect 513281 363427 513347 363430
rect 513281 362946 513347 362949
rect 509956 362944 513347 362946
rect 509956 362888 513286 362944
rect 513342 362888 513347 362944
rect 509956 362886 513347 362888
rect 513281 362883 513347 362886
rect 447225 362810 447291 362813
rect 447225 362808 450156 362810
rect 447225 362752 447230 362808
rect 447286 362752 450156 362808
rect 447225 362750 450156 362752
rect 447225 362747 447291 362750
rect 511993 362402 512059 362405
rect 509956 362400 512059 362402
rect 509956 362344 511998 362400
rect 512054 362344 512059 362400
rect 509956 362342 512059 362344
rect 511993 362339 512059 362342
rect 447133 362130 447199 362133
rect 447133 362128 450156 362130
rect 447133 362072 447138 362128
rect 447194 362072 450156 362128
rect 447133 362070 450156 362072
rect 447133 362067 447199 362070
rect 513097 361858 513163 361861
rect 509956 361856 513163 361858
rect 509956 361800 513102 361856
rect 513158 361800 513163 361856
rect 509956 361798 513163 361800
rect 513097 361795 513163 361798
rect 447225 361450 447291 361453
rect 447225 361448 450156 361450
rect 447225 361392 447230 361448
rect 447286 361392 450156 361448
rect 447225 361390 450156 361392
rect 447225 361387 447291 361390
rect 513281 361314 513347 361317
rect 509956 361312 513347 361314
rect 509956 361256 513286 361312
rect 513342 361256 513347 361312
rect 509956 361254 513347 361256
rect 513281 361251 513347 361254
rect 447133 360770 447199 360773
rect 510797 360770 510863 360773
rect 447133 360768 450156 360770
rect 447133 360712 447138 360768
rect 447194 360712 450156 360768
rect 447133 360710 450156 360712
rect 509956 360768 510863 360770
rect 509956 360712 510802 360768
rect 510858 360712 510863 360768
rect 509956 360710 510863 360712
rect 447133 360707 447199 360710
rect 510797 360707 510863 360710
rect 512545 360226 512611 360229
rect 509956 360224 512611 360226
rect 509956 360168 512550 360224
rect 512606 360168 512611 360224
rect 509956 360166 512611 360168
rect 512545 360163 512611 360166
rect 447225 360090 447291 360093
rect 447225 360088 450156 360090
rect 447225 360032 447230 360088
rect 447286 360032 450156 360088
rect 447225 360030 450156 360032
rect 447225 360027 447291 360030
rect 513281 359682 513347 359685
rect 509956 359680 513347 359682
rect 509956 359624 513286 359680
rect 513342 359624 513347 359680
rect 509956 359622 513347 359624
rect 513281 359619 513347 359622
rect 362217 359546 362283 359549
rect 359812 359544 362283 359546
rect 359812 359488 362222 359544
rect 362278 359488 362283 359544
rect 359812 359486 362283 359488
rect 362217 359483 362283 359486
rect 447133 359410 447199 359413
rect 447133 359408 450156 359410
rect 447133 359352 447138 359408
rect 447194 359352 450156 359408
rect 447133 359350 450156 359352
rect 447133 359347 447199 359350
rect 509374 358869 509434 359108
rect 450261 358866 450327 358869
rect 450261 358864 450370 358866
rect 450261 358808 450266 358864
rect 450322 358808 450370 358864
rect 450261 358803 450370 358808
rect 509374 358864 509483 358869
rect 509374 358808 509422 358864
rect 509478 358808 509483 358864
rect 509374 358806 509483 358808
rect 509417 358803 509483 358806
rect 450310 358700 450370 358803
rect 511993 358594 512059 358597
rect 509956 358592 512059 358594
rect -960 358458 480 358548
rect 509956 358536 511998 358592
rect 512054 358536 512059 358592
rect 509956 358534 512059 358536
rect 511993 358531 512059 358534
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 450077 358458 450143 358461
rect 450077 358456 450186 358458
rect 450077 358400 450082 358456
rect 450138 358400 450186 358456
rect 450077 358395 450186 358400
rect 450126 358020 450186 358395
rect 512085 358050 512151 358053
rect 509956 358048 512151 358050
rect 509956 357992 512090 358048
rect 512146 357992 512151 358048
rect 509956 357990 512151 357992
rect 512085 357987 512151 357990
rect 512085 357506 512151 357509
rect 509956 357504 512151 357506
rect 509956 357448 512090 357504
rect 512146 357448 512151 357504
rect 509956 357446 512151 357448
rect 512085 357443 512151 357446
rect 449617 357370 449683 357373
rect 449617 357368 450156 357370
rect 449617 357312 449622 357368
rect 449678 357312 450156 357368
rect 449617 357310 450156 357312
rect 449617 357307 449683 357310
rect 512729 356962 512795 356965
rect 509956 356960 512795 356962
rect 509956 356904 512734 356960
rect 512790 356904 512795 356960
rect 509956 356902 512795 356904
rect 512729 356899 512795 356902
rect 449433 356690 449499 356693
rect 449433 356688 450156 356690
rect 449433 356632 449438 356688
rect 449494 356632 450156 356688
rect 449433 356630 450156 356632
rect 449433 356627 449499 356630
rect 512085 356418 512151 356421
rect 509956 356416 512151 356418
rect 509956 356360 512090 356416
rect 512146 356360 512151 356416
rect 509956 356358 512151 356360
rect 512085 356355 512151 356358
rect 449709 356010 449775 356013
rect 449709 356008 450156 356010
rect 449709 355952 449714 356008
rect 449770 355952 450156 356008
rect 449709 355950 450156 355952
rect 449709 355947 449775 355950
rect 510889 355874 510955 355877
rect 509956 355872 510955 355874
rect 509956 355816 510894 355872
rect 510950 355816 510955 355872
rect 509956 355814 510955 355816
rect 510889 355811 510955 355814
rect 449341 355330 449407 355333
rect 513189 355330 513255 355333
rect 449341 355328 450156 355330
rect 449341 355272 449346 355328
rect 449402 355272 450156 355328
rect 449341 355270 450156 355272
rect 509956 355328 513255 355330
rect 509956 355272 513194 355328
rect 513250 355272 513255 355328
rect 509956 355270 513255 355272
rect 449341 355267 449407 355270
rect 513189 355267 513255 355270
rect 513281 354786 513347 354789
rect 509956 354784 513347 354786
rect 509956 354728 513286 354784
rect 513342 354728 513347 354784
rect 509956 354726 513347 354728
rect 513281 354723 513347 354726
rect 449065 354650 449131 354653
rect 449065 354648 450156 354650
rect 449065 354592 449070 354648
rect 449126 354592 450156 354648
rect 449065 354590 450156 354592
rect 449065 354587 449131 354590
rect 512085 354242 512151 354245
rect 509956 354240 512151 354242
rect 509956 354184 512090 354240
rect 512146 354184 512151 354240
rect 509956 354182 512151 354184
rect 512085 354179 512151 354182
rect 449525 353970 449591 353973
rect 449525 353968 450156 353970
rect 449525 353912 449530 353968
rect 449586 353912 450156 353968
rect 449525 353910 450156 353912
rect 449525 353907 449591 353910
rect 513281 353698 513347 353701
rect 509956 353696 513347 353698
rect 509956 353640 513286 353696
rect 513342 353640 513347 353696
rect 509956 353638 513347 353640
rect 513281 353635 513347 353638
rect 448973 353290 449039 353293
rect 448973 353288 450156 353290
rect 448973 353232 448978 353288
rect 449034 353232 450156 353288
rect 448973 353230 450156 353232
rect 448973 353227 449039 353230
rect 512913 353154 512979 353157
rect 509956 353152 512979 353154
rect 509956 353096 512918 353152
rect 512974 353096 512979 353152
rect 509956 353094 512979 353096
rect 512913 353091 512979 353094
rect 447593 352610 447659 352613
rect 510981 352610 511047 352613
rect 447593 352608 450156 352610
rect 447593 352552 447598 352608
rect 447654 352552 450156 352608
rect 447593 352550 450156 352552
rect 509956 352608 511047 352610
rect 509956 352552 510986 352608
rect 511042 352552 511047 352608
rect 509956 352550 511047 352552
rect 447593 352547 447659 352550
rect 510981 352547 511047 352550
rect 513281 352066 513347 352069
rect 509956 352064 513347 352066
rect 509956 352008 513286 352064
rect 513342 352008 513347 352064
rect 509956 352006 513347 352008
rect 513281 352003 513347 352006
rect 447133 351930 447199 351933
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 447133 351928 450156 351930
rect 447133 351872 447138 351928
rect 447194 351872 450156 351928
rect 447133 351870 450156 351872
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 447133 351867 447199 351870
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect 512821 351522 512887 351525
rect 509956 351520 512887 351522
rect 509956 351464 512826 351520
rect 512882 351464 512887 351520
rect 509956 351462 512887 351464
rect 512821 351459 512887 351462
rect 447409 351250 447475 351253
rect 447409 351248 450156 351250
rect 447409 351192 447414 351248
rect 447470 351192 450156 351248
rect 447409 351190 450156 351192
rect 447409 351187 447475 351190
rect 512085 350978 512151 350981
rect 509956 350976 512151 350978
rect 509956 350920 512090 350976
rect 512146 350920 512151 350976
rect 509956 350918 512151 350920
rect 512085 350915 512151 350918
rect 447133 350570 447199 350573
rect 447133 350568 450156 350570
rect 447133 350512 447138 350568
rect 447194 350512 450156 350568
rect 447133 350510 450156 350512
rect 447133 350507 447199 350510
rect 513005 350434 513071 350437
rect 509956 350432 513071 350434
rect 509956 350376 513010 350432
rect 513066 350376 513071 350432
rect 509956 350374 513071 350376
rect 513005 350371 513071 350374
rect 449709 349890 449775 349893
rect 449709 349888 450156 349890
rect 449709 349832 449714 349888
rect 449770 349832 450156 349888
rect 449709 349830 450156 349832
rect 449709 349827 449775 349830
rect 509558 349485 509618 349860
rect 509509 349480 509618 349485
rect 509509 349424 509514 349480
rect 509570 349424 509618 349480
rect 509509 349422 509618 349424
rect 509509 349419 509575 349422
rect 512085 349346 512151 349349
rect 509956 349344 512151 349346
rect 509956 349288 512090 349344
rect 512146 349288 512151 349344
rect 509956 349286 512151 349288
rect 512085 349283 512151 349286
rect 448421 349210 448487 349213
rect 448421 349208 450156 349210
rect 448421 349152 448426 349208
rect 448482 349152 450156 349208
rect 448421 349150 450156 349152
rect 448421 349147 448487 349150
rect 512821 348802 512887 348805
rect 509956 348800 512887 348802
rect 509956 348744 512826 348800
rect 512882 348744 512887 348800
rect 509956 348742 512887 348744
rect 512821 348739 512887 348742
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 447777 348530 447843 348533
rect 447777 348528 450156 348530
rect 447777 348472 447782 348528
rect 447838 348472 450156 348528
rect 447777 348470 450156 348472
rect 447777 348467 447843 348470
rect 512913 348258 512979 348261
rect 509956 348256 512979 348258
rect 509956 348200 512918 348256
rect 512974 348200 512979 348256
rect 509956 348198 512979 348200
rect 512913 348195 512979 348198
rect 447685 347850 447751 347853
rect 447685 347848 450156 347850
rect 447685 347792 447690 347848
rect 447746 347792 450156 347848
rect 447685 347790 450156 347792
rect 447685 347787 447751 347790
rect 512637 347714 512703 347717
rect 509956 347712 512703 347714
rect 509956 347656 512642 347712
rect 512698 347656 512703 347712
rect 509956 347654 512703 347656
rect 512637 347651 512703 347654
rect 447133 347170 447199 347173
rect 513281 347170 513347 347173
rect 447133 347168 450156 347170
rect 447133 347112 447138 347168
rect 447194 347112 450156 347168
rect 447133 347110 450156 347112
rect 509956 347168 513347 347170
rect 509956 347112 513286 347168
rect 513342 347112 513347 347168
rect 509956 347110 513347 347112
rect 447133 347107 447199 347110
rect 513281 347107 513347 347110
rect 449893 346898 449959 346901
rect 449893 346896 450186 346898
rect 449893 346840 449898 346896
rect 449954 346840 450186 346896
rect 449893 346838 450186 346840
rect 449893 346835 449959 346838
rect 450126 346460 450186 346838
rect 512821 346626 512887 346629
rect 509956 346624 512887 346626
rect 509956 346568 512826 346624
rect 512882 346568 512887 346624
rect 509956 346566 512887 346568
rect 512821 346563 512887 346566
rect 512085 346082 512151 346085
rect 509956 346080 512151 346082
rect 509956 346024 512090 346080
rect 512146 346024 512151 346080
rect 509956 346022 512151 346024
rect 512085 346019 512151 346022
rect 449801 345810 449867 345813
rect 449801 345808 450156 345810
rect 449801 345752 449806 345808
rect 449862 345752 450156 345808
rect 449801 345750 450156 345752
rect 449801 345747 449867 345750
rect 512085 345538 512151 345541
rect 509956 345536 512151 345538
rect -960 345402 480 345492
rect 509956 345480 512090 345536
rect 512146 345480 512151 345536
rect 509956 345478 512151 345480
rect 512085 345475 512151 345478
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 449801 345130 449867 345133
rect 449801 345128 450156 345130
rect 449801 345072 449806 345128
rect 449862 345072 450156 345128
rect 449801 345070 450156 345072
rect 449801 345067 449867 345070
rect 513281 344994 513347 344997
rect 509956 344992 513347 344994
rect 509956 344936 513286 344992
rect 513342 344936 513347 344992
rect 509956 344934 513347 344936
rect 513281 344931 513347 344934
rect 447593 344450 447659 344453
rect 512637 344450 512703 344453
rect 447593 344448 450156 344450
rect 447593 344392 447598 344448
rect 447654 344392 450156 344448
rect 447593 344390 450156 344392
rect 509956 344448 512703 344450
rect 509956 344392 512642 344448
rect 512698 344392 512703 344448
rect 509956 344390 512703 344392
rect 447593 344387 447659 344390
rect 512637 344387 512703 344390
rect 512821 343906 512887 343909
rect 509956 343904 512887 343906
rect 509956 343848 512826 343904
rect 512882 343848 512887 343904
rect 509956 343846 512887 343848
rect 512821 343843 512887 343846
rect 447317 343770 447383 343773
rect 447317 343768 450156 343770
rect 447317 343712 447322 343768
rect 447378 343712 450156 343768
rect 447317 343710 450156 343712
rect 447317 343707 447383 343710
rect 511533 343362 511599 343365
rect 509956 343360 511599 343362
rect 509956 343304 511538 343360
rect 511594 343304 511599 343360
rect 509956 343302 511599 343304
rect 511533 343299 511599 343302
rect 447869 343090 447935 343093
rect 449617 343090 449683 343093
rect 447869 343088 450156 343090
rect 447869 343032 447874 343088
rect 447930 343032 449622 343088
rect 449678 343032 450156 343088
rect 447869 343030 450156 343032
rect 447869 343027 447935 343030
rect 449617 343027 449683 343030
rect 511165 342818 511231 342821
rect 509956 342816 511231 342818
rect 509956 342760 511170 342816
rect 511226 342760 511231 342816
rect 509956 342758 511231 342760
rect 511165 342755 511231 342758
rect 449157 342410 449223 342413
rect 449157 342408 450156 342410
rect 449157 342352 449162 342408
rect 449218 342352 450156 342408
rect 449157 342350 450156 342352
rect 449157 342347 449223 342350
rect 512637 342274 512703 342277
rect 509956 342272 512703 342274
rect 509956 342216 512642 342272
rect 512698 342216 512703 342272
rect 509956 342214 512703 342216
rect 512637 342211 512703 342214
rect 447133 341730 447199 341733
rect 513281 341730 513347 341733
rect 447133 341728 450156 341730
rect 447133 341672 447138 341728
rect 447194 341672 450156 341728
rect 447133 341670 450156 341672
rect 509956 341728 513347 341730
rect 509956 341672 513286 341728
rect 513342 341672 513347 341728
rect 509956 341670 513347 341672
rect 447133 341667 447199 341670
rect 513281 341667 513347 341670
rect 513005 341186 513071 341189
rect 509956 341184 513071 341186
rect 509956 341128 513010 341184
rect 513066 341128 513071 341184
rect 509956 341126 513071 341128
rect 513005 341123 513071 341126
rect 447225 341050 447291 341053
rect 447225 341048 450156 341050
rect 447225 340992 447230 341048
rect 447286 340992 450156 341048
rect 447225 340990 450156 340992
rect 447225 340987 447291 340990
rect 513189 340642 513255 340645
rect 509956 340640 513255 340642
rect 509956 340584 513194 340640
rect 513250 340584 513255 340640
rect 509956 340582 513255 340584
rect 513189 340579 513255 340582
rect 447133 340370 447199 340373
rect 447133 340368 450156 340370
rect 447133 340312 447138 340368
rect 447194 340312 450156 340368
rect 447133 340310 450156 340312
rect 447133 340307 447199 340310
rect 513281 340098 513347 340101
rect 509956 340096 513347 340098
rect 509956 340040 513286 340096
rect 513342 340040 513347 340096
rect 509956 340038 513347 340040
rect 513281 340035 513347 340038
rect 447225 339690 447291 339693
rect 447225 339688 450156 339690
rect 447225 339632 447230 339688
rect 447286 339632 450156 339688
rect 447225 339630 450156 339632
rect 447225 339627 447291 339630
rect 513005 339554 513071 339557
rect 509956 339552 513071 339554
rect 509956 339496 513010 339552
rect 513066 339496 513071 339552
rect 509956 339494 513071 339496
rect 513005 339491 513071 339494
rect 447225 339010 447291 339013
rect 513189 339010 513255 339013
rect 447225 339008 450156 339010
rect 447225 338952 447230 339008
rect 447286 338952 450156 339008
rect 447225 338950 450156 338952
rect 509956 339008 513255 339010
rect 509956 338952 513194 339008
rect 513250 338952 513255 339008
rect 509956 338950 513255 338952
rect 447225 338947 447291 338950
rect 513189 338947 513255 338950
rect 513281 338466 513347 338469
rect 509956 338464 513347 338466
rect 509956 338408 513286 338464
rect 513342 338408 513347 338464
rect 583520 338452 584960 338692
rect 509956 338406 513347 338408
rect 513281 338403 513347 338406
rect 447133 338330 447199 338333
rect 447133 338328 450156 338330
rect 447133 338272 447138 338328
rect 447194 338272 450156 338328
rect 447133 338270 450156 338272
rect 447133 338267 447199 338270
rect 513189 337922 513255 337925
rect 509956 337920 513255 337922
rect 509956 337864 513194 337920
rect 513250 337864 513255 337920
rect 509956 337862 513255 337864
rect 513189 337859 513255 337862
rect 447225 337650 447291 337653
rect 447225 337648 450156 337650
rect 447225 337592 447230 337648
rect 447286 337592 450156 337648
rect 447225 337590 450156 337592
rect 447225 337587 447291 337590
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 513189 337378 513255 337381
rect 509956 337376 513255 337378
rect 509956 337320 513194 337376
rect 513250 337320 513255 337376
rect 509956 337318 513255 337320
rect 513189 337315 513255 337318
rect 447133 336970 447199 336973
rect 447133 336968 450156 336970
rect 447133 336912 447138 336968
rect 447194 336912 450156 336968
rect 447133 336910 450156 336912
rect 447133 336907 447199 336910
rect 513281 336834 513347 336837
rect 509956 336832 513347 336834
rect 509956 336776 513286 336832
rect 513342 336776 513347 336832
rect 509956 336774 513347 336776
rect 513281 336771 513347 336774
rect 447225 336290 447291 336293
rect 513189 336290 513255 336293
rect 447225 336288 450156 336290
rect 447225 336232 447230 336288
rect 447286 336232 450156 336288
rect 447225 336230 450156 336232
rect 509956 336288 513255 336290
rect 509956 336232 513194 336288
rect 513250 336232 513255 336288
rect 509956 336230 513255 336232
rect 447225 336227 447291 336230
rect 513189 336227 513255 336230
rect 513281 335746 513347 335749
rect 509956 335744 513347 335746
rect 509956 335688 513286 335744
rect 513342 335688 513347 335744
rect 509956 335686 513347 335688
rect 513281 335683 513347 335686
rect 447317 335610 447383 335613
rect 447317 335608 450156 335610
rect 447317 335552 447322 335608
rect 447378 335552 450156 335608
rect 447317 335550 450156 335552
rect 447317 335547 447383 335550
rect 513189 335202 513255 335205
rect 509956 335200 513255 335202
rect 509956 335144 513194 335200
rect 513250 335144 513255 335200
rect 509956 335142 513255 335144
rect 513189 335139 513255 335142
rect 447317 334930 447383 334933
rect 447317 334928 450156 334930
rect 447317 334872 447322 334928
rect 447378 334872 450156 334928
rect 447317 334870 450156 334872
rect 447317 334867 447383 334870
rect 510654 334658 510660 334660
rect 509956 334598 510660 334658
rect 510654 334596 510660 334598
rect 510724 334596 510730 334660
rect 420729 334522 420795 334525
rect 421046 334522 421052 334524
rect 420729 334520 421052 334522
rect 420729 334464 420734 334520
rect 420790 334464 421052 334520
rect 420729 334462 421052 334464
rect 420729 334459 420795 334462
rect 421046 334460 421052 334462
rect 421116 334460 421122 334524
rect 428089 334522 428155 334525
rect 428406 334522 428412 334524
rect 428089 334520 428412 334522
rect 428089 334464 428094 334520
rect 428150 334464 428412 334520
rect 428089 334462 428412 334464
rect 428089 334459 428155 334462
rect 428406 334460 428412 334462
rect 428476 334460 428482 334524
rect 447225 334250 447291 334253
rect 447225 334248 450156 334250
rect 447225 334192 447230 334248
rect 447286 334192 450156 334248
rect 447225 334190 450156 334192
rect 447225 334187 447291 334190
rect 513281 334114 513347 334117
rect 509956 334112 513347 334114
rect 509956 334056 513286 334112
rect 513342 334056 513347 334112
rect 509956 334054 513347 334056
rect 513281 334051 513347 334054
rect 447317 333570 447383 333573
rect 447317 333568 450156 333570
rect 447317 333512 447322 333568
rect 447378 333512 450156 333568
rect 447317 333510 450156 333512
rect 447317 333507 447383 333510
rect 509742 333165 509802 333540
rect 509742 333160 509851 333165
rect 509742 333104 509790 333160
rect 509846 333104 509851 333160
rect 509742 333102 509851 333104
rect 509785 333099 509851 333102
rect 510061 333026 510127 333029
rect 509956 333024 510127 333026
rect 509956 332968 510066 333024
rect 510122 332968 510127 333024
rect 509956 332966 510127 332968
rect 510061 332963 510127 332966
rect 432597 332890 432663 332893
rect 429916 332888 432663 332890
rect 429916 332832 432602 332888
rect 432658 332832 432663 332888
rect 429916 332830 432663 332832
rect 432597 332827 432663 332830
rect 447225 332890 447291 332893
rect 447225 332888 450156 332890
rect 447225 332832 447230 332888
rect 447286 332832 450156 332888
rect 447225 332830 450156 332832
rect 447225 332827 447291 332830
rect 511022 332482 511028 332484
rect -960 332196 480 332436
rect 509956 332422 511028 332482
rect 511022 332420 511028 332422
rect 511092 332420 511098 332484
rect 447501 332210 447567 332213
rect 447501 332208 450156 332210
rect 447501 332152 447506 332208
rect 447562 332152 450156 332208
rect 447501 332150 450156 332152
rect 447501 332147 447567 332150
rect 513281 331938 513347 331941
rect 509956 331936 513347 331938
rect 509956 331880 513286 331936
rect 513342 331880 513347 331936
rect 509956 331878 513347 331880
rect 513281 331875 513347 331878
rect 447225 331530 447291 331533
rect 447225 331528 450156 331530
rect 447225 331472 447230 331528
rect 447286 331472 450156 331528
rect 447225 331470 450156 331472
rect 447225 331467 447291 331470
rect 514150 331394 514156 331396
rect 509956 331334 514156 331394
rect 514150 331332 514156 331334
rect 514220 331332 514226 331396
rect 447317 330850 447383 330853
rect 512729 330850 512795 330853
rect 447317 330848 450156 330850
rect 447317 330792 447322 330848
rect 447378 330792 450156 330848
rect 447317 330790 450156 330792
rect 509956 330848 512795 330850
rect 509956 330792 512734 330848
rect 512790 330792 512795 330848
rect 509956 330790 512795 330792
rect 447317 330787 447383 330790
rect 512729 330787 512795 330790
rect 514702 330306 514708 330308
rect 509956 330246 514708 330306
rect 514702 330244 514708 330246
rect 514772 330244 514778 330308
rect 447225 330170 447291 330173
rect 447225 330168 450156 330170
rect 447225 330112 447230 330168
rect 447286 330112 450156 330168
rect 447225 330110 450156 330112
rect 447225 330107 447291 330110
rect 514886 329762 514892 329764
rect 509956 329702 514892 329762
rect 514886 329700 514892 329702
rect 514956 329700 514962 329764
rect 447225 329490 447291 329493
rect 447225 329488 450156 329490
rect 447225 329432 447230 329488
rect 447286 329432 450156 329488
rect 447225 329430 450156 329432
rect 447225 329427 447291 329430
rect 432781 329218 432847 329221
rect 510153 329218 510219 329221
rect 429916 329216 432847 329218
rect 429916 329160 432786 329216
rect 432842 329160 432847 329216
rect 429916 329158 432847 329160
rect 509956 329216 510219 329218
rect 509956 329160 510158 329216
rect 510214 329160 510219 329216
rect 509956 329158 510219 329160
rect 432781 329155 432847 329158
rect 510153 329155 510219 329158
rect 447225 328810 447291 328813
rect 448278 328810 448284 328812
rect 447225 328808 448284 328810
rect 447225 328752 447230 328808
rect 447286 328752 448284 328808
rect 447225 328750 448284 328752
rect 447225 328747 447291 328750
rect 448278 328748 448284 328750
rect 448348 328810 448354 328812
rect 448348 328750 450156 328810
rect 448348 328748 448354 328750
rect 515070 328674 515076 328676
rect 509956 328614 515076 328674
rect 515070 328612 515076 328614
rect 515140 328612 515146 328676
rect 447225 328130 447291 328133
rect 448094 328130 448100 328132
rect 447225 328128 448100 328130
rect 447225 328072 447230 328128
rect 447286 328072 448100 328128
rect 447225 328070 448100 328072
rect 447225 328067 447291 328070
rect 448094 328068 448100 328070
rect 448164 328130 448170 328132
rect 510245 328130 510311 328133
rect 448164 328070 450156 328130
rect 509956 328128 510311 328130
rect 509956 328072 510250 328128
rect 510306 328072 510311 328128
rect 509956 328070 510311 328072
rect 448164 328068 448170 328070
rect 510245 328067 510311 328070
rect 510838 327586 510844 327588
rect 509956 327526 510844 327586
rect 510838 327524 510844 327526
rect 510908 327524 510914 327588
rect 447317 327450 447383 327453
rect 447317 327448 450156 327450
rect 447317 327392 447322 327448
rect 447378 327392 450156 327448
rect 447317 327390 450156 327392
rect 447317 327387 447383 327390
rect 516174 327042 516180 327044
rect 509956 326982 516180 327042
rect 516174 326980 516180 326982
rect 516244 326980 516250 327044
rect 447225 326770 447291 326773
rect 448237 326770 448303 326773
rect 447225 326768 450156 326770
rect 447225 326712 447230 326768
rect 447286 326712 448242 326768
rect 448298 326712 450156 326768
rect 447225 326710 450156 326712
rect 447225 326707 447291 326710
rect 448237 326707 448303 326710
rect 362217 326498 362283 326501
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 359812 326438 362283 326440
rect 362217 326435 362283 326438
rect 509742 326093 509802 326468
rect 447317 326090 447383 326093
rect 447317 326088 450156 326090
rect 447317 326032 447322 326088
rect 447378 326032 450156 326088
rect 447317 326030 450156 326032
rect 509693 326088 509802 326093
rect 509693 326032 509698 326088
rect 509754 326032 509802 326088
rect 509693 326030 509802 326032
rect 447317 326027 447383 326030
rect 509693 326027 509759 326030
rect 514334 325954 514340 325956
rect 509956 325894 514340 325954
rect 514334 325892 514340 325894
rect 514404 325892 514410 325956
rect 432689 325546 432755 325549
rect 429916 325544 432755 325546
rect 429916 325488 432694 325544
rect 432750 325488 432755 325544
rect 429916 325486 432755 325488
rect 432689 325483 432755 325486
rect 448145 325410 448211 325413
rect 448421 325410 448487 325413
rect 512729 325410 512795 325413
rect 448145 325408 450156 325410
rect 448145 325352 448150 325408
rect 448206 325352 448426 325408
rect 448482 325352 450156 325408
rect 448145 325350 450156 325352
rect 509956 325408 512795 325410
rect 509956 325352 512734 325408
rect 512790 325352 512795 325408
rect 509956 325350 512795 325352
rect 448145 325347 448211 325350
rect 448421 325347 448487 325350
rect 512729 325347 512795 325350
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 517830 324866 517836 324868
rect 509956 324806 517836 324866
rect 517830 324804 517836 324806
rect 517900 324804 517906 324868
rect 447961 324730 448027 324733
rect 447961 324728 450156 324730
rect 447961 324672 447966 324728
rect 448022 324672 450156 324728
rect 447961 324670 450156 324672
rect 447961 324667 448027 324670
rect 511206 324322 511212 324324
rect 509956 324262 511212 324322
rect 511206 324260 511212 324262
rect 511276 324260 511282 324324
rect 449249 324186 449315 324189
rect 449249 324184 450738 324186
rect 449249 324128 449254 324184
rect 449310 324128 450738 324184
rect 449249 324126 450738 324128
rect 449249 324123 449315 324126
rect 450678 322965 450738 324126
rect 510470 323778 510476 323780
rect 509956 323718 510476 323778
rect 510470 323716 510476 323718
rect 510540 323716 510546 323780
rect 510286 323234 510292 323236
rect 509956 323174 510292 323234
rect 510286 323172 510292 323174
rect 510356 323172 510362 323236
rect 450678 322960 450787 322965
rect 450678 322904 450726 322960
rect 450782 322904 450787 322960
rect 450678 322902 450787 322904
rect 450721 322899 450787 322902
rect 506974 322900 506980 322964
rect 507044 322962 507050 322964
rect 510153 322962 510219 322965
rect 507044 322902 509066 322962
rect 507044 322900 507050 322902
rect 509006 322826 509066 322902
rect 509190 322960 510219 322962
rect 509190 322904 510158 322960
rect 510214 322904 510219 322960
rect 509190 322902 510219 322904
rect 509190 322826 509250 322902
rect 510153 322899 510219 322902
rect 509006 322766 509250 322826
rect 507301 322690 507367 322693
rect 510838 322690 510844 322692
rect 507301 322688 510844 322690
rect 507301 322632 507306 322688
rect 507362 322632 510844 322688
rect 507301 322630 510844 322632
rect 507301 322627 507367 322630
rect 510838 322628 510844 322630
rect 510908 322628 510914 322692
rect 507117 322554 507183 322557
rect 511022 322554 511028 322556
rect 507117 322552 511028 322554
rect 507117 322496 507122 322552
rect 507178 322496 511028 322552
rect 507117 322494 511028 322496
rect 507117 322491 507183 322494
rect 511022 322492 511028 322494
rect 511092 322492 511098 322556
rect 509182 322356 509188 322420
rect 509252 322418 509258 322420
rect 510286 322418 510292 322420
rect 509252 322358 510292 322418
rect 509252 322356 509258 322358
rect 510286 322356 510292 322358
rect 510356 322356 510362 322420
rect 432965 321874 433031 321877
rect 429916 321872 433031 321874
rect 429916 321816 432970 321872
rect 433026 321816 433031 321872
rect 429916 321814 433031 321816
rect 432965 321811 433031 321814
rect 446254 321812 446260 321876
rect 446324 321874 446330 321876
rect 460289 321874 460355 321877
rect 446324 321872 460355 321874
rect 446324 321816 460294 321872
rect 460350 321816 460355 321872
rect 446324 321814 460355 321816
rect 446324 321812 446330 321814
rect 460289 321811 460355 321814
rect 443494 321676 443500 321740
rect 443564 321738 443570 321740
rect 481541 321738 481607 321741
rect 443564 321736 481607 321738
rect 443564 321680 481546 321736
rect 481602 321680 481607 321736
rect 443564 321678 481607 321680
rect 443564 321676 443570 321678
rect 481541 321675 481607 321678
rect 442717 321602 442783 321605
rect 481817 321602 481883 321605
rect 442717 321600 481883 321602
rect 442717 321544 442722 321600
rect 442778 321544 481822 321600
rect 481878 321544 481883 321600
rect 442717 321542 481883 321544
rect 442717 321539 442783 321542
rect 481817 321539 481883 321542
rect 458633 321466 458699 321469
rect 559414 321466 559420 321468
rect 458633 321464 559420 321466
rect 458633 321408 458638 321464
rect 458694 321408 559420 321464
rect 458633 321406 559420 321408
rect 458633 321403 458699 321406
rect 559414 321404 559420 321406
rect 559484 321404 559490 321468
rect 449566 321268 449572 321332
rect 449636 321330 449642 321332
rect 480437 321330 480503 321333
rect 449636 321328 480503 321330
rect 449636 321272 480442 321328
rect 480498 321272 480503 321328
rect 449636 321270 480503 321272
rect 449636 321268 449642 321270
rect 480437 321267 480503 321270
rect 444230 321132 444236 321196
rect 444300 321194 444306 321196
rect 459737 321194 459803 321197
rect 444300 321192 459803 321194
rect 444300 321136 459742 321192
rect 459798 321136 459803 321192
rect 444300 321134 459803 321136
rect 444300 321132 444306 321134
rect 459737 321131 459803 321134
rect 444046 320996 444052 321060
rect 444116 321058 444122 321060
rect 460565 321058 460631 321061
rect 444116 321056 460631 321058
rect 444116 321000 460570 321056
rect 460626 321000 460631 321056
rect 444116 320998 460631 321000
rect 444116 320996 444122 320998
rect 460565 320995 460631 320998
rect 507669 320786 507735 320789
rect 514702 320786 514708 320788
rect 507669 320784 514708 320786
rect 507669 320728 507674 320784
rect 507730 320728 514708 320784
rect 507669 320726 514708 320728
rect 507669 320723 507735 320726
rect 514702 320724 514708 320726
rect 514772 320724 514778 320788
rect 446438 320044 446444 320108
rect 446508 320106 446514 320108
rect 471053 320106 471119 320109
rect 446508 320104 471119 320106
rect 446508 320048 471058 320104
rect 471114 320048 471119 320104
rect 446508 320046 471119 320048
rect 446508 320044 446514 320046
rect 471053 320043 471119 320046
rect 479609 320106 479675 320109
rect 529974 320106 529980 320108
rect 479609 320104 529980 320106
rect 479609 320048 479614 320104
rect 479670 320048 529980 320104
rect 479609 320046 529980 320048
rect 479609 320043 479675 320046
rect 529974 320044 529980 320046
rect 530044 320044 530050 320108
rect 450353 319970 450419 319973
rect 471605 319970 471671 319973
rect 450353 319968 471671 319970
rect 450353 319912 450358 319968
rect 450414 319912 471610 319968
rect 471666 319912 471671 319968
rect 450353 319910 471671 319912
rect 450353 319907 450419 319910
rect 471605 319907 471671 319910
rect 450486 319772 450492 319836
rect 450556 319834 450562 319836
rect 471329 319834 471395 319837
rect 450556 319832 471395 319834
rect 450556 319776 471334 319832
rect 471390 319776 471395 319832
rect 450556 319774 471395 319776
rect 450556 319772 450562 319774
rect 471329 319771 471395 319774
rect 497273 319426 497339 319429
rect 538806 319426 538812 319428
rect 497273 319424 538812 319426
rect -960 319290 480 319380
rect 497273 319368 497278 319424
rect 497334 319368 538812 319424
rect 497273 319366 538812 319368
rect 497273 319363 497339 319366
rect 538806 319364 538812 319366
rect 538876 319364 538882 319428
rect 3601 319290 3667 319293
rect -960 319288 3667 319290
rect -960 319232 3606 319288
rect 3662 319232 3667 319288
rect -960 319230 3667 319232
rect -960 319140 480 319230
rect 3601 319227 3667 319230
rect 432873 318202 432939 318205
rect 429916 318200 432939 318202
rect 429916 318144 432878 318200
rect 432934 318144 432939 318200
rect 429916 318142 432939 318144
rect 432873 318139 432939 318142
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 432137 314530 432203 314533
rect 429916 314528 432203 314530
rect 429916 314472 432142 314528
rect 432198 314472 432203 314528
rect 429916 314470 432203 314472
rect 432137 314467 432203 314470
rect 494973 313986 495039 313989
rect 542670 313986 542676 313988
rect 494973 313984 542676 313986
rect 494973 313928 494978 313984
rect 495034 313928 542676 313984
rect 494973 313926 542676 313928
rect 494973 313923 495039 313926
rect 542670 313924 542676 313926
rect 542740 313924 542746 313988
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 432597 310858 432663 310861
rect 429916 310856 432663 310858
rect 429916 310800 432602 310856
rect 432658 310800 432663 310856
rect 429916 310798 432663 310800
rect 432597 310795 432663 310798
rect 432229 307186 432295 307189
rect 429916 307184 432295 307186
rect 429916 307128 432234 307184
rect 432290 307128 432295 307184
rect 429916 307126 432295 307128
rect 432229 307123 432295 307126
rect 370497 306914 370563 306917
rect 514334 306914 514340 306916
rect 370497 306912 514340 306914
rect 370497 306856 370502 306912
rect 370558 306856 514340 306912
rect 370497 306854 514340 306856
rect 370497 306851 370563 306854
rect 514334 306852 514340 306854
rect 514404 306852 514410 306916
rect 380341 306778 380407 306781
rect 514886 306778 514892 306780
rect 380341 306776 514892 306778
rect 380341 306720 380346 306776
rect 380402 306720 514892 306776
rect 380341 306718 514892 306720
rect 380341 306715 380407 306718
rect 514886 306716 514892 306718
rect 514956 306716 514962 306780
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 376017 306234 376083 306237
rect 484485 306234 484551 306237
rect 376017 306232 484551 306234
rect 376017 306176 376022 306232
rect 376078 306176 484490 306232
rect 484546 306176 484551 306232
rect 376017 306174 484551 306176
rect 376017 306171 376083 306174
rect 484485 306171 484551 306174
rect 381813 306098 381879 306101
rect 510470 306098 510476 306100
rect 381813 306096 510476 306098
rect 381813 306040 381818 306096
rect 381874 306040 510476 306096
rect 381813 306038 510476 306040
rect 381813 306035 381879 306038
rect 510470 306036 510476 306038
rect 510540 306036 510546 306100
rect 381629 305962 381695 305965
rect 511206 305962 511212 305964
rect 381629 305960 511212 305962
rect 381629 305904 381634 305960
rect 381690 305904 511212 305960
rect 381629 305902 511212 305904
rect 381629 305899 381695 305902
rect 511206 305900 511212 305902
rect 511276 305900 511282 305964
rect 363597 305826 363663 305829
rect 512637 305826 512703 305829
rect 363597 305824 512703 305826
rect 363597 305768 363602 305824
rect 363658 305768 512642 305824
rect 512698 305768 512703 305824
rect 363597 305766 512703 305768
rect 363597 305763 363663 305766
rect 512637 305763 512703 305766
rect 381486 305628 381492 305692
rect 381556 305690 381562 305692
rect 508998 305690 509004 305692
rect 381556 305630 509004 305690
rect 381556 305628 381562 305630
rect 508998 305628 509004 305630
rect 509068 305628 509074 305692
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 382181 303106 382247 303109
rect 509693 303106 509759 303109
rect 382181 303104 509759 303106
rect 382181 303048 382186 303104
rect 382242 303048 509698 303104
rect 509754 303048 509759 303104
rect 382181 303046 509759 303048
rect 382181 303043 382247 303046
rect 509693 303043 509759 303046
rect 381445 302970 381511 302973
rect 511165 302970 511231 302973
rect 381445 302968 511231 302970
rect 381445 302912 381450 302968
rect 381506 302912 511170 302968
rect 511226 302912 511231 302968
rect 381445 302910 511231 302912
rect 381445 302907 381511 302910
rect 511165 302907 511231 302910
rect 379237 302834 379303 302837
rect 515489 302834 515555 302837
rect 379237 302832 515555 302834
rect 379237 302776 379242 302832
rect 379298 302776 515494 302832
rect 515550 302776 515555 302832
rect 379237 302774 515555 302776
rect 379237 302771 379303 302774
rect 515489 302771 515555 302774
rect 383009 300250 383075 300253
rect 518341 300250 518407 300253
rect 383009 300248 518407 300250
rect 383009 300192 383014 300248
rect 383070 300192 518346 300248
rect 518402 300192 518407 300248
rect 383009 300190 518407 300192
rect 383009 300187 383075 300190
rect 518341 300187 518407 300190
rect 373533 300114 373599 300117
rect 510245 300114 510311 300117
rect 373533 300112 510311 300114
rect 373533 300056 373538 300112
rect 373594 300056 510250 300112
rect 510306 300056 510311 300112
rect 373533 300054 510311 300056
rect 373533 300051 373599 300054
rect 510245 300051 510311 300054
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 371969 297802 372035 297805
rect 516174 297802 516180 297804
rect 371969 297800 516180 297802
rect 371969 297744 371974 297800
rect 372030 297744 516180 297800
rect 371969 297742 516180 297744
rect 371969 297739 372035 297742
rect 516174 297740 516180 297742
rect 516244 297740 516250 297804
rect 362401 297666 362467 297669
rect 510654 297666 510660 297668
rect 362401 297664 510660 297666
rect 362401 297608 362406 297664
rect 362462 297608 510660 297664
rect 362401 297606 510660 297608
rect 362401 297603 362467 297606
rect 510654 297604 510660 297606
rect 510724 297604 510730 297668
rect 365161 297530 365227 297533
rect 514150 297530 514156 297532
rect 365161 297528 514156 297530
rect 365161 297472 365166 297528
rect 365222 297472 514156 297528
rect 365161 297470 514156 297472
rect 365161 297467 365227 297470
rect 514150 297468 514156 297470
rect 514220 297468 514226 297532
rect 365345 297394 365411 297397
rect 517830 297394 517836 297396
rect 365345 297392 517836 297394
rect 365345 297336 365350 297392
rect 365406 297336 517836 297392
rect 365345 297334 517836 297336
rect 365345 297331 365411 297334
rect 517830 297332 517836 297334
rect 517900 297332 517906 297396
rect 372153 294538 372219 294541
rect 515070 294538 515076 294540
rect 372153 294536 515076 294538
rect 372153 294480 372158 294536
rect 372214 294480 515076 294536
rect 372153 294478 515076 294480
rect 372153 294475 372219 294478
rect 515070 294476 515076 294478
rect 515140 294476 515146 294540
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 384757 289098 384823 289101
rect 506974 289098 506980 289100
rect 384757 289096 506980 289098
rect 384757 289040 384762 289096
rect 384818 289040 506980 289096
rect 384757 289038 506980 289040
rect 384757 289035 384823 289038
rect 506974 289036 506980 289038
rect 507044 289036 507050 289100
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 362585 271418 362651 271421
rect 359812 271416 362651 271418
rect 359812 271360 362590 271416
rect 362646 271360 362651 271416
rect 359812 271358 362651 271360
rect 362585 271355 362651 271358
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 529289 261626 529355 261629
rect 529289 261624 529490 261626
rect 529289 261568 529294 261624
rect 529350 261568 529490 261624
rect 529289 261566 529490 261568
rect 529289 261563 529355 261566
rect 529430 261052 529490 261566
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 456793 248842 456859 248845
rect 456793 248840 460092 248842
rect 456793 248784 456798 248840
rect 456854 248784 460092 248840
rect 456793 248782 460092 248784
rect 456793 248779 456859 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 530117 243674 530183 243677
rect 529828 243672 530183 243674
rect 529828 243616 530122 243672
rect 530178 243616 530183 243672
rect 529828 243614 530183 243616
rect 530117 243611 530183 243614
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 457805 234970 457871 234973
rect 458081 234970 458147 234973
rect 457805 234968 460092 234970
rect 457805 234912 457810 234968
rect 457866 234912 458086 234968
rect 458142 234912 460092 234968
rect 457805 234910 460092 234912
rect 457805 234907 457871 234910
rect 458081 234907 458147 234910
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 459461 221098 459527 221101
rect 459461 221096 460092 221098
rect 459461 221040 459466 221096
rect 459522 221040 460092 221096
rect 459461 221038 460092 221040
rect 459461 221035 459527 221038
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 361665 216338 361731 216341
rect 359812 216336 361731 216338
rect 359812 216280 361670 216336
rect 361726 216280 361731 216336
rect 359812 216278 361731 216280
rect 361665 216275 361731 216278
rect -960 214978 480 215068
rect 3877 214978 3943 214981
rect -960 214976 3943 214978
rect -960 214920 3882 214976
rect 3938 214920 3943 214976
rect -960 214918 3943 214920
rect -960 214828 480 214918
rect 3877 214915 3943 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 456793 207226 456859 207229
rect 456793 207224 460092 207226
rect 456793 207168 456798 207224
rect 456854 207168 460092 207224
rect 456793 207166 460092 207168
rect 456793 207163 456859 207166
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 361757 194306 361823 194309
rect 359812 194304 361823 194306
rect 359812 194248 361762 194304
rect 361818 194248 361823 194304
rect 359812 194246 361823 194248
rect 361757 194243 361823 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 4061 188866 4127 188869
rect -960 188864 4127 188866
rect -960 188808 4066 188864
rect 4122 188808 4127 188864
rect -960 188806 4127 188808
rect -960 188716 480 188806
rect 4061 188803 4127 188806
rect 361757 183290 361823 183293
rect 359812 183288 361823 183290
rect 359812 183232 361762 183288
rect 361818 183232 361823 183288
rect 359812 183230 361823 183232
rect 361757 183227 361823 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361757 172274 361823 172277
rect 359812 172272 361823 172274
rect 359812 172216 361762 172272
rect 361818 172216 361823 172272
rect 359812 172214 361823 172216
rect 361757 172211 361823 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 421046 162692 421052 162756
rect 421116 162754 421122 162756
rect 421557 162754 421623 162757
rect 421116 162752 421623 162754
rect 421116 162696 421562 162752
rect 421618 162696 421623 162752
rect 421116 162694 421623 162696
rect 421116 162692 421122 162694
rect 421557 162691 421623 162694
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 451549 158266 451615 158269
rect 449788 158264 451615 158266
rect 449788 158208 451554 158264
rect 451610 158208 451615 158264
rect 449788 158206 451615 158208
rect 451549 158203 451615 158206
rect 451733 156906 451799 156909
rect 449788 156904 451799 156906
rect 449788 156848 451738 156904
rect 451794 156848 451799 156904
rect 449788 156846 451799 156848
rect 451733 156843 451799 156846
rect 452561 155546 452627 155549
rect 449788 155544 452627 155546
rect 449788 155488 452566 155544
rect 452622 155488 452627 155544
rect 449788 155486 452627 155488
rect 452561 155483 452627 155486
rect 451733 154186 451799 154189
rect 449788 154184 451799 154186
rect 449788 154128 451738 154184
rect 451794 154128 451799 154184
rect 449788 154126 451799 154128
rect 451733 154123 451799 154126
rect 451641 152826 451707 152829
rect 449788 152824 451707 152826
rect 449788 152768 451646 152824
rect 451702 152768 451707 152824
rect 449788 152766 451707 152768
rect 451641 152763 451707 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 451457 151466 451523 151469
rect 449788 151464 451523 151466
rect 449788 151408 451462 151464
rect 451518 151408 451523 151464
rect 449788 151406 451523 151408
rect 451457 151403 451523 151406
rect 362585 150242 362651 150245
rect 359812 150240 362651 150242
rect 359812 150184 362590 150240
rect 362646 150184 362651 150240
rect 359812 150182 362651 150184
rect 362585 150179 362651 150182
rect 452377 150106 452443 150109
rect 449788 150104 452443 150106
rect 449788 150048 452382 150104
rect 452438 150048 452443 150104
rect 449788 150046 452443 150048
rect 452377 150043 452443 150046
rect -960 149834 480 149924
rect 3233 149834 3299 149837
rect -960 149832 3299 149834
rect -960 149776 3238 149832
rect 3294 149776 3299 149832
rect -960 149774 3299 149776
rect -960 149684 480 149774
rect 3233 149771 3299 149774
rect 452193 148746 452259 148749
rect 449788 148744 452259 148746
rect 449788 148688 452198 148744
rect 452254 148688 452259 148744
rect 449788 148686 452259 148688
rect 452193 148683 452259 148686
rect 452561 147386 452627 147389
rect 449788 147384 452627 147386
rect 449788 147328 452566 147384
rect 452622 147328 452627 147384
rect 449788 147326 452627 147328
rect 452561 147323 452627 147326
rect 452561 146026 452627 146029
rect 449788 146024 452627 146026
rect 449788 145968 452566 146024
rect 452622 145968 452627 146024
rect 449788 145966 452627 145968
rect 452561 145963 452627 145966
rect 452561 144666 452627 144669
rect 449788 144664 452627 144666
rect 449788 144608 452566 144664
rect 452622 144608 452627 144664
rect 449788 144606 452627 144608
rect 452561 144603 452627 144606
rect 452561 143306 452627 143309
rect 449788 143304 452627 143306
rect 449788 143248 452566 143304
rect 452622 143248 452627 143304
rect 449788 143246 452627 143248
rect 452561 143243 452627 143246
rect 452561 141946 452627 141949
rect 449788 141944 452627 141946
rect 449788 141888 452566 141944
rect 452622 141888 452627 141944
rect 449788 141886 452627 141888
rect 452561 141883 452627 141886
rect 452561 140586 452627 140589
rect 449788 140584 452627 140586
rect 449788 140528 452566 140584
rect 452622 140528 452627 140584
rect 449788 140526 452627 140528
rect 452561 140523 452627 140526
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 451549 139226 451615 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 359812 139166 361823 139168
rect 449788 139224 451615 139226
rect 449788 139168 451554 139224
rect 451610 139168 451615 139224
rect 583520 139212 584960 139302
rect 449788 139166 451615 139168
rect 361757 139163 361823 139166
rect 451549 139163 451615 139166
rect 538949 138002 539015 138005
rect 538949 138000 539610 138002
rect 538949 137944 538954 138000
rect 539010 137944 539610 138000
rect 538949 137942 539610 137944
rect 538949 137939 539015 137942
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 539550 137428 539610 137942
rect -960 136778 480 136868
rect 3366 136778 3372 136780
rect -960 136718 3372 136778
rect -960 136628 480 136718
rect 3366 136716 3372 136718
rect 3436 136716 3442 136780
rect 539358 136716 539364 136780
rect 539428 136778 539434 136780
rect 542997 136778 543063 136781
rect 539428 136776 543063 136778
rect 539428 136720 543002 136776
rect 543058 136720 543063 136776
rect 539428 136718 543063 136720
rect 539428 136716 539434 136718
rect 542997 136715 543063 136718
rect 452561 136506 452627 136509
rect 449788 136504 452627 136506
rect 449788 136448 452566 136504
rect 452622 136448 452627 136504
rect 449788 136446 452627 136448
rect 452561 136443 452627 136446
rect 539317 135690 539383 135693
rect 539317 135688 539426 135690
rect 539317 135632 539322 135688
rect 539378 135632 539426 135688
rect 539317 135627 539426 135632
rect 539366 135388 539426 135627
rect 452561 135146 452627 135149
rect 449788 135144 452627 135146
rect 449788 135088 452566 135144
rect 452622 135088 452627 135144
rect 449788 135086 452627 135088
rect 452561 135083 452627 135086
rect 452561 133786 452627 133789
rect 449788 133784 452627 133786
rect 449788 133728 452566 133784
rect 452622 133728 452627 133784
rect 449788 133726 452627 133728
rect 452561 133723 452627 133726
rect 541525 133378 541591 133381
rect 539948 133376 541591 133378
rect 539948 133320 541530 133376
rect 541586 133320 541591 133376
rect 539948 133318 541591 133320
rect 541525 133315 541591 133318
rect 452193 132426 452259 132429
rect 449788 132424 452259 132426
rect 449788 132368 452198 132424
rect 452254 132368 452259 132424
rect 449788 132366 452259 132368
rect 452193 132363 452259 132366
rect 543181 131338 543247 131341
rect 539948 131336 543247 131338
rect 539948 131280 543186 131336
rect 543242 131280 543247 131336
rect 539948 131278 543247 131280
rect 543181 131275 543247 131278
rect 452377 131066 452443 131069
rect 449788 131064 452443 131066
rect 449788 131008 452382 131064
rect 452438 131008 452443 131064
rect 449788 131006 452443 131008
rect 452377 131003 452443 131006
rect 452285 129706 452351 129709
rect 449788 129704 452351 129706
rect 449788 129648 452290 129704
rect 452346 129648 452351 129704
rect 449788 129646 452351 129648
rect 452285 129643 452351 129646
rect 540329 129298 540395 129301
rect 539948 129296 540395 129298
rect 539948 129240 540334 129296
rect 540390 129240 540395 129296
rect 539948 129238 540395 129240
rect 540329 129235 540395 129238
rect 452009 128346 452075 128349
rect 449788 128344 452075 128346
rect 449788 128288 452014 128344
rect 452070 128288 452075 128344
rect 449788 128286 452075 128288
rect 452009 128283 452075 128286
rect 361757 128210 361823 128213
rect 359812 128208 361823 128210
rect 359812 128152 361762 128208
rect 361818 128152 361823 128208
rect 359812 128150 361823 128152
rect 361757 128147 361823 128150
rect 542905 127258 542971 127261
rect 539948 127256 542971 127258
rect 539948 127200 542910 127256
rect 542966 127200 542971 127256
rect 539948 127198 542971 127200
rect 542905 127195 542971 127198
rect 452377 126986 452443 126989
rect 449788 126984 452443 126986
rect 449788 126928 452382 126984
rect 452438 126928 452443 126984
rect 449788 126926 452443 126928
rect 452377 126923 452443 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 452101 125626 452167 125629
rect 449788 125624 452167 125626
rect 449788 125568 452106 125624
rect 452162 125568 452167 125624
rect 449788 125566 452167 125568
rect 452101 125563 452167 125566
rect 540237 125218 540303 125221
rect 539948 125216 540303 125218
rect 539948 125160 540242 125216
rect 540298 125160 540303 125216
rect 539948 125158 540303 125160
rect 540237 125155 540303 125158
rect 451917 124266 451983 124269
rect 449788 124264 451983 124266
rect 449788 124208 451922 124264
rect 451978 124208 451983 124264
rect 449788 124206 451983 124208
rect 451917 124203 451983 124206
rect -960 123572 480 123812
rect 543089 123178 543155 123181
rect 539948 123176 543155 123178
rect 539948 123120 543094 123176
rect 543150 123120 543155 123176
rect 539948 123118 543155 123120
rect 543089 123115 543155 123118
rect 451917 122906 451983 122909
rect 449788 122904 451983 122906
rect 449788 122848 451922 122904
rect 451978 122848 451983 122904
rect 449788 122846 451983 122848
rect 451917 122843 451983 122846
rect 451917 121546 451983 121549
rect 449788 121544 451983 121546
rect 449788 121488 451922 121544
rect 451978 121488 451983 121544
rect 449788 121486 451983 121488
rect 451917 121483 451983 121486
rect 542629 121138 542695 121141
rect 539948 121136 542695 121138
rect 539948 121080 542634 121136
rect 542690 121080 542695 121136
rect 539948 121078 542695 121080
rect 542629 121075 542695 121078
rect 539685 119642 539751 119645
rect 539685 119640 539794 119642
rect 539685 119584 539690 119640
rect 539746 119584 539794 119640
rect 539685 119579 539794 119584
rect 539734 119068 539794 119579
rect 361757 117194 361823 117197
rect 359812 117192 361823 117194
rect 359812 117136 361762 117192
rect 361818 117136 361823 117192
rect 359812 117134 361823 117136
rect 361757 117131 361823 117134
rect 540145 117058 540211 117061
rect 539948 117056 540211 117058
rect 539948 117000 540150 117056
rect 540206 117000 540211 117056
rect 539948 116998 540211 117000
rect 540145 116995 540211 116998
rect 541157 115018 541223 115021
rect 539948 115016 541223 115018
rect 539948 114960 541162 115016
rect 541218 114960 541223 115016
rect 539948 114958 541223 114960
rect 541157 114955 541223 114958
rect 539918 112845 539978 112948
rect 539918 112840 540027 112845
rect 539918 112784 539966 112840
rect 540022 112784 540027 112840
rect 539918 112782 540027 112784
rect 539961 112779 540027 112782
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 540053 111482 540119 111485
rect 539918 111480 540119 111482
rect 539918 111424 540058 111480
rect 540114 111424 540119 111480
rect 539918 111422 540119 111424
rect 539918 110908 539978 111422
rect 540053 111419 540119 111422
rect -960 110666 480 110756
rect 3550 110666 3556 110668
rect -960 110606 3556 110666
rect -960 110516 480 110606
rect 3550 110604 3556 110606
rect 3620 110604 3626 110668
rect 541065 108898 541131 108901
rect 539948 108896 541131 108898
rect 539948 108840 541070 108896
rect 541126 108840 541131 108896
rect 539948 108838 541131 108840
rect 541065 108835 541131 108838
rect 541433 106858 541499 106861
rect 539948 106856 541499 106858
rect 539948 106800 541438 106856
rect 541494 106800 541499 106856
rect 539948 106798 541499 106800
rect 541433 106795 541499 106798
rect 361757 106178 361823 106181
rect 359812 106176 361823 106178
rect 359812 106120 361762 106176
rect 361818 106120 361823 106176
rect 359812 106118 361823 106120
rect 361757 106115 361823 106118
rect 541249 104818 541315 104821
rect 539948 104816 541315 104818
rect 539948 104760 541254 104816
rect 541310 104760 541315 104816
rect 539948 104758 541315 104760
rect 541249 104755 541315 104758
rect 541341 102778 541407 102781
rect 539948 102776 541407 102778
rect 539948 102720 541346 102776
rect 541402 102720 541407 102776
rect 539948 102718 541407 102720
rect 541341 102715 541407 102718
rect 542997 100738 543063 100741
rect 539948 100736 543063 100738
rect 539948 100680 543002 100736
rect 543058 100680 543063 100736
rect 539948 100678 543063 100680
rect 542997 100675 543063 100678
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 539777 99242 539843 99245
rect 539734 99240 539843 99242
rect 539734 99184 539782 99240
rect 539838 99184 539843 99240
rect 539734 99179 539843 99184
rect 539734 98668 539794 99179
rect -960 97610 480 97700
rect 3693 97610 3759 97613
rect -960 97608 3759 97610
rect -960 97552 3698 97608
rect 3754 97552 3759 97608
rect -960 97550 3759 97552
rect -960 97460 480 97550
rect 3693 97547 3759 97550
rect 539593 97202 539659 97205
rect 539550 97200 539659 97202
rect 539550 97144 539598 97200
rect 539654 97144 539659 97200
rect 539550 97139 539659 97144
rect 539550 96628 539610 97139
rect 361757 95162 361823 95165
rect 359812 95160 361823 95162
rect 359812 95104 361762 95160
rect 361818 95104 361823 95160
rect 359812 95102 361823 95104
rect 361757 95099 361823 95102
rect 542813 94618 542879 94621
rect 539948 94616 542879 94618
rect 539948 94560 542818 94616
rect 542874 94560 542879 94616
rect 539948 94558 542879 94560
rect 542813 94555 542879 94558
rect 542537 92578 542603 92581
rect 539948 92576 542603 92578
rect 539948 92520 542542 92576
rect 542598 92520 542603 92576
rect 539948 92518 542603 92520
rect 542537 92515 542603 92518
rect 542445 90538 542511 90541
rect 539948 90536 542511 90538
rect 539948 90480 542450 90536
rect 542506 90480 542511 90536
rect 539948 90478 542511 90480
rect 542445 90475 542511 90478
rect 543273 88498 543339 88501
rect 539948 88496 543339 88498
rect 539948 88440 543278 88496
rect 543334 88440 543339 88496
rect 539948 88438 543339 88440
rect 543273 88435 543339 88438
rect 542721 86458 542787 86461
rect 539948 86456 542787 86458
rect 539948 86400 542726 86456
rect 542782 86400 542787 86456
rect 539948 86398 542787 86400
rect 542721 86395 542787 86398
rect 578877 86186 578943 86189
rect 583520 86186 584960 86276
rect 578877 86184 584960 86186
rect 578877 86128 578882 86184
rect 578938 86128 584960 86184
rect 578877 86126 584960 86128
rect 578877 86123 578943 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 542670 84418 542676 84420
rect 539948 84358 542676 84418
rect 542670 84356 542676 84358
rect 542740 84356 542746 84420
rect 361665 84146 361731 84149
rect 359812 84144 361731 84146
rect 359812 84088 361670 84144
rect 361726 84088 361731 84144
rect 359812 84086 361731 84088
rect 361665 84083 361731 84086
rect 540973 82378 541039 82381
rect 539948 82376 541039 82378
rect 539948 82320 540978 82376
rect 541034 82320 541039 82376
rect 539948 82318 541039 82320
rect 540973 82315 541039 82318
rect 20897 73674 20963 73677
rect 21449 73674 21515 73677
rect 20897 73672 21515 73674
rect 20897 73616 20902 73672
rect 20958 73616 21454 73672
rect 21510 73616 21515 73672
rect 20897 73614 21515 73616
rect 20897 73611 20963 73614
rect 21449 73611 21515 73614
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3141 71634 3207 71637
rect -960 71632 3207 71634
rect -960 71576 3146 71632
rect 3202 71576 3207 71632
rect -960 71574 3207 71576
rect -960 71484 480 71574
rect 3141 71571 3207 71574
rect 462313 67554 462379 67557
rect 462957 67554 463023 67557
rect 460828 67552 463023 67554
rect 460828 67496 462318 67552
rect 462374 67496 462962 67552
rect 463018 67496 463023 67552
rect 460828 67494 463023 67496
rect 462313 67491 462379 67494
rect 462957 67491 463023 67494
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3141 58578 3207 58581
rect -960 58576 3207 58578
rect -960 58520 3146 58576
rect 3202 58520 3207 58576
rect -960 58518 3207 58520
rect -960 58428 480 58518
rect 3141 58515 3207 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 18873 49602 18939 49605
rect 22318 49602 22324 49604
rect 18873 49600 22324 49602
rect 18873 49544 18878 49600
rect 18934 49544 22324 49600
rect 18873 49542 22324 49544
rect 18873 49539 18939 49542
rect 22318 49540 22324 49542
rect 22388 49540 22394 49604
rect 15193 48922 15259 48925
rect 22134 48922 22140 48924
rect 15193 48920 22140 48922
rect 15193 48864 15198 48920
rect 15254 48864 22140 48920
rect 15193 48862 22140 48864
rect 15193 48859 15259 48862
rect 22134 48860 22140 48862
rect 22204 48860 22210 48924
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3366 46956 3372 47020
rect 3436 47018 3442 47020
rect 384941 47018 385007 47021
rect 3436 47016 385007 47018
rect 3436 46960 384946 47016
rect 385002 46960 385007 47016
rect 3436 46958 385007 46960
rect 3436 46956 3442 46958
rect 384941 46955 385007 46958
rect 3550 46820 3556 46884
rect 3620 46882 3626 46884
rect 385953 46882 386019 46885
rect 3620 46880 386019 46882
rect 3620 46824 385958 46880
rect 386014 46824 386019 46880
rect 3620 46822 386019 46824
rect 3620 46820 3626 46822
rect 385953 46819 386019 46822
rect 20069 46746 20135 46749
rect 384573 46746 384639 46749
rect 20069 46744 384639 46746
rect 20069 46688 20074 46744
rect 20130 46688 384578 46744
rect 384634 46688 384639 46744
rect 20069 46686 384639 46688
rect 20069 46683 20135 46686
rect 384573 46683 384639 46686
rect 22134 46548 22140 46612
rect 22204 46610 22210 46612
rect 359825 46610 359891 46613
rect 22204 46608 359891 46610
rect 22204 46552 359830 46608
rect 359886 46552 359891 46608
rect 22204 46550 359891 46552
rect 22204 46548 22210 46550
rect 359825 46547 359891 46550
rect 22318 46412 22324 46476
rect 22388 46474 22394 46476
rect 359641 46474 359707 46477
rect 22388 46472 359707 46474
rect 22388 46416 359646 46472
rect 359702 46416 359707 46472
rect 22388 46414 359707 46416
rect 22388 46412 22394 46414
rect 359641 46411 359707 46414
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 6913 44842 6979 44845
rect 382181 44842 382247 44845
rect 6913 44840 382247 44842
rect 6913 44784 6918 44840
rect 6974 44784 382186 44840
rect 382242 44784 382247 44840
rect 6913 44782 382247 44784
rect 6913 44779 6979 44782
rect 382181 44779 382247 44782
rect 536833 41034 536899 41037
rect 536833 41032 540132 41034
rect 536833 40976 536838 41032
rect 536894 40976 540132 41032
rect 536833 40974 540132 40976
rect 536833 40971 536899 40974
rect 539869 33690 539935 33693
rect 539869 33688 540132 33690
rect 539869 33632 539874 33688
rect 539930 33632 540132 33688
rect 539869 33630 540132 33632
rect 539869 33627 539935 33630
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 5257 4042 5323 4045
rect 362217 4042 362283 4045
rect 5257 4040 362283 4042
rect 5257 3984 5262 4040
rect 5318 3984 362222 4040
rect 362278 3984 362283 4040
rect 5257 3982 362283 3984
rect 5257 3979 5323 3982
rect 362217 3979 362283 3982
rect 13537 3906 13603 3909
rect 372153 3906 372219 3909
rect 13537 3904 372219 3906
rect 13537 3848 13542 3904
rect 13598 3848 372158 3904
rect 372214 3848 372219 3904
rect 13537 3846 372219 3848
rect 13537 3843 13603 3846
rect 372153 3843 372219 3846
rect 8753 3770 8819 3773
rect 371969 3770 372035 3773
rect 8753 3768 372035 3770
rect 8753 3712 8758 3768
rect 8814 3712 371974 3768
rect 372030 3712 372035 3768
rect 8753 3710 372035 3712
rect 8753 3707 8819 3710
rect 371969 3707 372035 3710
rect 6453 3634 6519 3637
rect 370497 3634 370563 3637
rect 6453 3632 370563 3634
rect 6453 3576 6458 3632
rect 6514 3576 370502 3632
rect 370558 3576 370563 3632
rect 6453 3574 370563 3576
rect 6453 3571 6519 3574
rect 370497 3571 370563 3574
rect 1669 3498 1735 3501
rect 381813 3498 381879 3501
rect 1669 3496 381879 3498
rect 1669 3440 1674 3496
rect 1730 3440 381818 3496
rect 381874 3440 381879 3496
rect 1669 3438 381879 3440
rect 1669 3435 1735 3438
rect 381813 3435 381879 3438
rect 565 3362 631 3365
rect 381486 3362 381492 3364
rect 565 3360 381492 3362
rect 565 3304 570 3360
rect 626 3304 381492 3360
rect 565 3302 381492 3304
rect 565 3299 631 3302
rect 381486 3300 381492 3302
rect 381556 3300 381562 3364
<< via3 >>
rect 449572 700572 449636 700636
rect 444236 700436 444300 700500
rect 446260 700300 446324 700364
rect 455092 700300 455156 700364
rect 529980 699756 530044 699820
rect 559420 699756 559484 699820
rect 450492 687788 450556 687852
rect 446444 685068 446508 685132
rect 3556 683300 3620 683364
rect 3740 683164 3804 683228
rect 3372 682756 3436 682820
rect 3740 671196 3804 671260
rect 453252 669836 453316 669900
rect 459508 667932 459572 667996
rect 458036 665212 458100 665276
rect 459140 630668 459204 630732
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 474780 599660 474844 599724
rect 476436 599524 476500 599588
rect 474964 598164 475028 598228
rect 478828 595444 478892 595508
rect 459508 562940 459572 563004
rect 474412 541588 474476 541652
rect 458036 523636 458100 523700
rect 474596 522276 474660 522340
rect 472020 518060 472084 518124
rect 448284 516156 448348 516220
rect 448100 514176 448164 514180
rect 448100 514120 448114 514176
rect 448114 514120 448164 514176
rect 448100 514116 448164 514120
rect 448100 500244 448164 500308
rect 481772 496904 481836 496908
rect 481772 496848 481822 496904
rect 481822 496848 481836 496904
rect 481772 496844 481836 496848
rect 483060 496844 483124 496908
rect 448284 496028 448348 496092
rect 487108 453868 487172 453932
rect 455092 422860 455156 422924
rect 443500 421908 443564 421972
rect 444052 421772 444116 421836
rect 459140 410484 459204 410548
rect 483060 389812 483124 389876
rect 472020 388996 472084 389060
rect 474412 389056 474476 389060
rect 474412 389000 474426 389056
rect 474426 389000 474476 389056
rect 474412 388996 474476 389000
rect 474964 388996 475028 389060
rect 476436 388996 476500 389060
rect 478828 388996 478892 389060
rect 474596 388860 474660 388924
rect 474780 388860 474844 388924
rect 453252 387092 453316 387156
rect 481772 386956 481836 387020
rect 487108 385596 487172 385660
rect 510660 334596 510724 334660
rect 421052 334460 421116 334524
rect 428412 334460 428476 334524
rect 511028 332420 511092 332484
rect 514156 331332 514220 331396
rect 514708 330244 514772 330308
rect 514892 329700 514956 329764
rect 448284 328748 448348 328812
rect 515076 328612 515140 328676
rect 448100 328068 448164 328132
rect 510844 327524 510908 327588
rect 516180 326980 516244 327044
rect 514340 325892 514404 325956
rect 517836 324804 517900 324868
rect 511212 324260 511276 324324
rect 510476 323716 510540 323780
rect 510292 323172 510356 323236
rect 506980 322900 507044 322964
rect 510844 322628 510908 322692
rect 511028 322492 511092 322556
rect 509188 322356 509252 322420
rect 510292 322356 510356 322420
rect 446260 321812 446324 321876
rect 443500 321676 443564 321740
rect 559420 321404 559484 321468
rect 449572 321268 449636 321332
rect 444236 321132 444300 321196
rect 444052 320996 444116 321060
rect 514708 320724 514772 320788
rect 446444 320044 446508 320108
rect 529980 320044 530044 320108
rect 450492 319772 450556 319836
rect 538812 319364 538876 319428
rect 542676 313924 542740 313988
rect 514340 306852 514404 306916
rect 514892 306716 514956 306780
rect 510476 306036 510540 306100
rect 511212 305900 511276 305964
rect 381492 305628 381556 305692
rect 509004 305628 509068 305692
rect 516180 297740 516244 297804
rect 510660 297604 510724 297668
rect 514156 297468 514220 297532
rect 517836 297332 517900 297396
rect 515076 294476 515140 294540
rect 506980 289036 507044 289100
rect 421052 162692 421116 162756
rect 428412 162692 428476 162756
rect 3372 136716 3436 136780
rect 539364 136716 539428 136780
rect 3556 110604 3620 110668
rect 542676 84356 542740 84420
rect 22324 49540 22388 49604
rect 22140 48860 22204 48924
rect 3372 46956 3436 47020
rect 3556 46820 3620 46884
rect 22140 46548 22204 46612
rect 22324 46412 22388 46476
rect 381492 3300 381556 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3555 683364 3621 683365
rect 3555 683300 3556 683364
rect 3620 683300 3621 683364
rect 3555 683299 3621 683300
rect 3371 682820 3437 682821
rect 3371 682756 3372 682820
rect 3436 682756 3437 682820
rect 3371 682755 3437 682756
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682755
rect 3558 619173 3618 683299
rect 3739 683228 3805 683229
rect 3739 683164 3740 683228
rect 3804 683164 3805 683228
rect 3739 683163 3805 683164
rect 3742 671261 3802 683163
rect 3739 671260 3805 671261
rect 3739 671196 3740 671260
rect 3804 671196 3805 671260
rect 3739 671195 3805 671196
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3371 136780 3437 136781
rect 3371 136716 3372 136780
rect 3436 136716 3437 136780
rect 3371 136715 3437 136716
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 47021 3434 136715
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3555 110668 3621 110669
rect 3555 110604 3556 110668
rect 3620 110604 3621 110668
rect 3555 110603 3621 110604
rect 3371 47020 3437 47021
rect 3371 46956 3372 47020
rect 3436 46956 3437 47020
rect 3371 46955 3437 46956
rect 3558 46885 3618 110603
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3555 46884 3621 46885
rect 3555 46820 3556 46884
rect 3620 46820 3621 46884
rect 3555 46819 3621 46820
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674393 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674393 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674393 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674393 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 674393 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674393 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674393 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674393 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674393 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 674393 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674393 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674393 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674393 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674393 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 674393 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674393 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674393 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674393 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674393 157574 698058
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 674393 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674393 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674393 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674393 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 674393 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674393 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674393 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674393 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674393 229574 698058
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 674393 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674393 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674393 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674393 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674393 265574 698058
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 674393 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674393 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674393 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674393 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674393 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674393 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674393 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674393 337574 698058
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 674393 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22323 49604 22389 49605
rect 22323 49540 22324 49604
rect 22388 49540 22389 49604
rect 22323 49539 22389 49540
rect 22139 48924 22205 48925
rect 22139 48860 22140 48924
rect 22204 48860 22205 48924
rect 22139 48859 22205 48860
rect 22142 46613 22202 48859
rect 22139 46612 22205 46613
rect 22139 46548 22140 46612
rect 22204 46548 22205 46612
rect 22139 46547 22205 46548
rect 22326 46477 22386 49539
rect 22323 46476 22389 46477
rect 22323 46412 22324 46476
rect 22388 46412 22389 46476
rect 22323 46411 22389 46412
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 49367
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 49367
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 49367
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 49367
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 49367
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 49367
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 49367
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 49367
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 49367
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 49367
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 49367
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 49367
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 49367
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 49367
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 49367
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 49367
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 49367
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 49367
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 49367
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 49367
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 49367
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 49367
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 49367
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 49367
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 49367
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 49367
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 49367
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 49367
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 49367
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 49367
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 49367
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 49367
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 49367
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 49367
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 49367
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 49367
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 49367
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 49367
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 49367
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 49367
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 49367
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 49367
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 49367
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 49367
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 49367
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 49367
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 49367
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 49367
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 49367
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 49367
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 49367
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 49367
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 49367
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 49367
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 49367
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 49367
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 49367
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 49367
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 49367
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 49367
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 49367
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 49367
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 49367
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 49367
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 49367
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 49367
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 49367
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 49367
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 49367
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 381491 305692 381557 305693
rect 381491 305628 381492 305692
rect 381556 305628 381557 305692
rect 381491 305627 381557 305628
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 381494 3365 381554 305627
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 92137 388454 100938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 92137 398414 110898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 92137 402134 114618
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 104460 405854 118338
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 92137 409574 122058
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444235 700500 444301 700501
rect 444235 700436 444236 700500
rect 444300 700436 444301 700500
rect 444235 700435 444301 700436
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 157249 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421051 334524 421117 334525
rect 421051 334460 421052 334524
rect 421116 334460 421117 334524
rect 421051 334459 421117 334460
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 157249 420734 169218
rect 421054 162757 421114 334459
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 428411 334524 428477 334525
rect 428411 334460 428412 334524
rect 428476 334460 428477 334524
rect 428411 334459 428477 334460
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421051 162756 421117 162757
rect 421051 162692 421052 162756
rect 421116 162692 421117 162756
rect 421051 162691 421117 162692
rect 423834 157249 424454 172938
rect 428414 162757 428474 334459
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 157249 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 157249 438134 186618
rect 441234 406894 441854 422599
rect 443499 421972 443565 421973
rect 443499 421908 443500 421972
rect 443564 421908 443565 421972
rect 443499 421907 443565 421908
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 443502 321741 443562 421907
rect 444051 421836 444117 421837
rect 444051 421772 444052 421836
rect 444116 421772 444117 421836
rect 444051 421771 444117 421772
rect 443499 321740 443565 321741
rect 443499 321676 443500 321740
rect 443564 321676 443565 321740
rect 443499 321675 443565 321676
rect 444054 321061 444114 421771
rect 444238 321197 444298 700435
rect 444954 698614 445574 707162
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 446259 700364 446325 700365
rect 446259 700300 446260 700364
rect 446324 700300 446325 700364
rect 446259 700299 446325 700300
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 321196 444301 321197
rect 444235 321132 444236 321196
rect 444300 321132 444301 321196
rect 444235 321131 444301 321132
rect 444051 321060 444117 321061
rect 444051 320996 444052 321060
rect 444116 320996 444117 321060
rect 444051 320995 444117 320996
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 157249 441854 190338
rect 444954 302614 445574 338058
rect 446262 321877 446322 700299
rect 446443 685132 446509 685133
rect 446443 685068 446444 685132
rect 446508 685068 446509 685132
rect 446443 685067 446509 685068
rect 446259 321876 446325 321877
rect 446259 321812 446260 321876
rect 446324 321812 446325 321876
rect 446259 321811 446325 321812
rect 446446 320109 446506 685067
rect 448674 666334 449294 708122
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 449571 700636 449637 700637
rect 449571 700572 449572 700636
rect 449636 700572 449637 700636
rect 449571 700571 449637 700572
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448283 516220 448349 516221
rect 448283 516156 448284 516220
rect 448348 516156 448349 516220
rect 448283 516155 448349 516156
rect 448099 514180 448165 514181
rect 448099 514116 448100 514180
rect 448164 514116 448165 514180
rect 448099 514115 448165 514116
rect 448102 500309 448162 514115
rect 448099 500308 448165 500309
rect 448099 500244 448100 500308
rect 448164 500244 448165 500308
rect 448099 500243 448165 500244
rect 448102 328133 448162 500243
rect 448286 496093 448346 516155
rect 448283 496092 448349 496093
rect 448283 496028 448284 496092
rect 448348 496028 448349 496092
rect 448283 496027 448349 496028
rect 448286 328813 448346 496027
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448283 328812 448349 328813
rect 448283 328748 448284 328812
rect 448348 328748 448349 328812
rect 448283 328747 448349 328748
rect 448099 328132 448165 328133
rect 448099 328068 448100 328132
rect 448164 328068 448165 328132
rect 448099 328067 448165 328068
rect 446443 320108 446509 320109
rect 446443 320044 446444 320108
rect 446508 320044 446509 320108
rect 446443 320043 446509 320044
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 159644 445574 194058
rect 448674 306334 449294 341778
rect 449574 321333 449634 700571
rect 450491 687852 450557 687853
rect 450491 687788 450492 687852
rect 450556 687788 450557 687852
rect 450491 687787 450557 687788
rect 449571 321332 449637 321333
rect 449571 321268 449572 321332
rect 449636 321268 449637 321332
rect 449571 321267 449637 321268
rect 450494 319837 450554 687787
rect 452394 670054 453014 709082
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 455091 700364 455157 700365
rect 455091 700300 455092 700364
rect 455156 700300 455157 700364
rect 455091 700299 455157 700300
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 453251 669900 453317 669901
rect 453251 669836 453252 669900
rect 453316 669836 453317 669900
rect 453251 669835 453317 669836
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 453254 387157 453314 669835
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 455094 422925 455154 700299
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 669073 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 669073 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 669073 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 669073 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 669073 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 669073 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 669073 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 669073 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 669073 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 669073 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 669073 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 669073 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 459507 667996 459573 667997
rect 459507 667932 459508 667996
rect 459572 667932 459573 667996
rect 459507 667931 459573 667932
rect 458035 665276 458101 665277
rect 458035 665212 458036 665276
rect 458100 665212 458101 665276
rect 458035 665211 458101 665212
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 458038 523701 458098 665211
rect 459139 630732 459205 630733
rect 459139 630668 459140 630732
rect 459204 630668 459205 630732
rect 459139 630667 459205 630668
rect 458035 523700 458101 523701
rect 458035 523636 458036 523700
rect 458100 523636 458101 523700
rect 458035 523635 458101 523636
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 455091 422924 455157 422925
rect 455091 422860 455092 422924
rect 455156 422860 455157 422924
rect 455091 422859 455157 422860
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 453251 387156 453317 387157
rect 453251 387092 453252 387156
rect 453316 387092 453317 387156
rect 453251 387091 453317 387092
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 385774 456734 421218
rect 459142 410549 459202 630667
rect 459510 563005 459570 667931
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 459834 569494 460454 601103
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459507 563004 459573 563005
rect 459507 562940 459508 563004
rect 459572 562940 459573 563004
rect 459507 562939 459573 562940
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 517884 460454 532938
rect 469794 579454 470414 601103
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 473514 583174 474134 601103
rect 474779 599724 474845 599725
rect 474779 599660 474780 599724
rect 474844 599660 474845 599724
rect 474779 599659 474845 599660
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 472019 518124 472085 518125
rect 472019 518060 472020 518124
rect 472084 518060 472085 518124
rect 472019 518059 472085 518060
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459139 410548 459205 410549
rect 459139 410484 459140 410548
rect 459204 410484 459205 410548
rect 459139 410483 459205 410484
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450491 319836 450557 319837
rect 450491 319772 450492 319836
rect 450556 319772 450557 319836
rect 450491 319771 450557 319772
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 92137 413294 125778
rect 416394 94054 417014 127767
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 92137 417014 93498
rect 420114 97774 420734 127767
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 92137 420734 97218
rect 423834 101494 424454 127767
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 92137 424454 100938
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 92137 449294 125778
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 92137 453014 93498
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 92137 456734 97218
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 389061 472082 518059
rect 473514 511174 474134 546618
rect 474411 541652 474477 541653
rect 474411 541588 474412 541652
rect 474476 541588 474477 541652
rect 474411 541587 474477 541588
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 541587
rect 474595 522340 474661 522341
rect 474595 522276 474596 522340
rect 474660 522276 474661 522340
rect 474595 522275 474661 522276
rect 472019 389060 472085 389061
rect 472019 388996 472020 389060
rect 472084 388996 472085 389060
rect 472019 388995 472085 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 474598 388925 474658 522275
rect 474782 388925 474842 599659
rect 476435 599588 476501 599589
rect 476435 599524 476436 599588
rect 476500 599524 476501 599588
rect 476435 599523 476501 599524
rect 474963 598228 475029 598229
rect 474963 598164 474964 598228
rect 475028 598164 475029 598228
rect 474963 598163 475029 598164
rect 474966 389061 475026 598163
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 476438 389061 476498 599523
rect 477234 586894 477854 601103
rect 478827 595508 478893 595509
rect 478827 595444 478828 595508
rect 478892 595444 478893 595508
rect 478827 595443 478893 595444
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 474963 389060 475029 389061
rect 474963 388996 474964 389060
rect 475028 388996 475029 389060
rect 474963 388995 475029 388996
rect 476435 389060 476501 389061
rect 476435 388996 476436 389060
rect 476500 388996 476501 389060
rect 476435 388995 476501 388996
rect 474595 388924 474661 388925
rect 474595 388860 474596 388924
rect 474660 388860 474661 388924
rect 474595 388859 474661 388860
rect 474779 388924 474845 388925
rect 474779 388860 474780 388924
rect 474844 388860 474845 388924
rect 474779 388859 474845 388860
rect 477234 385225 477854 406338
rect 478830 389061 478890 595443
rect 480954 590614 481574 601103
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 601103
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 601103
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 601103
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 481771 496908 481837 496909
rect 481771 496844 481772 496908
rect 481836 496844 481837 496908
rect 481771 496843 481837 496844
rect 483059 496908 483125 496909
rect 483059 496844 483060 496908
rect 483124 496844 483125 496908
rect 483059 496843 483125 496844
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 481774 387021 481834 496843
rect 483062 389877 483122 496843
rect 484674 486334 485294 500068
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 488394 490054 489014 500068
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 487107 453932 487173 453933
rect 487107 453868 487108 453932
rect 487172 453868 487173 453932
rect 487107 453867 487173 453868
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 483059 389876 483125 389877
rect 483059 389812 483060 389876
rect 483124 389812 483125 389876
rect 483059 389811 483125 389812
rect 481771 387020 481837 387021
rect 481771 386956 481772 387020
rect 481836 386956 481837 387020
rect 481771 386955 481837 386956
rect 484674 385580 485294 413778
rect 487110 385661 487170 453867
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 487107 385660 487173 385661
rect 487107 385596 487108 385660
rect 487172 385596 487173 385660
rect 487107 385595 487173 385596
rect 492114 385225 492734 421218
rect 495834 569494 496454 601103
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 385225 496454 388938
rect 505794 579454 506414 601103
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 385225 506414 398898
rect 509514 583174 510134 601103
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 509514 331174 510134 366618
rect 513234 586894 513854 601103
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 510659 334660 510725 334661
rect 510659 334596 510660 334660
rect 510724 334596 510725 334660
rect 510659 334595 510725 334596
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 506979 322964 507045 322965
rect 506979 322900 506980 322964
rect 507044 322900 507045 322964
rect 506979 322899 507045 322900
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 469794 291454 470414 321879
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 248401 470414 254898
rect 473514 295174 474134 321879
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 248401 474134 258618
rect 477234 298894 477854 321879
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 248401 477854 262338
rect 480954 302614 481574 321879
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 480954 248401 481574 266058
rect 484674 306334 485294 321879
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 248401 485294 269778
rect 488394 310054 489014 321879
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 248401 489014 273498
rect 492114 313774 492734 321879
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 248401 492734 277218
rect 495834 317494 496454 321879
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 495834 248401 496454 280938
rect 505794 291454 506414 321879
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 506982 289101 507042 322899
rect 509006 322630 509250 322690
rect 509006 305693 509066 322630
rect 509190 322421 509250 322630
rect 509187 322420 509253 322421
rect 509187 322356 509188 322420
rect 509252 322356 509253 322420
rect 509187 322355 509253 322356
rect 509003 305692 509069 305693
rect 509003 305628 509004 305692
rect 509068 305628 509069 305692
rect 509003 305627 509069 305628
rect 509514 295174 510134 330618
rect 510475 323780 510541 323781
rect 510475 323716 510476 323780
rect 510540 323716 510541 323780
rect 510475 323715 510541 323716
rect 510291 323236 510357 323237
rect 510291 323172 510292 323236
rect 510356 323172 510357 323236
rect 510291 323171 510357 323172
rect 510294 322421 510354 323171
rect 510291 322420 510357 322421
rect 510291 322356 510292 322420
rect 510356 322356 510357 322420
rect 510291 322355 510357 322356
rect 510478 306101 510538 323715
rect 510475 306100 510541 306101
rect 510475 306036 510476 306100
rect 510540 306036 510541 306100
rect 510475 306035 510541 306036
rect 510662 297669 510722 334595
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 511027 332484 511093 332485
rect 511027 332420 511028 332484
rect 511092 332420 511093 332484
rect 511027 332419 511093 332420
rect 510843 327588 510909 327589
rect 510843 327524 510844 327588
rect 510908 327524 510909 327588
rect 510843 327523 510909 327524
rect 510846 322693 510906 327523
rect 510843 322692 510909 322693
rect 510843 322628 510844 322692
rect 510908 322628 510909 322692
rect 510843 322627 510909 322628
rect 511030 322557 511090 332419
rect 511211 324324 511277 324325
rect 511211 324260 511212 324324
rect 511276 324260 511277 324324
rect 511211 324259 511277 324260
rect 511027 322556 511093 322557
rect 511027 322492 511028 322556
rect 511092 322492 511093 322556
rect 511027 322491 511093 322492
rect 511214 305965 511274 324259
rect 511211 305964 511277 305965
rect 511211 305900 511212 305964
rect 511276 305900 511277 305964
rect 511211 305899 511277 305900
rect 513234 298894 513854 334338
rect 516954 590614 517574 601103
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 514155 331396 514221 331397
rect 514155 331332 514156 331396
rect 514220 331332 514221 331396
rect 514155 331331 514221 331332
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 510659 297668 510725 297669
rect 510659 297604 510660 297668
rect 510724 297604 510725 297668
rect 510659 297603 510725 297604
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 506979 289100 507045 289101
rect 506979 289036 506980 289100
rect 507044 289036 507045 289100
rect 506979 289035 507045 289036
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 248401 506414 254898
rect 509514 259174 510134 294618
rect 513234 262894 513854 298338
rect 514158 297533 514218 331331
rect 514707 330308 514773 330309
rect 514707 330244 514708 330308
rect 514772 330244 514773 330308
rect 514707 330243 514773 330244
rect 514339 325956 514405 325957
rect 514339 325892 514340 325956
rect 514404 325892 514405 325956
rect 514339 325891 514405 325892
rect 514342 306917 514402 325891
rect 514710 320789 514770 330243
rect 514891 329764 514957 329765
rect 514891 329700 514892 329764
rect 514956 329700 514957 329764
rect 514891 329699 514957 329700
rect 514707 320788 514773 320789
rect 514707 320724 514708 320788
rect 514772 320724 514773 320788
rect 514707 320723 514773 320724
rect 514339 306916 514405 306917
rect 514339 306852 514340 306916
rect 514404 306852 514405 306916
rect 514339 306851 514405 306852
rect 514894 306781 514954 329699
rect 515075 328676 515141 328677
rect 515075 328612 515076 328676
rect 515140 328612 515141 328676
rect 515075 328611 515141 328612
rect 514891 306780 514957 306781
rect 514891 306716 514892 306780
rect 514956 306716 514957 306780
rect 514891 306715 514957 306716
rect 514155 297532 514221 297533
rect 514155 297468 514156 297532
rect 514220 297468 514221 297532
rect 514155 297467 514221 297468
rect 515078 294541 515138 328611
rect 516179 327044 516245 327045
rect 516179 326980 516180 327044
rect 516244 326980 516245 327044
rect 516179 326979 516245 326980
rect 516182 297805 516242 326979
rect 516954 302614 517574 338058
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 517835 324868 517901 324869
rect 517835 324804 517836 324868
rect 517900 324804 517901 324868
rect 517835 324803 517901 324804
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516179 297804 516245 297805
rect 516179 297740 516180 297804
rect 516244 297740 516245 297804
rect 516179 297739 516245 297740
rect 515075 294540 515141 294541
rect 515075 294476 515076 294540
rect 515140 294476 515141 294540
rect 515075 294475 515141 294476
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 248401 510134 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 513234 248401 513854 262338
rect 516954 266614 517574 302058
rect 517838 297397 517898 324803
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 517835 297396 517901 297397
rect 517835 297332 517836 297396
rect 517900 297332 517901 297396
rect 517835 297331 517901 297332
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 248401 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 248401 521294 269778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 529979 699820 530045 699821
rect 529979 699756 529980 699820
rect 530044 699756 530045 699820
rect 529979 699755 530045 699756
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 248401 525014 273498
rect 528114 421774 528734 457218
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 529982 320109 530042 699755
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 529979 320108 530045 320109
rect 529979 320044 529980 320108
rect 530044 320044 530045 320108
rect 529979 320043 530045 320044
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 528114 248401 528734 277218
rect 531834 317494 532454 352938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 538811 319428 538877 319429
rect 538811 319364 538812 319428
rect 538876 319364 538877 319428
rect 538811 319363 538877 319364
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 405568 79174 405888 79206
rect 405568 78938 405610 79174
rect 405846 78938 405888 79174
rect 405568 78854 405888 78938
rect 405568 78618 405610 78854
rect 405846 78618 405888 78854
rect 405568 78586 405888 78618
rect 436288 79174 436608 79206
rect 436288 78938 436330 79174
rect 436566 78938 436608 79174
rect 436288 78854 436608 78938
rect 436288 78618 436330 78854
rect 436566 78618 436608 78854
rect 436288 78586 436608 78618
rect 390208 75454 390528 75486
rect 390208 75218 390250 75454
rect 390486 75218 390528 75454
rect 390208 75134 390528 75218
rect 390208 74898 390250 75134
rect 390486 74898 390528 75134
rect 390208 74866 390528 74898
rect 420928 75454 421248 75486
rect 420928 75218 420970 75454
rect 421206 75218 421248 75454
rect 420928 75134 421248 75218
rect 420928 74898 420970 75134
rect 421206 74898 421248 75134
rect 420928 74866 421248 74898
rect 451648 75454 451968 75486
rect 451648 75218 451690 75454
rect 451926 75218 451968 75454
rect 451648 75134 451968 75218
rect 451648 74898 451690 75134
rect 451926 74898 451968 75134
rect 451648 74866 451968 74898
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 405568 43174 405888 43206
rect 405568 42938 405610 43174
rect 405846 42938 405888 43174
rect 405568 42854 405888 42938
rect 405568 42618 405610 42854
rect 405846 42618 405888 42854
rect 405568 42586 405888 42618
rect 436288 43174 436608 43206
rect 436288 42938 436330 43174
rect 436566 42938 436608 43174
rect 436288 42854 436608 42938
rect 436288 42618 436330 42854
rect 436566 42618 436608 42854
rect 436288 42586 436608 42618
rect 390208 39454 390528 39486
rect 390208 39218 390250 39454
rect 390486 39218 390528 39454
rect 390208 39134 390528 39218
rect 390208 38898 390250 39134
rect 390486 38898 390528 39134
rect 390208 38866 390528 38898
rect 420928 39454 421248 39486
rect 420928 39218 420970 39454
rect 421206 39218 421248 39454
rect 420928 39134 421248 39218
rect 420928 38898 420970 39134
rect 421206 38898 421248 39134
rect 420928 38866 421248 38898
rect 451648 39454 451968 39486
rect 451648 39218 451690 39454
rect 451926 39218 451968 39454
rect 451648 39134 451968 39218
rect 451648 38898 451690 39134
rect 451926 38898 451968 39134
rect 451648 38866 451968 38898
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 381491 3364 381557 3365
rect 381491 3300 381492 3364
rect 381556 3300 381557 3364
rect 381491 3299 381557 3300
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 32599
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 3454 398414 32599
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 32599
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 30068
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 32599
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 32599
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 32599
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 32599
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 32599
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 32599
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 32599
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 32599
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 32599
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 32599
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 32599
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 32599
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 207495
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 207495
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 207495
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 207495
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 207495
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 488394 202054 489014 207495
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 166054 489014 201498
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 139281 489014 165498
rect 492114 205774 492734 207495
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 139281 492734 169218
rect 505794 183454 506414 207495
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139281 506414 146898
rect 509514 187174 510134 207495
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139281 510134 150618
rect 513234 190894 513854 207495
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139281 513854 154338
rect 516954 194614 517574 207495
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139281 517574 158058
rect 520674 198334 521294 207495
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139281 521294 161778
rect 524394 202054 525014 207495
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139281 525014 165498
rect 528114 205774 528734 207495
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 139281 528734 169218
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139281 532454 172938
rect 538814 151830 538874 319363
rect 541794 291454 542414 326898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 542675 313988 542741 313989
rect 542675 313924 542676 313988
rect 542740 313924 542741 313988
rect 542675 313923 542741 313924
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 538814 151770 539426 151830
rect 539366 136781 539426 151770
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 539363 136780 539429 136781
rect 539363 136716 539364 136780
rect 539428 136716 539429 136780
rect 539363 136715 539429 136716
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 58054 489014 82599
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 82599
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 82599
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 82599
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 82599
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 82599
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 82599
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 82599
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 82599
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 82599
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 82599
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 542678 84421 542738 313923
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 542675 84420 542741 84421
rect 542675 84356 542676 84420
rect 542740 84356 542741 84420
rect 542675 84355 542741 84356
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 559419 699820 559485 699821
rect 559419 699756 559420 699820
rect 559484 699756 559485 699820
rect 559419 699755 559485 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 559422 321469 559482 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 559419 321468 559485 321469
rect 559419 321404 559420 321468
rect 559484 321404 559485 321468
rect 559419 321403 559485 321404
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 405610 78938 405846 79174
rect 405610 78618 405846 78854
rect 436330 78938 436566 79174
rect 436330 78618 436566 78854
rect 390250 75218 390486 75454
rect 390250 74898 390486 75134
rect 420970 75218 421206 75454
rect 420970 74898 421206 75134
rect 451690 75218 451926 75454
rect 451690 74898 451926 75134
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 405610 42938 405846 43174
rect 405610 42618 405846 42854
rect 436330 42938 436566 43174
rect 436330 42618 436566 42854
rect 390250 39218 390486 39454
rect 390250 38898 390486 39134
rect 420970 39218 421206 39454
rect 420970 38898 421206 39134
rect 451690 39218 451926 39454
rect 451690 38898 451926 39134
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 479610 259174
rect 479846 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 479610 258854
rect 479846 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 494970 255454
rect 495206 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 494970 255134
rect 495206 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 405610 79174
rect 405846 78938 436330 79174
rect 436566 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 405610 78854
rect 405846 78618 436330 78854
rect 436566 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 390250 75454
rect 390486 75218 420970 75454
rect 421206 75218 451690 75454
rect 451926 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 390250 75134
rect 390486 74898 420970 75134
rect 421206 74898 451690 75134
rect 451926 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 405610 43174
rect 405846 42938 436330 43174
rect 436566 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 405610 42854
rect 405846 42618 436330 42854
rect 436566 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 390250 39454
rect 390486 39218 420970 39454
rect 421206 39218 451690 39454
rect 451926 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 390250 39134
rect 390486 38898 420970 39134
rect 421206 38898 451690 39134
rect 451926 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
use wrapped_vgatest  wrapped_vgatest
timestamp 0
transform 1 0 386000 0 1 30000
box 658 2128 75000 75000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 674393 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 674393 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 674393 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 674393 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 674393 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 674393 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 674393 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 674393 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 674393 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 32599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 92137 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 32599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 157249 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 207495 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 248401 470414 321879 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 669073 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 82599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139281 506414 207495 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 248401 506414 321879 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 385225 506414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 669073 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 674393 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 674393 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 674393 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 674393 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 674393 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 674393 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 674393 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 674393 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 674393 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 30068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 104460 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 32599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 157249 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 207495 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 248401 477854 321879 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 385225 477854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 669073 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 82599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139281 513854 207495 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 248401 513854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 669073 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 32599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 92137 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 32599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 92137 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 207495 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 248401 485294 321879 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 601103 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 82599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139281 521294 207495 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 248401 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 32599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 92137 420734 127767 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 157249 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 32599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 92137 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 139281 492734 207495 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 248401 492734 321879 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 385225 492734 601103 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 669073 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 139281 528734 207495 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 248401 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 32599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 92137 417014 127767 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 157249 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 32599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 92137 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 139281 489014 207495 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 248401 489014 321879 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 601103 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 669073 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139281 525014 207495 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 248401 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 674393 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 674393 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 674393 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 674393 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 674393 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 674393 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 674393 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 674393 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 32599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 92137 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 32599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 92137 424454 127767 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 157249 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 669073 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 248401 496454 321879 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 385225 496454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 669073 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139281 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 674393 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 674393 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 674393 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 674393 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 674393 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 674393 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 674393 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 674393 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 674393 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 32599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 92137 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 32599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 157249 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 207495 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 248401 474134 321879 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 669073 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 82599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139281 510134 207495 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 248401 510134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 669073 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 674393 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 674393 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 674393 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 674393 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 674393 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 674393 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 674393 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 32599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 92137 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 32599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 159644 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 207495 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 248401 481574 321879 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 669073 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 82599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139281 517574 207495 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 248401 517574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 669073 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 451808 75336 451808 75336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 521144 666216 521144 666216 0 vdda1
rlabel via4 456584 97656 456584 97656 0 vdda2
rlabel via4 452864 93936 452864 93936 0 vssa1
rlabel via4 460304 101376 460304 101376 0 vssa2
rlabel via4 436448 79056 436448 79056 0 vssd1
rlabel via4 481424 122496 481424 122496 0 vssd2
rlabel metal1 423062 447542 423062 447542 0 design_clk
rlabel metal2 411578 159868 411578 159868 0 dsi_all\[0\]
rlabel metal1 446660 331194 446660 331194 0 dsi_all\[10\]
rlabel metal1 445464 331262 445464 331262 0 dsi_all\[11\]
rlabel metal3 448830 332180 448830 332180 0 dsi_all\[12\]
rlabel metal2 447258 332741 447258 332741 0 dsi_all\[13\]
rlabel metal2 447350 333115 447350 333115 0 dsi_all\[14\]
rlabel metal2 447258 334101 447258 334101 0 dsi_all\[15\]
rlabel metal1 445556 334050 445556 334050 0 dsi_all\[16\]
rlabel metal1 444820 335478 444820 335478 0 dsi_all\[17\]
rlabel metal2 447258 335801 447258 335801 0 dsi_all\[18\]
rlabel metal2 447166 336855 447166 336855 0 dsi_all\[19\]
rlabel metal3 450156 503589 450156 503589 0 dsi_all\[1\]
rlabel metal1 445556 336838 445556 336838 0 dsi_all\[20\]
rlabel metal2 447166 338249 447166 338249 0 dsi_all\[21\]
rlabel metal2 385802 316030 385802 316030 0 dsi_all\[22\]
rlabel metal1 444820 339558 444820 339558 0 dsi_all\[23\]
rlabel metal2 447166 339915 447166 339915 0 dsi_all\[24\]
rlabel metal2 444130 338504 444130 338504 0 dsi_all\[25\]
rlabel metal2 447166 341309 447166 341309 0 dsi_all\[26\]
rlabel metal3 449658 342380 449658 342380 0 dsi_all\[27\]
rlabel metal3 450156 505395 450156 505395 0 dsi_all\[2\]
rlabel metal2 447350 326553 447350 326553 0 dsi_all\[3\]
rlabel metal2 425040 159994 425040 159994 0 dsi_all\[4\]
rlabel metal2 428184 159868 428184 159868 0 dsi_all\[5\]
rlabel metal2 431496 159868 431496 159868 0 dsi_all\[6\]
rlabel metal3 448692 328780 448692 328780 0 dsi_all\[7\]
rlabel metal2 447258 329273 447258 329273 0 dsi_all\[8\]
rlabel metal3 448692 330140 448692 330140 0 dsi_all\[9\]
rlabel metal2 451950 121839 451950 121839 0 dso_6502\[0\]
rlabel via2 452594 135133 452594 135133 0 dso_6502\[10\]
rlabel via2 452594 136493 452594 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel metal2 451582 139281 451582 139281 0 dso_6502\[13\]
rlabel metal2 452594 140607 452594 140607 0 dso_6502\[14\]
rlabel via2 452594 141933 452594 141933 0 dso_6502\[15\]
rlabel metal1 473386 274006 473386 274006 0 dso_6502\[16\]
rlabel metal1 474858 275366 474858 275366 0 dso_6502\[17\]
rlabel via2 452594 146013 452594 146013 0 dso_6502\[18\]
rlabel metal1 474306 276794 474306 276794 0 dso_6502\[19\]
rlabel metal2 451950 123131 451950 123131 0 dso_6502\[1\]
rlabel metal3 451022 148716 451022 148716 0 dso_6502\[20\]
rlabel metal3 451114 150076 451114 150076 0 dso_6502\[21\]
rlabel metal1 473386 272510 473386 272510 0 dso_6502\[22\]
rlabel metal2 451674 152983 451674 152983 0 dso_6502\[23\]
rlabel metal2 451766 154343 451766 154343 0 dso_6502\[24\]
rlabel via2 452594 155533 452594 155533 0 dso_6502\[25\]
rlabel metal2 451766 157097 451766 157097 0 dso_6502\[26\]
rlabel metal1 469936 311270 469936 311270 0 dso_6502\[2\]
rlabel metal3 450976 125596 450976 125596 0 dso_6502\[3\]
rlabel via2 452410 126939 452410 126939 0 dso_6502\[4\]
rlabel metal1 470442 309842 470442 309842 0 dso_6502\[5\]
rlabel metal1 470626 271150 470626 271150 0 dso_6502\[6\]
rlabel metal1 471316 308414 471316 308414 0 dso_6502\[7\]
rlabel via2 452226 132413 452226 132413 0 dso_6502\[8\]
rlabel via2 452594 133773 452594 133773 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 387862 505310 387862 0 dso_LCD\[2\]
rlabel metal2 506046 388576 506046 388576 0 dso_LCD\[3\]
rlabel metal2 506637 385900 506637 385900 0 dso_LCD\[4\]
rlabel metal2 507281 385900 507281 385900 0 dso_LCD\[5\]
rlabel metal2 508109 385900 508109 385900 0 dso_LCD\[6\]
rlabel metal2 508799 385900 508799 385900 0 dso_LCD\[7\]
rlabel metal3 540492 82348 540492 82348 0 dso_as1802\[0\]
rlabel metal3 540676 102748 540676 102748 0 dso_as1802\[10\]
rlabel metal3 540630 104788 540630 104788 0 dso_as1802\[11\]
rlabel metal3 540722 106828 540722 106828 0 dso_as1802\[12\]
rlabel metal3 540538 108868 540538 108868 0 dso_as1802\[13\]
rlabel metal3 539948 111195 539948 111195 0 dso_as1802\[14\]
rlabel metal3 539948 112865 539948 112865 0 dso_as1802\[15\]
rlabel metal3 540584 114988 540584 114988 0 dso_as1802\[16\]
rlabel metal3 540078 117028 540078 117028 0 dso_as1802\[17\]
rlabel via2 539741 119612 539741 119612 0 dso_as1802\[18\]
rlabel metal3 541320 121108 541320 121108 0 dso_as1802\[19\]
rlabel metal3 541343 84388 541343 84388 0 dso_as1802\[1\]
rlabel metal1 541006 138550 541006 138550 0 dso_as1802\[20\]
rlabel metal2 499974 297019 499974 297019 0 dso_as1802\[21\]
rlabel metal1 500250 319090 500250 319090 0 dso_as1802\[22\]
rlabel metal2 501170 316686 501170 316686 0 dso_as1802\[23\]
rlabel metal2 501446 320902 501446 320902 0 dso_as1802\[24\]
rlabel metal3 540768 133348 540768 133348 0 dso_as1802\[25\]
rlabel via2 539373 135660 539373 135660 0 dso_as1802\[26\]
rlabel metal3 541366 86428 541366 86428 0 dso_as1802\[2\]
rlabel metal3 541642 88468 541642 88468 0 dso_as1802\[3\]
rlabel metal3 541228 90508 541228 90508 0 dso_as1802\[4\]
rlabel metal3 541274 92548 541274 92548 0 dso_as1802\[5\]
rlabel metal3 541412 94588 541412 94588 0 dso_as1802\[6\]
rlabel via2 539603 97172 539603 97172 0 dso_as1802\[7\]
rlabel via2 539787 99212 539787 99212 0 dso_as1802\[8\]
rlabel metal3 541504 100708 541504 100708 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal1 465152 541654 465152 541654 0 dso_as2650\[10\]
rlabel metal2 471217 385900 471217 385900 0 dso_as2650\[11\]
rlabel metal2 472091 385900 472091 385900 0 dso_as2650\[12\]
rlabel metal2 472926 387471 472926 387471 0 dso_as2650\[13\]
rlabel metal3 459747 635460 459747 635460 0 dso_as2650\[14\]
rlabel metal3 459701 637908 459701 637908 0 dso_as2650\[15\]
rlabel metal3 459517 640356 459517 640356 0 dso_as2650\[16\]
rlabel metal3 459563 643212 459563 643212 0 dso_as2650\[17\]
rlabel metal2 461610 494598 461610 494598 0 dso_as2650\[18\]
rlabel metal2 477342 387471 477342 387471 0 dso_as2650\[19\]
rlabel metal2 463903 385900 463903 385900 0 dso_as2650\[1\]
rlabel metal2 469890 494258 469890 494258 0 dso_as2650\[20\]
rlabel metal2 468510 493510 468510 493510 0 dso_as2650\[21\]
rlabel metal3 459640 655724 459640 655724 0 dso_as2650\[22\]
rlabel metal2 480286 387318 480286 387318 0 dso_as2650\[23\]
rlabel metal2 481022 387182 481022 387182 0 dso_as2650\[24\]
rlabel metal2 481758 387216 481758 387216 0 dso_as2650\[25\]
rlabel metal2 482494 387284 482494 387284 0 dso_as2650\[26\]
rlabel metal2 464593 385900 464593 385900 0 dso_as2650\[2\]
rlabel metal2 465329 385900 465329 385900 0 dso_as2650\[3\]
rlabel metal2 466065 385900 466065 385900 0 dso_as2650\[4\]
rlabel metal2 466801 385900 466801 385900 0 dso_as2650\[5\]
rlabel metal2 467583 385900 467583 385900 0 dso_as2650\[6\]
rlabel metal2 468510 387284 468510 387284 0 dso_as2650\[7\]
rlabel metal2 469246 387522 469246 387522 0 dso_as2650\[8\]
rlabel metal2 469982 387046 469982 387046 0 dso_as2650\[9\]
rlabel metal2 444038 367778 444038 367778 0 dso_as512512512\[0\]
rlabel metal2 447258 372045 447258 372045 0 dso_as512512512\[10\]
rlabel metal2 447166 372419 447166 372419 0 dso_as512512512\[11\]
rlabel metal2 447258 373439 447258 373439 0 dso_as512512512\[12\]
rlabel metal2 447166 373813 447166 373813 0 dso_as512512512\[13\]
rlabel metal2 411930 449854 411930 449854 0 dso_as512512512\[14\]
rlabel metal2 447166 375173 447166 375173 0 dso_as512512512\[15\]
rlabel metal2 447258 376193 447258 376193 0 dso_as512512512\[16\]
rlabel metal2 447166 376499 447166 376499 0 dso_as512512512\[17\]
rlabel metal2 367770 473348 367770 473348 0 dso_as512512512\[18\]
rlabel metal2 370530 478856 370530 478856 0 dso_as512512512\[19\]
rlabel metal1 444820 365602 444820 365602 0 dso_as512512512\[1\]
rlabel metal2 371910 485078 371910 485078 0 dso_as512512512\[20\]
rlabel metal2 447166 379253 447166 379253 0 dso_as512512512\[21\]
rlabel metal2 410550 496774 410550 496774 0 dso_as512512512\[22\]
rlabel metal2 447166 380647 447166 380647 0 dso_as512512512\[23\]
rlabel metal2 407790 508470 407790 508470 0 dso_as512512512\[24\]
rlabel metal2 447166 382007 447166 382007 0 dso_as512512512\[25\]
rlabel metal2 406410 519860 406410 519860 0 dso_as512512512\[26\]
rlabel metal2 447166 383401 447166 383401 0 dso_as512512512\[27\]
rlabel metal2 447258 366571 447258 366571 0 dso_as512512512\[2\]
rlabel metal2 447166 366945 447166 366945 0 dso_as512512512\[3\]
rlabel metal1 444774 368390 444774 368390 0 dso_as512512512\[4\]
rlabel metal1 445418 368458 445418 368458 0 dso_as512512512\[5\]
rlabel metal2 447258 369359 447258 369359 0 dso_as512512512\[6\]
rlabel metal2 447166 369665 447166 369665 0 dso_as512512512\[7\]
rlabel metal2 447258 370719 447258 370719 0 dso_as512512512\[8\]
rlabel metal2 447166 371025 447166 371025 0 dso_as512512512\[9\]
rlabel metal2 483177 385900 483177 385900 0 dso_as5401\[0\]
rlabel metal2 490590 389256 490590 389256 0 dso_as5401\[10\]
rlabel metal2 491326 386451 491326 386451 0 dso_as5401\[11\]
rlabel metal2 491825 385900 491825 385900 0 dso_as5401\[12\]
rlabel metal2 537779 425068 537779 425068 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 483775 385900 483775 385900 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498449 385900 498449 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406164 522330 406164 0 dso_as5401\[22\]
rlabel metal2 499921 385900 499921 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387352 500894 387352 0 dso_as5401\[24\]
rlabel metal2 501393 385900 501393 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387318 502366 387318 0 dso_as5401\[26\]
rlabel metal2 484702 387420 484702 387420 0 dso_as5401\[2\]
rlabel metal2 485438 387284 485438 387284 0 dso_as5401\[3\]
rlabel metal2 485983 385900 485983 385900 0 dso_as5401\[4\]
rlabel metal2 486910 387250 486910 387250 0 dso_as5401\[5\]
rlabel metal2 487409 385900 487409 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387182 488382 387182 0 dso_as5401\[7\]
rlabel metal2 488881 385900 488881 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387216 489854 387216 0 dso_as5401\[9\]
rlabel metal2 523710 368628 523710 368628 0 dso_counter\[0\]
rlabel metal2 565570 359526 565570 359526 0 dso_counter\[10\]
rlabel metal2 567042 359458 567042 359458 0 dso_counter\[11\]
rlabel metal2 547170 368730 547170 368730 0 dso_counter\[1\]
rlabel metal2 544410 369308 544410 369308 0 dso_counter\[2\]
rlabel metal3 511052 380324 511052 380324 0 dso_counter\[3\]
rlabel metal3 511190 380868 511190 380868 0 dso_counter\[4\]
rlabel metal2 558210 359594 558210 359594 0 dso_counter\[5\]
rlabel metal2 559682 359254 559682 359254 0 dso_counter\[6\]
rlabel metal2 561154 359322 561154 359322 0 dso_counter\[7\]
rlabel metal2 519662 370532 519662 370532 0 dso_counter\[8\]
rlabel metal2 522330 370396 522330 370396 0 dso_counter\[9\]
rlabel metal2 456734 387522 456734 387522 0 dso_diceroll\[0\]
rlabel metal2 457233 385900 457233 385900 0 dso_diceroll\[1\]
rlabel metal1 467590 429930 467590 429930 0 dso_diceroll\[2\]
rlabel metal2 458705 385900 458705 385900 0 dso_diceroll\[3\]
rlabel metal2 463634 390660 463634 390660 0 dso_diceroll\[4\]
rlabel metal2 484978 430994 484978 430994 0 dso_diceroll\[5\]
rlabel metal2 461097 385900 461097 385900 0 dso_diceroll\[6\]
rlabel metal2 461695 385900 461695 385900 0 dso_diceroll\[7\]
rlabel metal3 448876 352580 448876 352580 0 dso_mc14500\[0\]
rlabel metal3 449566 353260 449566 353260 0 dso_mc14500\[1\]
rlabel metal3 449842 353940 449842 353940 0 dso_mc14500\[2\]
rlabel metal3 449612 354620 449612 354620 0 dso_mc14500\[3\]
rlabel metal2 484902 500140 484902 500140 0 dso_mc14500\[4\]
rlabel metal2 486190 500140 486190 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 488766 500140 488766 500140 0 dso_mc14500\[7\]
rlabel via2 450133 358428 450133 358428 0 dso_mc14500\[8\]
rlabel metal2 450793 385900 450793 385900 0 dso_multiplier\[0\]
rlabel metal2 451437 385900 451437 385900 0 dso_multiplier\[1\]
rlabel metal2 452081 385900 452081 385900 0 dso_multiplier\[2\]
rlabel metal2 452955 385900 452955 385900 0 dso_multiplier\[3\]
rlabel metal2 453790 387522 453790 387522 0 dso_multiplier\[4\]
rlabel metal2 454335 385900 454335 385900 0 dso_multiplier\[5\]
rlabel metal2 455071 385900 455071 385900 0 dso_multiplier\[6\]
rlabel metal2 461058 498518 461058 498518 0 dso_multiplier\[7\]
rlabel metal1 507978 307122 507978 307122 0 dso_posit\[0\]
rlabel metal3 530004 226236 530004 226236 0 dso_posit\[1\]
rlabel metal3 530004 243644 530004 243644 0 dso_posit\[2\]
rlabel metal3 529391 261596 529391 261596 0 dso_posit\[3\]
rlabel metal2 447166 359091 447166 359091 0 dso_tbb1143\[0\]
rlabel metal2 447258 359465 447258 359465 0 dso_tbb1143\[1\]
rlabel metal2 447166 360485 447166 360485 0 dso_tbb1143\[2\]
rlabel metal1 444866 360298 444866 360298 0 dso_tbb1143\[3\]
rlabel metal2 447166 361845 447166 361845 0 dso_tbb1143\[4\]
rlabel metal1 445464 361658 445464 361658 0 dso_tbb1143\[5\]
rlabel metal1 444774 363018 444774 363018 0 dso_tbb1143\[6\]
rlabel metal2 447166 363545 447166 363545 0 dso_tbb1143\[7\]
rlabel metal1 502550 319464 502550 319464 0 dso_tune
rlabel metal2 502366 318087 502366 318087 0 dso_vgatest\[0\]
rlabel metal2 407806 104924 407806 104924 0 dso_vgatest\[1\]
rlabel metal2 503010 319124 503010 319124 0 dso_vgatest\[2\]
rlabel metal2 450754 211208 450754 211208 0 dso_vgatest\[3\]
rlabel metal2 426680 104924 426680 104924 0 dso_vgatest\[4\]
rlabel metal2 504206 316652 504206 316652 0 dso_vgatest\[5\]
rlabel metal2 450662 211276 450662 211276 0 dso_vgatest\[6\]
rlabel metal2 445172 104924 445172 104924 0 dso_vgatest\[7\]
rlabel metal2 451198 104924 451198 104924 0 dso_vgatest\[8\]
rlabel metal2 505257 322116 505257 322116 0 dso_vgatest\[9\]
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal3 582046 458116 582046 458116 0 io_in[10]
rlabel metal2 580198 510969 580198 510969 0 io_in[11]
rlabel metal3 582000 564332 582000 564332 0 io_in[12]
rlabel metal3 581954 617508 581954 617508 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal3 559567 699788 559567 699788 0 io_in[15]
rlabel via2 444245 422076 444245 422076 0 io_in[16]
rlabel metal2 429870 701940 429870 701940 0 io_in[17]
rlabel metal2 365010 702212 365010 702212 0 io_in[18]
rlabel metal4 444268 510816 444268 510816 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 235198 702144 235198 702144 0 io_in[20]
rlabel metal4 446292 511088 446292 511088 0 io_in[21]
rlabel metal3 444245 421804 444245 421804 0 io_in[22]
rlabel metal2 40526 701974 40526 701974 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 2016 632060 2016 632060 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal2 3542 678436 3542 678436 0 io_in[28]
rlabel metal3 2016 423572 2016 423572 0 io_in[29]
rlabel metal3 581218 86156 581218 86156 0 io_in[2]
rlabel metal1 4600 218042 4600 218042 0 io_in[30]
rlabel metal1 4324 259386 4324 259386 0 io_in[31]
rlabel metal3 1924 267172 1924 267172 0 io_in[32]
rlabel metal3 2108 214948 2108 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1947 110636 1947 110636 0 io_in[35]
rlabel metal3 1740 71604 1740 71604 0 io_in[36]
rlabel metal3 1924 32436 1924 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 461610 308754 461610 308754 0 io_in[7]
rlabel metal3 582138 351900 582138 351900 0 io_in[8]
rlabel metal3 582092 404940 582092 404940 0 io_in[9]
rlabel metal2 565110 171428 565110 171428 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 519570 428366 519570 428366 0 io_oeb[11]
rlabel metal2 579646 590835 579646 590835 0 io_oeb[12]
rlabel metal3 581218 644028 581218 644028 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 527206 701685 527206 701685 0 io_oeb[15]
rlabel metal1 446430 322422 446430 322422 0 io_oeb[16]
rlabel metal2 446522 510850 446522 510850 0 io_oeb[17]
rlabel metal2 332534 702093 332534 702093 0 io_oeb[18]
rlabel metal2 442566 328474 442566 328474 0 io_oeb[19]
rlabel metal2 544410 181050 544410 181050 0 io_oeb[1]
rlabel metal2 445326 503030 445326 503030 0 io_oeb[20]
rlabel metal2 137862 702076 137862 702076 0 io_oeb[21]
rlabel metal3 443831 421940 443831 421940 0 io_oeb[22]
rlabel metal2 442750 328831 442750 328831 0 io_oeb[23]
rlabel metal3 1740 658172 1740 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal3 2200 553860 2200 553860 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1878 449548 1878 449548 0 io_oeb[28]
rlabel metal2 465750 272034 465750 272034 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal3 1924 345372 1924 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 2062 241060 2062 241060 0 io_oeb[32]
rlabel metal3 2200 188836 2200 188836 0 io_oeb[33]
rlabel metal3 1855 136748 1855 136748 0 io_oeb[34]
rlabel metal3 1740 84660 1740 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580014 232781 580014 232781 0 io_oeb[5]
rlabel metal2 580198 272697 580198 272697 0 io_oeb[6]
rlabel metal2 580198 324785 580198 324785 0 io_oeb[7]
rlabel metal2 579646 378301 579646 378301 0 io_oeb[8]
rlabel metal2 579646 431103 579646 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 467774 321956 467774 321956 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 579646 577269 579646 577269 0 io_out[12]
rlabel metal2 468602 321718 468602 321718 0 io_out[13]
rlabel metal2 468878 320970 468878 320970 0 io_out[14]
rlabel metal2 469154 321038 469154 321038 0 io_out[15]
rlabel metal1 446016 423402 446016 423402 0 io_out[16]
rlabel metal2 449190 328984 449190 328984 0 io_out[17]
rlabel metal2 347806 693811 347806 693811 0 io_out[18]
rlabel metal2 446614 511564 446614 511564 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 218454 703596 218454 703596 0 io_out[20]
rlabel metal2 154146 702110 154146 702110 0 io_out[21]
rlabel metal4 446476 502588 446476 502588 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 2039 671228 2039 671228 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal1 3772 678538 3772 678538 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal2 422878 192916 422878 192916 0 io_out[30]
rlabel metal3 2016 306204 2016 306204 0 io_out[31]
rlabel metal3 1970 254116 1970 254116 0 io_out[32]
rlabel metal3 2154 201892 2154 201892 0 io_out[33]
rlabel metal3 1786 149804 1786 149804 0 io_out[34]
rlabel metal3 2016 97580 2016 97580 0 io_out[35]
rlabel metal3 1740 58548 1740 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal2 580198 219215 580198 219215 0 io_out[5]
rlabel metal2 466617 322116 466617 322116 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 467682 322031 467682 322031 0 io_out[9]
rlabel metal2 451582 158321 451582 158321 0 oeb_6502
rlabel metal3 539281 137972 539281 137972 0 oeb_as1802
rlabel metal2 462477 385900 462477 385900 0 oeb_as2650
rlabel metal2 447166 384421 447166 384421 0 oeb_as512512512
rlabel metal2 502865 385900 502865 385900 0 oeb_as5401
rlabel via2 450317 358836 450317 358836 0 oeb_mc14500
rlabel metal2 448010 159868 448010 159868 0 rst_6502
rlabel metal2 427478 446070 427478 446070 0 rst_LCD
rlabel metal3 449980 345100 449980 345100 0 rst_as1802
rlabel metal3 449980 345780 449980 345780 0 rst_as2650
rlabel metal2 447166 347429 447166 347429 0 rst_as512512512
rlabel metal3 450041 346868 450041 346868 0 rst_as5401
rlabel metal3 448922 347820 448922 347820 0 rst_counter
rlabel metal3 448968 348500 448968 348500 0 rst_diceroll
rlabel metal3 449290 349180 449290 349180 0 rst_mc14500
rlabel metal3 449934 349860 449934 349860 0 rst_posit
rlabel via2 447166 350557 447166 350557 0 rst_tbb1143
rlabel metal3 448784 351220 448784 351220 0 rst_tune
rlabel via2 447166 351917 447166 351917 0 rst_vgatest
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1911 1702 1911 0 wb_rst_i
rlabel metal2 2898 1214 2898 1214 0 wbs_ack_o
rlabel metal3 194580 44812 194580 44812 0 wbs_adr_i[0]
rlabel metal2 47649 340 47649 340 0 wbs_adr_i[10]
rlabel metal2 51237 340 51237 340 0 wbs_adr_i[11]
rlabel metal1 216476 44982 216476 44982 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 65313 340 65313 340 0 wbs_adr_i[15]
rlabel metal1 222686 45254 222686 45254 0 wbs_adr_i[16]
rlabel metal1 224020 44778 224020 44778 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 373566 171071 373566 171071 0 wbs_adr_i[1]
rlabel metal2 83076 16560 83076 16560 0 wbs_adr_i[20]
rlabel metal2 370990 171428 370990 171428 0 wbs_adr_i[21]
rlabel metal2 370806 171394 370806 171394 0 wbs_adr_i[22]
rlabel metal2 93978 3627 93978 3627 0 wbs_adr_i[23]
rlabel metal2 97060 16560 97060 16560 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 367770 171496 367770 171496 0 wbs_adr_i[26]
rlabel metal2 368046 171462 368046 171462 0 wbs_adr_i[27]
rlabel metal2 367954 171428 367954 171428 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 1894 17066 1894 0 wbs_adr_i[2]
rlabel metal2 118818 3627 118818 3627 0 wbs_adr_i[30]
rlabel metal2 121900 16560 121900 16560 0 wbs_adr_i[31]
rlabel metal2 21298 16560 21298 16560 0 wbs_adr_i[3]
rlabel metal2 507794 309230 507794 309230 0 wbs_adr_i[4]
rlabel metal1 195730 39610 195730 39610 0 wbs_adr_i[5]
rlabel metal1 198444 39678 198444 39678 0 wbs_adr_i[6]
rlabel metal2 37214 1248 37214 1248 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 1282 44298 1282 0 wbs_adr_i[9]
rlabel metal2 3857 340 3857 340 0 wbs_cyc_i
rlabel metal2 372002 150756 372002 150756 0 wbs_dat_i[0]
rlabel metal2 365010 150722 365010 150722 0 wbs_dat_i[10]
rlabel metal1 208150 39746 208150 39746 0 wbs_dat_i[11]
rlabel metal2 55660 16560 55660 16560 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal2 365470 167314 365470 167314 0 wbs_dat_i[15]
rlabel metal2 366482 165682 366482 165682 0 wbs_dat_i[16]
rlabel metal2 369242 165648 369242 165648 0 wbs_dat_i[17]
rlabel metal2 77418 2132 77418 2132 0 wbs_dat_i[18]
rlabel metal2 80500 16560 80500 16560 0 wbs_dat_i[19]
rlabel metal2 372186 149192 372186 149192 0 wbs_dat_i[1]
rlabel metal2 373382 165886 373382 165886 0 wbs_dat_i[20]
rlabel metal2 372278 165886 372278 165886 0 wbs_dat_i[21]
rlabel metal2 519018 328576 519018 328576 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102212 16560 102212 16560 0 wbs_dat_i[25]
rlabel metal2 518926 330276 518926 330276 0 wbs_dat_i[26]
rlabel metal2 109197 340 109197 340 0 wbs_dat_i[27]
rlabel metal2 507518 307462 507518 307462 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18117 340 18117 340 0 wbs_dat_i[2]
rlabel metal2 119370 16560 119370 16560 0 wbs_dat_i[30]
rlabel metal2 123273 340 123273 340 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 385802 147662 385802 147662 0 wbs_dat_i[4]
rlabel metal2 386354 163098 386354 163098 0 wbs_dat_i[5]
rlabel metal2 520674 314466 520674 314466 0 wbs_dat_i[6]
rlabel metal2 38410 1996 38410 1996 0 wbs_dat_i[7]
rlabel metal2 41676 16560 41676 16560 0 wbs_dat_i[8]
rlabel metal2 45257 340 45257 340 0 wbs_dat_i[9]
rlabel metal2 507334 306153 507334 306153 0 wbs_dat_o[0]
rlabel metal2 366666 161738 366666 161738 0 wbs_dat_o[10]
rlabel metal2 53774 2098 53774 2098 0 wbs_dat_o[11]
rlabel metal2 57033 340 57033 340 0 wbs_dat_o[12]
rlabel metal2 60858 15766 60858 15766 0 wbs_dat_o[13]
rlabel metal2 63940 16560 63940 16560 0 wbs_dat_o[14]
rlabel metal2 522054 320654 522054 320654 0 wbs_dat_o[15]
rlabel metal2 519110 321538 519110 321538 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78377 340 78377 340 0 wbs_dat_o[18]
rlabel metal2 82110 2166 82110 2166 0 wbs_dat_o[19]
rlabel metal2 384790 160055 384790 160055 0 wbs_dat_o[1]
rlabel metal2 85698 2234 85698 2234 0 wbs_dat_o[20]
rlabel metal2 385894 167960 385894 167960 0 wbs_dat_o[21]
rlabel metal2 92637 340 92637 340 0 wbs_dat_o[22]
rlabel metal2 96278 2200 96278 2200 0 wbs_dat_o[23]
rlabel metal2 99636 16560 99636 16560 0 wbs_dat_o[24]
rlabel metal2 103362 1860 103362 1860 0 wbs_dat_o[25]
rlabel metal2 369150 160412 369150 160412 0 wbs_dat_o[26]
rlabel metal2 110538 1792 110538 1792 0 wbs_dat_o[27]
rlabel metal2 113620 16560 113620 16560 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19412 16560 19412 16560 0 wbs_dat_o[2]
rlabel metal2 121118 1792 121118 1792 0 wbs_dat_o[30]
rlabel metal1 446108 386410 446108 386410 0 wbs_dat_o[31]
rlabel metal2 24242 1928 24242 1928 0 wbs_dat_o[3]
rlabel metal2 386170 157454 386170 157454 0 wbs_dat_o[4]
rlabel metal2 522330 310964 522330 310964 0 wbs_dat_o[5]
rlabel metal2 35972 16560 35972 16560 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal2 46690 2030 46690 2030 0 wbs_dat_o[9]
rlabel metal2 5290 2183 5290 2183 0 wbs_stb_i
rlabel metal2 6486 1979 6486 1979 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
