magic
tech sky130B
magscale 1 2
timestamp 1680173551
<< nwell >>
rect 1066 56837 58918 57403
rect 1066 55749 58918 56315
rect 1066 54661 58918 55227
rect 1066 53573 58918 54139
rect 1066 52485 58918 53051
rect 1066 51397 58918 51963
rect 1066 50309 58918 50875
rect 1066 49221 58918 49787
rect 1066 48133 58918 48699
rect 1066 47045 58918 47611
rect 1066 45957 58918 46523
rect 1066 44869 58918 45435
rect 1066 43781 58918 44347
rect 1066 42693 58918 43259
rect 1066 41605 58918 42171
rect 1066 40517 58918 41083
rect 1066 39429 58918 39995
rect 1066 38341 58918 38907
rect 1066 37253 58918 37819
rect 1066 36165 58918 36731
rect 1066 35077 58918 35643
rect 1066 33989 58918 34555
rect 1066 32901 58918 33467
rect 1066 31813 58918 32379
rect 1066 30725 58918 31291
rect 1066 29637 58918 30203
rect 1066 28549 58918 29115
rect 1066 27461 58918 28027
rect 1066 26373 58918 26939
rect 1066 25285 58918 25851
rect 1066 24197 58918 24763
rect 1066 23109 58918 23675
rect 1066 22021 58918 22587
rect 1066 20933 58918 21499
rect 1066 19845 58918 20411
rect 1066 18757 58918 19323
rect 1066 17669 58918 18235
rect 1066 16581 58918 17147
rect 1066 15493 58918 16059
rect 1066 14405 58918 14971
rect 1066 13317 58918 13883
rect 1066 12229 58918 12795
rect 1066 11141 58918 11707
rect 1066 10053 58918 10619
rect 1066 8965 58918 9531
rect 1066 7877 58918 8443
rect 1066 6789 58918 7355
rect 1066 5701 58918 6267
rect 1066 4613 58918 5179
rect 1066 3525 58918 4091
rect 1066 2437 58918 3003
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 2128 58880 57712
<< metal2 >>
rect 2226 59200 2282 60000
rect 6182 59200 6238 60000
rect 10138 59200 10194 60000
rect 14094 59200 14150 60000
rect 18050 59200 18106 60000
rect 22006 59200 22062 60000
rect 25962 59200 26018 60000
rect 29918 59200 29974 60000
rect 33874 59200 33930 60000
rect 37830 59200 37886 60000
rect 41786 59200 41842 60000
rect 45742 59200 45798 60000
rect 49698 59200 49754 60000
rect 53654 59200 53710 60000
rect 57610 59200 57666 60000
<< obsm2 >>
rect 1952 59144 2170 59200
rect 2338 59144 6126 59200
rect 6294 59144 10082 59200
rect 10250 59144 14038 59200
rect 14206 59144 17994 59200
rect 18162 59144 21950 59200
rect 22118 59144 25906 59200
rect 26074 59144 29862 59200
rect 30030 59144 33818 59200
rect 33986 59144 37774 59200
rect 37942 59144 41730 59200
rect 41898 59144 45686 59200
rect 45854 59144 49642 59200
rect 49810 59144 53598 59200
rect 53766 59144 57554 59200
rect 57722 59144 58492 59200
rect 1952 2139 58492 59144
<< metal3 >>
rect 59200 57400 60000 57520
rect 59200 55360 60000 55480
rect 59200 53320 60000 53440
rect 59200 51280 60000 51400
rect 59200 49240 60000 49360
rect 59200 47200 60000 47320
rect 59200 45160 60000 45280
rect 59200 43120 60000 43240
rect 59200 41080 60000 41200
rect 59200 39040 60000 39160
rect 59200 37000 60000 37120
rect 59200 34960 60000 35080
rect 59200 32920 60000 33040
rect 59200 30880 60000 31000
rect 59200 28840 60000 28960
rect 59200 26800 60000 26920
rect 59200 24760 60000 24880
rect 59200 22720 60000 22840
rect 59200 20680 60000 20800
rect 59200 18640 60000 18760
rect 59200 16600 60000 16720
rect 59200 14560 60000 14680
rect 59200 12520 60000 12640
rect 59200 10480 60000 10600
rect 59200 8440 60000 8560
rect 59200 6400 60000 6520
rect 59200 4360 60000 4480
rect 59200 2320 60000 2440
<< obsm3 >>
rect 3325 57600 59200 57697
rect 3325 57320 59120 57600
rect 3325 55560 59200 57320
rect 3325 55280 59120 55560
rect 3325 53520 59200 55280
rect 3325 53240 59120 53520
rect 3325 51480 59200 53240
rect 3325 51200 59120 51480
rect 3325 49440 59200 51200
rect 3325 49160 59120 49440
rect 3325 47400 59200 49160
rect 3325 47120 59120 47400
rect 3325 45360 59200 47120
rect 3325 45080 59120 45360
rect 3325 43320 59200 45080
rect 3325 43040 59120 43320
rect 3325 41280 59200 43040
rect 3325 41000 59120 41280
rect 3325 39240 59200 41000
rect 3325 38960 59120 39240
rect 3325 37200 59200 38960
rect 3325 36920 59120 37200
rect 3325 35160 59200 36920
rect 3325 34880 59120 35160
rect 3325 33120 59200 34880
rect 3325 32840 59120 33120
rect 3325 31080 59200 32840
rect 3325 30800 59120 31080
rect 3325 29040 59200 30800
rect 3325 28760 59120 29040
rect 3325 27000 59200 28760
rect 3325 26720 59120 27000
rect 3325 24960 59200 26720
rect 3325 24680 59120 24960
rect 3325 22920 59200 24680
rect 3325 22640 59120 22920
rect 3325 20880 59200 22640
rect 3325 20600 59120 20880
rect 3325 18840 59200 20600
rect 3325 18560 59120 18840
rect 3325 16800 59200 18560
rect 3325 16520 59120 16800
rect 3325 14760 59200 16520
rect 3325 14480 59120 14760
rect 3325 12720 59200 14480
rect 3325 12440 59120 12720
rect 3325 10680 59200 12440
rect 3325 10400 59120 10680
rect 3325 8640 59200 10400
rect 3325 8360 59120 8640
rect 3325 6600 59200 8360
rect 3325 6320 59120 6600
rect 3325 4560 59200 6320
rect 3325 4280 59120 4560
rect 3325 2520 59200 4280
rect 3325 2240 59120 2520
rect 3325 2143 59200 2240
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 7603 4659 19488 57221
rect 19968 4659 34848 57221
rect 35328 4659 50208 57221
rect 50688 4659 53669 57221
<< labels >>
rlabel metal2 s 53654 59200 53710 60000 6 clk
port 1 nsew signal input
rlabel metal2 s 2226 59200 2282 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 41786 59200 41842 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 45742 59200 45798 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 49698 59200 49754 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 6182 59200 6238 60000 6 io_in[1]
port 6 nsew signal input
rlabel metal2 s 10138 59200 10194 60000 6 io_in[2]
port 7 nsew signal input
rlabel metal2 s 14094 59200 14150 60000 6 io_in[3]
port 8 nsew signal input
rlabel metal2 s 18050 59200 18106 60000 6 io_in[4]
port 9 nsew signal input
rlabel metal2 s 22006 59200 22062 60000 6 io_in[5]
port 10 nsew signal input
rlabel metal2 s 25962 59200 26018 60000 6 io_in[6]
port 11 nsew signal input
rlabel metal2 s 29918 59200 29974 60000 6 io_in[7]
port 12 nsew signal input
rlabel metal2 s 33874 59200 33930 60000 6 io_in[8]
port 13 nsew signal input
rlabel metal2 s 37830 59200 37886 60000 6 io_in[9]
port 14 nsew signal input
rlabel metal3 s 59200 57400 60000 57520 6 io_oeb
port 15 nsew signal output
rlabel metal3 s 59200 2320 60000 2440 6 io_out[0]
port 16 nsew signal output
rlabel metal3 s 59200 22720 60000 22840 6 io_out[10]
port 17 nsew signal output
rlabel metal3 s 59200 24760 60000 24880 6 io_out[11]
port 18 nsew signal output
rlabel metal3 s 59200 26800 60000 26920 6 io_out[12]
port 19 nsew signal output
rlabel metal3 s 59200 28840 60000 28960 6 io_out[13]
port 20 nsew signal output
rlabel metal3 s 59200 30880 60000 31000 6 io_out[14]
port 21 nsew signal output
rlabel metal3 s 59200 32920 60000 33040 6 io_out[15]
port 22 nsew signal output
rlabel metal3 s 59200 34960 60000 35080 6 io_out[16]
port 23 nsew signal output
rlabel metal3 s 59200 37000 60000 37120 6 io_out[17]
port 24 nsew signal output
rlabel metal3 s 59200 39040 60000 39160 6 io_out[18]
port 25 nsew signal output
rlabel metal3 s 59200 41080 60000 41200 6 io_out[19]
port 26 nsew signal output
rlabel metal3 s 59200 4360 60000 4480 6 io_out[1]
port 27 nsew signal output
rlabel metal3 s 59200 43120 60000 43240 6 io_out[20]
port 28 nsew signal output
rlabel metal3 s 59200 45160 60000 45280 6 io_out[21]
port 29 nsew signal output
rlabel metal3 s 59200 47200 60000 47320 6 io_out[22]
port 30 nsew signal output
rlabel metal3 s 59200 49240 60000 49360 6 io_out[23]
port 31 nsew signal output
rlabel metal3 s 59200 51280 60000 51400 6 io_out[24]
port 32 nsew signal output
rlabel metal3 s 59200 53320 60000 53440 6 io_out[25]
port 33 nsew signal output
rlabel metal3 s 59200 55360 60000 55480 6 io_out[26]
port 34 nsew signal output
rlabel metal3 s 59200 6400 60000 6520 6 io_out[2]
port 35 nsew signal output
rlabel metal3 s 59200 8440 60000 8560 6 io_out[3]
port 36 nsew signal output
rlabel metal3 s 59200 10480 60000 10600 6 io_out[4]
port 37 nsew signal output
rlabel metal3 s 59200 12520 60000 12640 6 io_out[5]
port 38 nsew signal output
rlabel metal3 s 59200 14560 60000 14680 6 io_out[6]
port 39 nsew signal output
rlabel metal3 s 59200 16600 60000 16720 6 io_out[7]
port 40 nsew signal output
rlabel metal3 s 59200 18640 60000 18760 6 io_out[8]
port 41 nsew signal output
rlabel metal3 s 59200 20680 60000 20800 6 io_out[9]
port 42 nsew signal output
rlabel metal2 s 57610 59200 57666 60000 6 rst
port 43 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10009644
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS1802/runs/23_03_30_12_39/results/signoff/wrapped_as1802.magic.gds
string GDS_START 1237642
<< end >>

