VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_6502
  CLASS BLOCK ;
  FOREIGN wrapped_6502 ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 225.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 221.000 195.410 225.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 221.000 11.410 225.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 221.000 29.810 225.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 221.000 48.210 225.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 221.000 66.610 225.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 221.000 85.010 225.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 221.000 103.410 225.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 221.000 121.810 225.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 221.000 140.210 225.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 221.000 158.610 225.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 221.000 177.010 225.000 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 212.880 225.000 213.480 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 10.920 225.000 11.520 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 85.720 225.000 86.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 93.200 225.000 93.800 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 100.680 225.000 101.280 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 108.160 225.000 108.760 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 115.640 225.000 116.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 123.120 225.000 123.720 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 130.600 225.000 131.200 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 138.080 225.000 138.680 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 145.560 225.000 146.160 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 153.040 225.000 153.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 18.400 225.000 19.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 160.520 225.000 161.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 168.000 225.000 168.600 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 175.480 225.000 176.080 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 182.960 225.000 183.560 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 190.440 225.000 191.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 197.920 225.000 198.520 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 205.400 225.000 206.000 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 25.880 225.000 26.480 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 33.360 225.000 33.960 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 40.840 225.000 41.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 48.320 225.000 48.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 55.800 225.000 56.400 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 63.280 225.000 63.880 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 70.760 225.000 71.360 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.000 78.240 225.000 78.840 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 221.000 213.810 225.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 212.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 212.400 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 208.025 219.610 210.855 ;
        RECT 5.330 202.585 219.610 205.415 ;
        RECT 5.330 197.145 219.610 199.975 ;
        RECT 5.330 191.705 219.610 194.535 ;
        RECT 5.330 186.265 219.610 189.095 ;
        RECT 5.330 180.825 219.610 183.655 ;
        RECT 5.330 175.385 219.610 178.215 ;
        RECT 5.330 169.945 219.610 172.775 ;
        RECT 5.330 164.505 219.610 167.335 ;
        RECT 5.330 159.065 219.610 161.895 ;
        RECT 5.330 153.625 219.610 156.455 ;
        RECT 5.330 148.185 219.610 151.015 ;
        RECT 5.330 142.745 219.610 145.575 ;
        RECT 5.330 137.305 219.610 140.135 ;
        RECT 5.330 131.865 219.610 134.695 ;
        RECT 5.330 126.425 219.610 129.255 ;
        RECT 5.330 120.985 219.610 123.815 ;
        RECT 5.330 115.545 219.610 118.375 ;
        RECT 5.330 110.105 219.610 112.935 ;
        RECT 5.330 104.665 219.610 107.495 ;
        RECT 5.330 99.225 219.610 102.055 ;
        RECT 5.330 93.785 219.610 96.615 ;
        RECT 5.330 88.345 219.610 91.175 ;
        RECT 5.330 82.905 219.610 85.735 ;
        RECT 5.330 77.465 219.610 80.295 ;
        RECT 5.330 72.025 219.610 74.855 ;
        RECT 5.330 66.585 219.610 69.415 ;
        RECT 5.330 61.145 219.610 63.975 ;
        RECT 5.330 55.705 219.610 58.535 ;
        RECT 5.330 50.265 219.610 53.095 ;
        RECT 5.330 44.825 219.610 47.655 ;
        RECT 5.330 39.385 219.610 42.215 ;
        RECT 5.330 33.945 219.610 36.775 ;
        RECT 5.330 28.505 219.610 31.335 ;
        RECT 5.330 23.065 219.610 25.895 ;
        RECT 5.330 17.625 219.610 20.455 ;
        RECT 5.330 12.185 219.610 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 219.420 212.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 220.270 220.620 ;
      LAYER met2 ;
        RECT 11.690 220.720 29.250 221.000 ;
        RECT 30.090 220.720 47.650 221.000 ;
        RECT 48.490 220.720 66.050 221.000 ;
        RECT 66.890 220.720 84.450 221.000 ;
        RECT 85.290 220.720 102.850 221.000 ;
        RECT 103.690 220.720 121.250 221.000 ;
        RECT 122.090 220.720 139.650 221.000 ;
        RECT 140.490 220.720 158.050 221.000 ;
        RECT 158.890 220.720 176.450 221.000 ;
        RECT 177.290 220.720 194.850 221.000 ;
        RECT 195.690 220.720 213.250 221.000 ;
        RECT 214.090 220.720 220.250 221.000 ;
        RECT 11.140 10.695 220.250 220.720 ;
      LAYER met3 ;
        RECT 21.050 212.480 220.600 213.345 ;
        RECT 21.050 206.400 221.000 212.480 ;
        RECT 21.050 205.000 220.600 206.400 ;
        RECT 21.050 198.920 221.000 205.000 ;
        RECT 21.050 197.520 220.600 198.920 ;
        RECT 21.050 191.440 221.000 197.520 ;
        RECT 21.050 190.040 220.600 191.440 ;
        RECT 21.050 183.960 221.000 190.040 ;
        RECT 21.050 182.560 220.600 183.960 ;
        RECT 21.050 176.480 221.000 182.560 ;
        RECT 21.050 175.080 220.600 176.480 ;
        RECT 21.050 169.000 221.000 175.080 ;
        RECT 21.050 167.600 220.600 169.000 ;
        RECT 21.050 161.520 221.000 167.600 ;
        RECT 21.050 160.120 220.600 161.520 ;
        RECT 21.050 154.040 221.000 160.120 ;
        RECT 21.050 152.640 220.600 154.040 ;
        RECT 21.050 146.560 221.000 152.640 ;
        RECT 21.050 145.160 220.600 146.560 ;
        RECT 21.050 139.080 221.000 145.160 ;
        RECT 21.050 137.680 220.600 139.080 ;
        RECT 21.050 131.600 221.000 137.680 ;
        RECT 21.050 130.200 220.600 131.600 ;
        RECT 21.050 124.120 221.000 130.200 ;
        RECT 21.050 122.720 220.600 124.120 ;
        RECT 21.050 116.640 221.000 122.720 ;
        RECT 21.050 115.240 220.600 116.640 ;
        RECT 21.050 109.160 221.000 115.240 ;
        RECT 21.050 107.760 220.600 109.160 ;
        RECT 21.050 101.680 221.000 107.760 ;
        RECT 21.050 100.280 220.600 101.680 ;
        RECT 21.050 94.200 221.000 100.280 ;
        RECT 21.050 92.800 220.600 94.200 ;
        RECT 21.050 86.720 221.000 92.800 ;
        RECT 21.050 85.320 220.600 86.720 ;
        RECT 21.050 79.240 221.000 85.320 ;
        RECT 21.050 77.840 220.600 79.240 ;
        RECT 21.050 71.760 221.000 77.840 ;
        RECT 21.050 70.360 220.600 71.760 ;
        RECT 21.050 64.280 221.000 70.360 ;
        RECT 21.050 62.880 220.600 64.280 ;
        RECT 21.050 56.800 221.000 62.880 ;
        RECT 21.050 55.400 220.600 56.800 ;
        RECT 21.050 49.320 221.000 55.400 ;
        RECT 21.050 47.920 220.600 49.320 ;
        RECT 21.050 41.840 221.000 47.920 ;
        RECT 21.050 40.440 220.600 41.840 ;
        RECT 21.050 34.360 221.000 40.440 ;
        RECT 21.050 32.960 220.600 34.360 ;
        RECT 21.050 26.880 221.000 32.960 ;
        RECT 21.050 25.480 220.600 26.880 ;
        RECT 21.050 19.400 221.000 25.480 ;
        RECT 21.050 18.000 220.600 19.400 ;
        RECT 21.050 11.920 221.000 18.000 ;
        RECT 21.050 10.715 220.600 11.920 ;
      LAYER met4 ;
        RECT 40.775 89.255 97.440 207.225 ;
        RECT 99.840 89.255 174.240 207.225 ;
        RECT 176.640 89.255 195.665 207.225 ;
  END
END wrapped_6502
END LIBRARY

