* NGSPICE file created from wrapped_as1802.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt wrapped_as1802 clk io_in[0] io_in[10] io_in[11] io_in[12] io_in[1] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24]
+ io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst vccd1 vssd1
X_3155_ _3209_/A _3209_/B _4157_/B _4184_/B vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__o31a_1
X_3086_ _3086_/A _3086_/B vssd1 vssd1 vccd1 vccd1 _3086_/X sky130_fd_sc_hd__or2_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3988_ _4620_/Q _3991_/B _3988_/C vssd1 vssd1 vccd1 vccd1 _3989_/C sky130_fd_sc_hd__and3_1
X_2939_ _3209_/A _2940_/A _2995_/A vssd1 vssd1 vccd1 vccd1 _2942_/A sky130_fd_sc_hd__o21a_1
X_4609_ _4630_/CLK _4609_/D vssd1 vssd1 vccd1 vccd1 _4609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_as1802_287 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_287/HI io_out[12] sky130_fd_sc_hd__conb_1
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3911_ _4127_/A _4132_/A vssd1 vssd1 vccd1 vccd1 _3911_/Y sky130_fd_sc_hd__nor2_2
X_3842_ _4635_/Q _3802_/B _3836_/A vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _3771_/X _3772_/X _3773_/S vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__mux2_1
X_2724_ _2722_/X _2723_/X _2889_/A vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__mux2_2
X_2655_ _3185_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _2655_/Y sky130_fd_sc_hd__nor2_4
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2586_ _2644_/S _2583_/X _2585_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__o211a_2
X_4325_ _4689_/Q _4336_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4689_/D sky130_fd_sc_hd__mux2_1
Xfanout138 _3632_/X vssd1 vssd1 vccd1 vccd1 _3747_/B2 sky130_fd_sc_hd__buf_4
Xfanout105 _3140_/S vssd1 vssd1 vccd1 vccd1 _3089_/S sky130_fd_sc_hd__clkbuf_8
Xfanout116 _2931_/C1 vssd1 vssd1 vccd1 vccd1 _3139_/A sky130_fd_sc_hd__buf_6
Xfanout127 _2424_/X vssd1 vssd1 vccd1 vccd1 _2846_/S sky130_fd_sc_hd__buf_4
X_4256_ _4256_/A1 _4254_/X _4255_/Y vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__a21o_1
Xfanout149 _2863_/B vssd1 vssd1 vccd1 vccd1 _2927_/B sky130_fd_sc_hd__buf_4
X_4187_ _3908_/B _4161_/Y _4213_/A vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__o21ba_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3207_ _3194_/X _3199_/X _3206_/X _3257_/A1 vssd1 vssd1 vccd1 vccd1 _3283_/A sky130_fd_sc_hd__o22a_4
X_3138_ _4505_/Q _4561_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3139_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3287_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _4644_/Q _2440_/B _2440_/C vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__nand3b_2
X_2371_ _3629_/A _3832_/B _2371_/C _2384_/D vssd1 vssd1 vccd1 vccd1 _3185_/A sky130_fd_sc_hd__and4_4
X_4110_ _4059_/A _3072_/B _4109_/Y vssd1 vssd1 vccd1 vccd1 _4110_/X sky130_fd_sc_hd__a21o_1
X_4041_ _2351_/C _3396_/B _4040_/X _3608_/A vssd1 vssd1 vccd1 vccd1 _4054_/B sky130_fd_sc_hd__a31o_1
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3825_ _4629_/Q _4605_/Q _3827_/S vssd1 vssd1 vccd1 vccd1 _3826_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3756_ _3989_/B _3755_/X _4184_/B _3632_/X vssd1 vssd1 vccd1 vccd1 _3756_/X sky130_fd_sc_hd__a2bb2o_1
X_2707_ _2938_/A1 _2702_/X _2706_/X _2697_/X _2698_/X vssd1 vssd1 vccd1 vccd1 _2848_/A
+ sky130_fd_sc_hd__o32ai_4
X_3687_ _3731_/A1 _2848_/A _3739_/B _3685_/X _3686_/Y vssd1 vssd1 vccd1 vccd1 _3687_/X
+ sky130_fd_sc_hd__a221o_2
X_2638_ _2933_/C1 _2633_/X _2635_/X _2637_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2638_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2569_ _4484_/Q _4485_/Q _4486_/Q vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__o21a_1
X_4308_ _4062_/A _4307_/X _4270_/X vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4239_ _4239_/A _4239_/B _4232_/X vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__or3b_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4590_ _4692_/CLK _4590_/D vssd1 vssd1 vccd1 vccd1 _4590_/Q sky130_fd_sc_hd__dfxtp_4
X_3610_ _2360_/A _2473_/B _3847_/B _2356_/B vssd1 vssd1 vccd1 vccd1 _3610_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3541_ _4552_/Q _3541_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4552_/D sky130_fd_sc_hd__mux2_1
X_3472_ _4491_/Q _3544_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4491_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2423_ _2424_/A _2424_/B vssd1 vssd1 vccd1 vccd1 _3020_/S sky130_fd_sc_hd__nor2_8
X_2354_ _2354_/A _2354_/B vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__or2_4
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2285_ _3581_/B _3581_/D vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__nand2_2
X_4024_ _4665_/Q _4649_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3808_ _3689_/A input7/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4618_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3739_ _3739_/A _3739_/B vssd1 vssd1 vccd1 vccd1 _3739_/X sky130_fd_sc_hd__or2_1
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2972_ _4685_/Q _2971_/B _2389_/A vssd1 vssd1 vccd1 vccd1 _2972_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4642_ _4702_/CLK _4642_/D vssd1 vssd1 vccd1 vccd1 _4642_/Q sky130_fd_sc_hd__dfxtp_1
X_4573_ _4573_/CLK _4573_/D vssd1 vssd1 vccd1 vccd1 _4573_/Q sky130_fd_sc_hd__dfxtp_1
X_3524_ _4537_/Q _3569_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4537_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3455_ _3572_/A _3536_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _3463_/S sky130_fd_sc_hd__and3_4
X_2406_ _2404_/A _2406_/B vssd1 vssd1 vccd1 vccd1 _2406_/Y sky130_fd_sc_hd__nand2b_1
X_3386_ _2290_/B _3640_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3833_/A sky130_fd_sc_hd__o21a_1
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2337_ _2904_/A _2337_/B _2337_/C vssd1 vssd1 vccd1 vccd1 _2861_/A sky130_fd_sc_hd__or3_2
X_2268_ _4062_/A _2268_/B _3384_/B vssd1 vssd1 vccd1 vccd1 _2268_/X sky130_fd_sc_hd__and3_1
X_4007_ _4011_/A _4006_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4007_/X sky130_fd_sc_hd__a21bo_1
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _2195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3226_/X _3236_/X _3239_/X vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3751_/B vssd1 vssd1 vccd1 vccd1 _3273_/C sky130_fd_sc_hd__inv_2
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2955_ _2549_/A _2954_/X _2898_/A vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__a21o_1
X_2886_ _2886_/A _2940_/A vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__nor2_1
X_4625_ _4629_/CLK _4625_/D vssd1 vssd1 vccd1 vccd1 _4625_/Q sky130_fd_sc_hd__dfxtp_1
X_4556_ _4580_/CLK _4556_/D vssd1 vssd1 vccd1 vccd1 _4556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3507_ _4522_/Q _3570_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4522_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4487_ _4551_/CLK _4487_/D vssd1 vssd1 vccd1 vccd1 _4487_/Q sky130_fd_sc_hd__dfxtp_2
X_3438_ _4460_/Q _3537_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4460_/D sky130_fd_sc_hd__mux2_1
X_3369_ _4423_/Q _3567_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4423_/D sky130_fd_sc_hd__mux2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput31 _4702_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_4
Xoutput20 _4610_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_4
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _3020_/S _2734_/X _2739_/X vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__a21o_1
X_2671_ _2834_/A _2671_/B vssd1 vssd1 vccd1 vccd1 _2678_/B sky130_fd_sc_hd__or2_1
X_4410_ _4587_/CLK _4410_/D vssd1 vssd1 vccd1 vccd1 _4410_/Q sky130_fd_sc_hd__dfxtp_1
X_4341_ _4341_/A _4341_/B vssd1 vssd1 vccd1 vccd1 _4342_/S sky130_fd_sc_hd__nand2_1
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4272_ _3855_/B _4271_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4663_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3223_ _3223_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__xor2_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3154_ _3212_/A _3185_/C _3288_/A vssd1 vssd1 vccd1 vccd1 _3154_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3085_ _4568_/Q _4528_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3086_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _3987_/A _3987_/B vssd1 vssd1 vccd1 vccd1 _3987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ _2938_/A1 _2933_/X _2937_/X _2924_/X _2929_/X vssd1 vssd1 vccd1 vccd1 _2995_/A
+ sky130_fd_sc_hd__o32ai_4
X_2869_ _4564_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__and3_1
X_4608_ _4630_/CLK _4608_/D vssd1 vssd1 vccd1 vccd1 _4608_/Q sky130_fd_sc_hd__dfxtp_1
X_4539_ _4576_/CLK _4539_/D vssd1 vssd1 vccd1 vccd1 _4539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _4177_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _3910_/X sky130_fd_sc_hd__or2_2
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3841_ _3849_/A _3841_/B _3840_/X vssd1 vssd1 vccd1 vccd1 _4634_/D sky130_fd_sc_hd__or3b_1
XFILLER_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3772_ _4691_/Q _4017_/S _3770_/X _2331_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__o22a_1
X_2723_ _4473_/Q _4465_/Q _4457_/Q _4449_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2723_/X sky130_fd_sc_hd__mux4_1
X_2654_ _2885_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__or2_1
X_2585_ _4487_/Q _2811_/S _2584_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__a211o_1
X_4324_ _4688_/Q _4335_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4688_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout106 _3201_/S vssd1 vssd1 vccd1 vccd1 _3140_/S sky130_fd_sc_hd__buf_6
Xfanout117 _2931_/C1 vssd1 vssd1 vccd1 vccd1 _3252_/S sky130_fd_sc_hd__buf_4
Xfanout128 _2370_/X vssd1 vssd1 vccd1 vccd1 _2389_/A sky130_fd_sc_hd__buf_6
X_4255_ _4256_/A1 _2848_/C _4081_/A vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__o21ai_1
Xfanout139 _2927_/C vssd1 vssd1 vccd1 vccd1 _2804_/C sky130_fd_sc_hd__buf_4
X_4186_ _3907_/B _4161_/Y _4205_/A vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__o21a_1
X_3206_ _3202_/X _3205_/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3137_ _3086_/A _3134_/X _3136_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__o211a_1
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3068_ _3068_/A _3068_/B vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__nor2_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2370_ _2372_/C _4013_/S vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__or2_2
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _4050_/A _4040_/B vssd1 vssd1 vccd1 vccd1 _4040_/X sky130_fd_sc_hd__or2_1
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3824_ _3828_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _4628_/D sky130_fd_sc_hd__nand2_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3755_ _4689_/Q _2242_/X _3691_/C _3754_/X vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__o31a_1
X_2706_ _2814_/A1 _2703_/X _2705_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__o211a_1
X_3686_ _3680_/B _3739_/B _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3686_/Y sky130_fd_sc_hd__o21bai_1
X_2637_ _2805_/C1 _2636_/X _2937_/C1 vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__o21a_1
X_2568_ _3938_/A _2618_/B _3160_/B1 _2567_/X vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4307_ _3855_/B _4278_/Y _4306_/X _4278_/B vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__a22o_1
X_2499_ _4429_/Q _4421_/Q _2661_/S vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__mux2_1
X_4238_ _4238_/A _4238_/B _4238_/C _4237_/X vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__or4b_1
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _4157_/Y _4168_/X _4256_/A1 vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3540_ _4551_/Q _3540_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4551_/D sky130_fd_sc_hd__mux2_1
X_3471_ _4490_/Q _3543_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4490_/D sky130_fd_sc_hd__mux2_1
X_2422_ _2422_/A _2422_/B vssd1 vssd1 vccd1 vccd1 _2422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2353_ _2400_/B _2907_/A vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__or2_2
X_2284_ _2284_/A _2284_/B _2284_/C vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__and3_4
X_4023_ _4037_/A _4023_/B vssd1 vssd1 vccd1 vccd1 _4648_/D sky130_fd_sc_hd__and2_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3807_ _4057_/B input6/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4617_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3738_ _3068_/B _3631_/X _3989_/B _3737_/X vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__o22a_1
X_3669_ _3668_/X _4594_/Q _4329_/S vssd1 vssd1 vccd1 vccd1 _4594_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ _4685_/Q _2971_/B vssd1 vssd1 vccd1 vccd1 _3080_/C sky130_fd_sc_hd__or2_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4641_ _4702_/CLK _4641_/D vssd1 vssd1 vccd1 vccd1 _4641_/Q sky130_fd_sc_hd__dfxtp_1
X_4572_ _4572_/CLK _4572_/D vssd1 vssd1 vccd1 vccd1 _4572_/Q sky130_fd_sc_hd__dfxtp_1
X_3523_ _4536_/Q _3568_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4536_/D sky130_fd_sc_hd__mux2_1
X_3454_ _4475_/Q _3544_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4475_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2405_ _4572_/Q _4516_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _2406_/B sky130_fd_sc_hd__mux2_1
X_3385_ _4011_/A _3385_/B vssd1 vssd1 vccd1 vccd1 _3385_/Y sky130_fd_sc_hd__nand2_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2336_ _2337_/C vssd1 vssd1 vccd1 vccd1 _2844_/A sky130_fd_sc_hd__inv_2
X_2267_ _2473_/A _2293_/A vssd1 vssd1 vccd1 vccd1 _3385_/B sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_49_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4006_ _2373_/B _4005_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2198_ _2889_/A vssd1 vssd1 vccd1 vccd1 _3269_/S sky130_fd_sc_hd__clkinv_4
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _4670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3164_/X _3166_/X _3169_/X _3270_/A vssd1 vssd1 vccd1 vccd1 _3751_/B sky130_fd_sc_hd__o22a_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2954_ _4365_/Q _4694_/Q _4685_/Q _4413_/Q _2892_/S _2954_/S1 vssd1 vssd1 vccd1 vccd1
+ _2954_/X sky130_fd_sc_hd__mux4_2
X_2885_ _2885_/A _2885_/B _2885_/C _2940_/A vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__and4_4
X_4624_ _4691_/CLK _4624_/D vssd1 vssd1 vccd1 vccd1 _4624_/Q sky130_fd_sc_hd__dfxtp_1
X_4555_ _4555_/CLK _4555_/D vssd1 vssd1 vccd1 vccd1 _4555_/Q sky130_fd_sc_hd__dfxtp_1
X_3506_ _4521_/Q _3569_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4521_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4486_ _4490_/CLK _4486_/D vssd1 vssd1 vccd1 vccd1 _4486_/Q sky130_fd_sc_hd__dfxtp_4
X_3437_ _3536_/A _3446_/C _4330_/C vssd1 vssd1 vccd1 vccd1 _3445_/S sky130_fd_sc_hd__and3_4
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3368_ _4422_/Q _3566_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4422_/D sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2319_ _4011_/A _4062_/A vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__nand2_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3318_/A _3299_/B vssd1 vssd1 vccd1 vccd1 _4330_/B sky130_fd_sc_hd__nor2_4
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput21 _4611_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_4
Xoutput32 _4670_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_4
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _2670_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _2671_/B sky130_fd_sc_hd__nor2_1
X_4340_ _4044_/X _4339_/X _4042_/X _4043_/X vssd1 vssd1 vccd1 vccd1 _4341_/B sky130_fd_sc_hd__o211a_1
X_4271_ _4240_/A _4256_/X _4269_/X _4270_/X vssd1 vssd1 vccd1 vccd1 _4271_/X sky130_fd_sc_hd__a31o_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3222_ _3270_/A _3221_/X _3218_/X vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__o21ai_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3153_ _3287_/A _3287_/B _4157_/B _4184_/B vssd1 vssd1 vccd1 vccd1 _3185_/C sky130_fd_sc_hd__a31o_1
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _4359_/Q _4314_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4359_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _4084_/A _3983_/X _3985_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__o211a_1
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2937_ _2937_/A1 _2934_/X _2936_/X _2937_/C1 vssd1 vssd1 vccd1 vccd1 _2937_/X sky130_fd_sc_hd__o211a_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2868_ _4556_/Q _2932_/S _2867_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__a211o_1
X_4607_ _4691_/CLK _4607_/D vssd1 vssd1 vccd1 vccd1 _4607_/Q sky130_fd_sc_hd__dfxtp_1
X_2799_ _4547_/Q _2800_/S _2798_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2799_/X sky130_fd_sc_hd__a211o_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4538_ _4581_/CLK _4538_/D vssd1 vssd1 vccd1 vccd1 _4538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _4667_/CLK _4469_/D vssd1 vssd1 vccd1 vccd1 _4469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3840_ _3617_/B _4692_/Q _3802_/A _3618_/A vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3771_ _3272_/Y _3770_/X _3771_/S vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__mux2_1
X_2722_ _4553_/Q _4497_/Q _4489_/Q _4481_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2722_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2653_ _2885_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2584_ _4479_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__and3_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4323_ _4687_/Q _4334_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4687_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout118 _2438_/Y vssd1 vssd1 vccd1 vccd1 _2931_/C1 sky130_fd_sc_hd__buf_6
Xfanout129 _2370_/X vssd1 vssd1 vccd1 vccd1 _2571_/A sky130_fd_sc_hd__clkbuf_4
Xfanout107 _3254_/S vssd1 vssd1 vccd1 vccd1 _3247_/S sky130_fd_sc_hd__buf_6
X_4254_ _4059_/A _3286_/B _4252_/X _4253_/X vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4185_ _4205_/A _4205_/B _4185_/C vssd1 vssd1 vccd1 vccd1 _4185_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3205_ _3203_/X _3204_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__mux2_1
X_3136_ _4361_/Q _3201_/S _3135_/X _3252_/S vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__a211o_1
X_3067_ _3068_/B vssd1 vssd1 vccd1 vccd1 _3067_/Y sky130_fd_sc_hd__inv_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _3972_/A _4119_/B vssd1 vssd1 vccd1 vccd1 _4082_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3823_ _2183_/Y _2184_/Y _3827_/S vssd1 vssd1 vccd1 vccd1 _3824_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _3754_/A1 _3752_/Y _3753_/X _3773_/S vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2705_ _4457_/Q _2809_/S _2704_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__a211o_1
X_3685_ _3666_/B1 _3684_/X _2848_/A _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3685_/X sky130_fd_sc_hd__a2bb2o_1
X_2636_ _4520_/Q _4576_/Q _2636_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2567_ _3288_/A _2541_/Y _2566_/Y _2363_/B vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__a211o_1
X_4306_ _4647_/Q _2367_/Y _3629_/Y _4655_/Q vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__a22o_1
X_2498_ _2661_/S _4533_/Q _2404_/A vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__a21bo_1
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _3905_/X _4201_/X _4263_/S _4117_/B vssd1 vssd1 vccd1 vccd1 _4237_/X sky130_fd_sc_hd__a211o_1
X_4168_ _3935_/A _4672_/Q _4057_/X _4167_/X _4224_/A vssd1 vssd1 vccd1 vccd1 _4168_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4099_ _3899_/C _4119_/A _3894_/C _3927_/B vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3119_ _3119_/A _3119_/B _3273_/B vssd1 vssd1 vccd1 vccd1 _3173_/A sky130_fd_sc_hd__or3_4
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _4489_/Q _3542_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4489_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2421_ _2904_/A _2421_/B vssd1 vssd1 vccd1 vccd1 _2422_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2352_ _2352_/A _2352_/B vssd1 vssd1 vccd1 vccd1 _3232_/S sky130_fd_sc_hd__or2_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2283_ _4632_/Q _2230_/B _2300_/A vssd1 vssd1 vccd1 vccd1 _2284_/C sky130_fd_sc_hd__a21oi_2
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4022_ _4664_/Q _4648_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4023_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3806_ _4057_/A input5/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4616_/D sky130_fd_sc_hd__mux2_1
X_3737_ _4687_/Q _3762_/B _3691_/C _3736_/X vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__o31a_1
X_3668_ _2669_/C _3749_/A1 _3667_/X _4003_/B vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__o22a_1
X_2619_ _2616_/X _2817_/A vssd1 vssd1 vccd1 vccd1 _2622_/B sky130_fd_sc_hd__and2b_1
X_3599_ _3593_/X _3595_/X _3598_/X _3618_/A vssd1 vssd1 vccd1 vccd1 _3799_/S sky130_fd_sc_hd__a31o_4
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2970_ _2943_/X _2944_/Y _2969_/X vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__o21a_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4643_/CLK _4640_/D vssd1 vssd1 vccd1 vccd1 _4640_/Q sky130_fd_sc_hd__dfxtp_1
X_4571_ _4683_/CLK _4571_/D vssd1 vssd1 vccd1 vccd1 _4571_/Q sky130_fd_sc_hd__dfxtp_1
X_3522_ _4535_/Q _3567_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4535_/D sky130_fd_sc_hd__mux2_1
X_3453_ _4474_/Q _3543_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4474_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2404_ _2404_/A _2404_/B vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3384_ _3384_/A _3384_/B vssd1 vssd1 vccd1 vccd1 _3384_/Y sky130_fd_sc_hd__nor2_2
X_2335_ _3581_/B _3581_/C _2335_/C _2384_/D vssd1 vssd1 vccd1 vccd1 _2337_/C sky130_fd_sc_hd__and4_2
XFILLER_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2266_ _2473_/A _2293_/A vssd1 vssd1 vccd1 vccd1 _3384_/B sky130_fd_sc_hd__nor2_4
X_4005_ _4664_/Q _4672_/Q _4013_/S vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__mux2_1
X_2197_ _4484_/Q vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 _4671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _2953_/A _2953_/B vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__and2_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ _3209_/A _2940_/A _2883_/X vssd1 vssd1 vccd1 vccd1 _2916_/A sky130_fd_sc_hd__a21boi_1
X_4623_ _4626_/CLK _4623_/D vssd1 vssd1 vccd1 vccd1 _4623_/Q sky130_fd_sc_hd__dfxtp_1
X_4554_ _4684_/CLK _4554_/D vssd1 vssd1 vccd1 vccd1 _4554_/Q sky130_fd_sc_hd__dfxtp_1
X_3505_ _4520_/Q _3568_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4520_/D sky130_fd_sc_hd__mux2_1
X_4485_ _4490_/CLK _4485_/D vssd1 vssd1 vccd1 vccd1 _4485_/Q sky130_fd_sc_hd__dfxtp_4
X_3436_ _4459_/Q _3571_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4459_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3367_ _4421_/Q _3565_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4421_/D sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2318_ _4011_/A _3581_/C vssd1 vssd1 vccd1 vccd1 _2351_/C sky130_fd_sc_hd__nand2_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3298_ _3328_/A _3298_/B vssd1 vssd1 vccd1 vccd1 _3563_/C sky130_fd_sc_hd__nor2_8
X_2249_ _3846_/A _4615_/Q vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__nand2b_4
XFILLER_26_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput22 _4612_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_4
Xoutput33 _4671_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_4
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4270_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__and2_1
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3221_ _3219_/X _3220_/X _3269_/S vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3152_ _3287_/A _3287_/B _3287_/C vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__nand3_2
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3083_ _3078_/X _3079_/X _3082_/X vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3985_ _3985_/A _3993_/D _4228_/B _3985_/D vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__or4_1
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _4405_/Q _2934_/S _2935_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__a211o_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2867_ _4500_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__and3_1
X_4606_ _4626_/CLK _4606_/D vssd1 vssd1 vccd1 vccd1 _4606_/Q sky130_fd_sc_hd__dfxtp_2
X_2798_ _4539_/Q _2798_/B _2798_/C vssd1 vssd1 vccd1 vccd1 _2798_/X sky130_fd_sc_hd__and3_1
X_4537_ _4537_/CLK _4537_/D vssd1 vssd1 vccd1 vccd1 _4537_/Q sky130_fd_sc_hd__dfxtp_1
X_4468_ _4553_/CLK _4468_/D vssd1 vssd1 vccd1 vccd1 _4468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3419_ _3572_/A _3563_/B _3446_/C vssd1 vssd1 vccd1 vccd1 _3427_/S sky130_fd_sc_hd__and3_4
X_4399_ _4679_/CLK _4399_/D vssd1 vssd1 vccd1 vccd1 _4399_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ _3286_/B _3272_/Y _3770_/S vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__mux2_1
X_2721_ _2953_/A _2720_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2652_ _2652_/A _2652_/B vssd1 vssd1 vccd1 vccd1 _2652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _4495_/Q _4551_/Q _2811_/S vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4322_ _4686_/Q _4333_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4686_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _3855_/B _3857_/B _4057_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__o31a_1
Xfanout108 _3254_/S vssd1 vssd1 vccd1 vccd1 _3204_/S sky130_fd_sc_hd__clkbuf_4
Xfanout119 _3144_/S vssd1 vssd1 vccd1 vccd1 _2937_/A1 sky130_fd_sc_hd__buf_6
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3204_ _4402_/Q _4410_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4224_/A _4184_/B vssd1 vssd1 vccd1 vccd1 _4184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3135_ _4585_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__and3_1
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3066_ _3257_/A1 _3065_/X _3058_/X vssd1 vssd1 vccd1 vccd1 _3068_/B sky130_fd_sc_hd__o21a_4
XFILLER_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _2178_/Y _3941_/A _3967_/Y vssd1 vssd1 vccd1 vccd1 _4119_/B sky130_fd_sc_hd__o21ai_4
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2919_ _2971_/B _2918_/Y _2916_/Y vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__a21oi_2
X_3899_ _4161_/A _4127_/A _3899_/C _3899_/D vssd1 vssd1 vccd1 vccd1 _3899_/X sky130_fd_sc_hd__or4_2
XFILLER_100_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3822_ _3826_/A _3822_/B vssd1 vssd1 vccd1 vccd1 _4627_/D sky130_fd_sc_hd__or2_1
X_3753_ _3751_/B _3752_/Y _3761_/A vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__mux2_1
X_2704_ _4449_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2704_/X sky130_fd_sc_hd__and3_1
X_3684_ _4489_/Q _3762_/B _3691_/C _3683_/X vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__o31a_1
X_2635_ _2635_/A _2635_/B vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__or2_1
X_4305_ _4304_/X _3933_/B _4309_/S vssd1 vssd1 vccd1 vccd1 _4674_/D sky130_fd_sc_hd__mux2_1
X_2566_ _3288_/A _2566_/B vssd1 vssd1 vccd1 vccd1 _2566_/Y sky130_fd_sc_hd__nor2_1
X_2497_ _2661_/S _4541_/Q vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__and2b_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4236_ _3905_/A _4201_/X _4216_/B vssd1 vssd1 vccd1 vccd1 _4263_/S sky130_fd_sc_hd__a21oi_2
X_4167_ _4221_/A _4167_/B _4167_/C _4167_/D vssd1 vssd1 vccd1 vccd1 _4167_/X sky130_fd_sc_hd__or4_1
X_3118_ _3176_/A _3273_/B vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__or2_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _4119_/A _3894_/C _3899_/C vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ _3183_/A _3049_/B vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 _3256_/S vssd1 vssd1 vccd1 vccd1 _2645_/S sky130_fd_sc_hd__buf_8
X_2420_ _2418_/Y _2419_/X _3276_/B vssd1 vssd1 vccd1 vccd1 _2421_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2351_ _3581_/B _2351_/B _2351_/C _2352_/B vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__nor4_4
X_2282_ _2280_/X _2281_/X _2277_/X _4091_/B vssd1 vssd1 vccd1 vccd1 _2284_/B sky130_fd_sc_hd__o211ai_4
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4021_ _4017_/S _3401_/Y _3833_/X _3395_/B vssd1 vssd1 vccd1 vccd1 _4036_/S sky130_fd_sc_hd__a211o_4
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3805_ _2373_/B input1/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4615_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3736_ _3634_/Y _3734_/X _3735_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__o22a_1
X_3667_ _2432_/B _2591_/X _3666_/X _3384_/B vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__o22a_1
X_2618_ _3936_/A _2618_/B vssd1 vssd1 vccd1 vccd1 _2618_/Y sky130_fd_sc_hd__nor2_1
X_3598_ _3598_/A _3598_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__and3_1
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2549_ _2549_/A _2549_/B vssd1 vssd1 vccd1 vccd1 _2549_/Y sky130_fd_sc_hd__nand2_2
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4219_ _4248_/A _4213_/B _4261_/B _3585_/Y vssd1 vssd1 vccd1 vccd1 _4219_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout280 _3849_/A vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__buf_8
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4570_ _4570_/CLK _4570_/D vssd1 vssd1 vccd1 vccd1 _4570_/Q sky130_fd_sc_hd__dfxtp_1
X_3521_ _4534_/Q _3566_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4534_/D sky130_fd_sc_hd__mux2_1
X_3452_ _4473_/Q _3542_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4473_/D sky130_fd_sc_hd__mux2_1
X_3383_ _4631_/Q _3383_/B vssd1 vssd1 vccd1 vccd1 _3602_/B sky130_fd_sc_hd__nand2_2
X_2403_ _4508_/Q _4348_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _2404_/B sky130_fd_sc_hd__mux2_1
X_2334_ _2349_/B _2327_/Y _2612_/S _2332_/X vssd1 vssd1 vccd1 vccd1 _2337_/B sky130_fd_sc_hd__a211o_1
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2265_ _2268_/B vssd1 vssd1 vccd1 vccd1 _2265_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4004_ _2367_/Y _3834_/B _4003_/X _3397_/Y vssd1 vssd1 vccd1 vccd1 _4019_/S sky130_fd_sc_hd__o211a_4
X_2196_ _4662_/Q vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__inv_2
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4699_ _4700_/CLK _4699_/D vssd1 vssd1 vccd1 vccd1 _4699_/Q sky130_fd_sc_hd__dfxtp_1
X_3719_ _4685_/Q _3691_/C _3717_/Y _2331_/A vssd1 vssd1 vccd1 vccd1 _3719_/X sky130_fd_sc_hd__o22a_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _4668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2952_ _4381_/Q _4389_/Q _4405_/Q _4397_/Q _2950_/S _2893_/A vssd1 vssd1 vccd1 vccd1
+ _2953_/B sky130_fd_sc_hd__mux4_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _3209_/A _2940_/A _2882_/X _2377_/Y vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__o22a_1
X_4622_ _4674_/CLK _4622_/D vssd1 vssd1 vccd1 vccd1 _4622_/Q sky130_fd_sc_hd__dfxtp_1
X_4553_ _4553_/CLK _4553_/D vssd1 vssd1 vccd1 vccd1 _4553_/Q sky130_fd_sc_hd__dfxtp_1
X_3504_ _4519_/Q _3567_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4519_/D sky130_fd_sc_hd__mux2_1
X_4484_ _4551_/CLK _4484_/D vssd1 vssd1 vccd1 vccd1 _4484_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3435_ _4458_/Q _3570_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4458_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3366_ _4420_/Q _3564_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4420_/D sky130_fd_sc_hd__mux2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2284_/A _2284_/B _2284_/C _2315_/X vssd1 vssd1 vccd1 vccd1 _2335_/C sky130_fd_sc_hd__a31oi_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _4363_/Q _3580_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4363_/D sky130_fd_sc_hd__mux2_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _4643_/Q _2384_/B vssd1 vssd1 vccd1 vccd1 _2248_/Y sky130_fd_sc_hd__nand2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2179_ _4050_/A vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__inv_2
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput23 _4613_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_4
Xoutput34 _4672_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_4
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3220_ _4370_/Q _4699_/Q _4690_/Q _4418_/Q _3264_/S _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3220_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3151_ _4157_/B _4184_/B vssd1 vssd1 vccd1 vccd1 _3287_/C sky130_fd_sc_hd__and2_2
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3082_ _3239_/A _3130_/B _3082_/C vssd1 vssd1 vccd1 vccd1 _3082_/X sky130_fd_sc_hd__and3_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3984_ _3927_/A _3993_/C _3950_/X _2225_/Y vssd1 vssd1 vccd1 vccd1 _3985_/D sky130_fd_sc_hd__a22o_1
X_2935_ _4397_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2935_/X sky130_fd_sc_hd__and3_1
X_2866_ _2937_/A1 _2865_/X _2864_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__o211a_2
X_4605_ _4691_/CLK _4605_/D vssd1 vssd1 vccd1 vccd1 _4605_/Q sky130_fd_sc_hd__dfxtp_2
X_2797_ _4354_/Q _3570_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4354_/D sky130_fd_sc_hd__mux2_1
X_4536_ _4544_/CLK _4536_/D vssd1 vssd1 vccd1 vccd1 _4536_/Q sky130_fd_sc_hd__dfxtp_1
X_4467_ _4555_/CLK _4467_/D vssd1 vssd1 vccd1 vccd1 _4467_/Q sky130_fd_sc_hd__dfxtp_1
X_3418_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4443_/D sky130_fd_sc_hd__and2_1
X_4398_ _4678_/CLK _4398_/D vssd1 vssd1 vccd1 vccd1 _4398_/Q sky130_fd_sc_hd__dfxtp_1
X_3349_ _4405_/Q _4312_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4405_/D sky130_fd_sc_hd__mux2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _4577_/Q _4521_/Q _4513_/Q _4353_/Q _2824_/S _2404_/A vssd1 vssd1 vccd1 vccd1
+ _2720_/X sky130_fd_sc_hd__mux4_1
X_2651_ _3935_/A _2712_/B _2768_/B1 _2650_/Y vssd1 vssd1 vccd1 vccd1 _2685_/A sky130_fd_sc_hd__o211a_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2582_ _2937_/C1 _2579_/X _2581_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__a31o_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _4685_/Q _4332_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4685_/D sky130_fd_sc_hd__mux2_1
X_4252_ _4104_/A _4244_/Y _4246_/Y _2225_/Y _4251_/X vssd1 vssd1 vccd1 vccd1 _4252_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout109 _3201_/S vssd1 vssd1 vccd1 vccd1 _3254_/S sky130_fd_sc_hd__buf_6
X_3203_ _4394_/Q _4386_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__mux2_1
X_4183_ _3935_/A _4182_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4660_/D sky130_fd_sc_hd__mux2_1
X_3134_ _4681_/Q _4377_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3134_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3065_ _3061_/X _3064_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3065_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _4063_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _3967_/Y sky130_fd_sc_hd__nand2_2
X_2918_ _4684_/Q _2917_/B _2389_/A vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__a21oi_1
X_3898_ _3952_/A _3903_/A vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_30_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4626_/CLK sky130_fd_sc_hd__clkbuf_16
X_2849_ _2885_/A _2885_/B _2885_/C vssd1 vssd1 vccd1 vccd1 _2886_/A sky130_fd_sc_hd__and3_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4519_ _4543_/CLK _4519_/D vssd1 vssd1 vccd1 vccd1 _4519_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4665_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ _4627_/Q _4603_/Q _3827_/S vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3752_ _3770_/S _4184_/B _3751_/Y vssd1 vssd1 vccd1 vccd1 _3752_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_12_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2703_ _4465_/Q _4473_/Q _2809_/S vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__mux2_1
X_3683_ _3754_/A1 _3681_/Y _3682_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__o22a_1
X_2634_ _4352_/Q _4512_/Q _2636_/S vssd1 vssd1 vccd1 vccd1 _2635_/B sky130_fd_sc_hd__mux2_1
X_2565_ _3290_/A _2566_/B _2564_/X vssd1 vssd1 vccd1 vccd1 _2565_/Y sky130_fd_sc_hd__o21bai_1
X_4304_ _4062_/A _4303_/X _4241_/Y vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__a21bo_1
X_2496_ _4657_/Q _2495_/Y _2618_/B vssd1 vssd1 vccd1 vccd1 _2496_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4235_ _4235_/A _4235_/B _4265_/S vssd1 vssd1 vccd1 vccd1 _4238_/C sky130_fd_sc_hd__and3_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4166_ _4161_/Y _4162_/X _4165_/X _4159_/X vssd1 vssd1 vccd1 vccd1 _4167_/D sky130_fd_sc_hd__o211ai_1
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3117_ _3739_/A _3742_/B vssd1 vssd1 vccd1 vccd1 _3273_/B sky130_fd_sc_hd__nand2_1
X_4097_ _3972_/A _4096_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4657_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3048_ _3183_/A _3048_/B _3048_/C vssd1 vssd1 vccd1 vccd1 _3048_/X sky130_fd_sc_hd__or3_1
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout91 _3256_/S vssd1 vssd1 vccd1 vccd1 _3065_/S sky130_fd_sc_hd__buf_6
Xfanout80 _2847_/A1 vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ _2350_/A _2352_/B vssd1 vssd1 vccd1 vccd1 _2907_/A sky130_fd_sc_hd__nor2_4
XFILLER_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2281_ _4086_/A _4637_/Q _2178_/Y _2384_/B vssd1 vssd1 vccd1 vccd1 _2281_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4347_/A _4020_/B vssd1 vssd1 vccd1 vccd1 _4647_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4576_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _3836_/A _3804_/B vssd1 vssd1 vccd1 vccd1 _3812_/S sky130_fd_sc_hd__nor2_8
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3735_ _3739_/A _3734_/X _3771_/S vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__mux2_1
X_3666_ _2591_/X _3631_/X _3666_/B1 _3665_/X vssd1 vssd1 vccd1 vccd1 _3666_/X sky130_fd_sc_hd__o22a_1
X_3597_ _4625_/Q _4601_/Q vssd1 vssd1 vccd1 vccd1 _3598_/C sky130_fd_sc_hd__xnor2_1
X_2617_ _4061_/B _2617_/B _2617_/C _2617_/D vssd1 vssd1 vccd1 vccd1 _2817_/A sky130_fd_sc_hd__or4_4
X_2548_ _4550_/Q _4494_/Q _4486_/Q _4478_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2549_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _3855_/B _4267_/A2 _4267_/B1 _3934_/A vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__a22o_1
X_2479_ _4509_/Q _2636_/S _2478_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__a211o_1
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4149_ _4260_/B _4149_/B vssd1 vssd1 vccd1 vccd1 _4149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout281 input14/X vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__buf_6
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout270 _4003_/B vssd1 vssd1 vccd1 vccd1 _3384_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3520_ _4533_/Q _3565_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4533_/D sky130_fd_sc_hd__mux2_1
X_3451_ _4472_/Q _3541_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4472_/D sky130_fd_sc_hd__mux2_1
X_2402_ _4428_/Q _4420_/Q _4540_/Q _4532_/Q _2661_/S _2825_/B2 vssd1 vssd1 vccd1 vccd1
+ _2402_/X sky130_fd_sc_hd__mux4_1
X_3382_ _4435_/Q _3571_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4435_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2333_ _3629_/A _2333_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _3230_/A sky130_fd_sc_hd__or3_4
X_2264_ _3629_/A _2264_/B vssd1 vssd1 vccd1 vccd1 _2268_/B sky130_fd_sc_hd__xnor2_4
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2195_ _3836_/A vssd1 vssd1 vccd1 vccd1 _2195_/Y sky130_fd_sc_hd__inv_2
X_4003_ _4003_/A _4003_/B _4619_/Q vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__or3b_1
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4698_ _4698_/CLK _4698_/D vssd1 vssd1 vccd1 vccd1 _4698_/Q sky130_fd_sc_hd__dfxtp_1
X_3718_ _3716_/B _3717_/Y _3727_/S vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__mux2_1
X_3649_ _3643_/B _3749_/A1 _4329_/S vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__o21ba_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _2195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _2948_/X _2949_/X _2950_/X _2893_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2951_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4621_ _4674_/CLK _4621_/D vssd1 vssd1 vccd1 vccd1 _4621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2882_ _3966_/B _3259_/B _3160_/B1 _3288_/A vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__o211a_1
X_4552_ _4552_/CLK _4552_/D vssd1 vssd1 vccd1 vccd1 _4552_/Q sky130_fd_sc_hd__dfxtp_1
X_3503_ _4518_/Q _3566_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4518_/D sky130_fd_sc_hd__mux2_1
X_4483_ _4555_/CLK _4483_/D vssd1 vssd1 vccd1 vccd1 _4483_/Q sky130_fd_sc_hd__dfxtp_1
X_3434_ _4457_/Q _3569_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4457_/D sky130_fd_sc_hd__mux2_1
X_3365_ _3563_/B _4310_/A _4330_/C vssd1 vssd1 vccd1 vccd1 _3373_/S sky130_fd_sc_hd__and3_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _3836_/A _2316_/B _2316_/C vssd1 vssd1 vccd1 vccd1 _4436_/D sky130_fd_sc_hd__or3_1
XFILLER_85_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3291_/X _3293_/X _3295_/X vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__a21oi_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _3846_/A _4615_/Q vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__nand2_2
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2178_ _4643_/Q vssd1 vssd1 vccd1 vccd1 _2178_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput24 _4669_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_4
Xoutput35 _4673_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_4
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _3249_/C1 _3137_/X _3141_/X _3149_/X vssd1 vssd1 vccd1 vccd1 _4184_/B sky130_fd_sc_hd__o31ai_4
X_3081_ _4686_/Q _3080_/C _4687_/Q vssd1 vssd1 vccd1 vccd1 _3082_/C sky130_fd_sc_hd__o21ai_1
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3983_ _3980_/A _3980_/Y _4258_/B vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2934_ _4389_/Q _4381_/Q _2934_/S vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__mux2_1
X_2865_ _4676_/Q _4372_/Q _2932_/S vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__mux2_1
X_4604_ _4691_/CLK _4604_/D vssd1 vssd1 vccd1 vccd1 _4604_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4535_ _4543_/CLK _4535_/D vssd1 vssd1 vccd1 vccd1 _4535_/Q sky130_fd_sc_hd__dfxtp_1
X_2796_ _2854_/B _2795_/Y _2793_/Y vssd1 vssd1 vccd1 vccd1 _2796_/Y sky130_fd_sc_hd__a21oi_2
X_4466_ _4553_/CLK _4466_/D vssd1 vssd1 vccd1 vccd1 _4466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3417_ _4667_/Q _3416_/X _3417_/S vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__mux2_1
X_4397_ _4695_/CLK _4397_/D vssd1 vssd1 vccd1 vccd1 _4397_/Q sky130_fd_sc_hd__dfxtp_1
X_3348_ _4404_/Q _4331_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4404_/D sky130_fd_sc_hd__mux2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _4675_/Q _3278_/A _2425_/Y _3278_/Y vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__a211o_1
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ _2655_/B _2652_/B _2618_/B vssd1 vssd1 vccd1 vccd1 _2650_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2581_ _4575_/Q _2932_/S _2580_/X _2937_/A1 vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__a211o_1
X_4320_ _4684_/Q _4320_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4684_/D sky130_fd_sc_hd__mux2_1
X_4251_ _4215_/A _4264_/A _4247_/X _4250_/X vssd1 vssd1 vccd1 vccd1 _4251_/X sky130_fd_sc_hd__a31o_1
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3202_ _3200_/X _3201_/X _3252_/S vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__mux2_1
X_4182_ _4240_/A _4170_/Y _4181_/X _4270_/B input8/X vssd1 vssd1 vccd1 vccd1 _4182_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3133_ _4360_/Q _3577_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4360_/D sky130_fd_sc_hd__mux2_1
X_3064_ _3062_/X _3063_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _4643_/Q _3966_/B vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__xnor2_2
X_2917_ _4684_/Q _2917_/B vssd1 vssd1 vccd1 vccd1 _2971_/B sky130_fd_sc_hd__or2_2
X_3897_ _3952_/A _3903_/A vssd1 vssd1 vccd1 vccd1 _4213_/B sky130_fd_sc_hd__nor2_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2848_ _2848_/A _2848_/B _2848_/C vssd1 vssd1 vccd1 vccd1 _2885_/C sky130_fd_sc_hd__and3_1
X_2779_ _2898_/A _2777_/X _2774_/X vssd1 vssd1 vccd1 vccd1 _3690_/B sky130_fd_sc_hd__o21ai_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4518_ _4574_/CLK _4518_/D vssd1 vssd1 vccd1 vccd1 _4518_/Q sky130_fd_sc_hd__dfxtp_1
X_4449_ _4555_/CLK _4449_/D vssd1 vssd1 vccd1 vccd1 _4449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _3826_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _4626_/D sky130_fd_sc_hd__or2_1
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3751_ _3770_/S _3751_/B vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__nand2_1
X_2702_ _2644_/S _2699_/X _2701_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2702_/X sky130_fd_sc_hd__o211a_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3682_ _3680_/B _3681_/Y _3727_/S vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__mux2_1
X_2633_ _2631_/X _2632_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__mux2_1
X_2564_ _2377_/Y _2541_/Y _2563_/Y _2847_/A1 _2746_/A1 vssd1 vssd1 vccd1 vccd1 _2564_/X
+ sky130_fd_sc_hd__a221o_1
X_4303_ _4662_/Q _4278_/Y _4302_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4303_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2495_ _2655_/B _2517_/S vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__xnor2_1
X_4234_ _3956_/A _4233_/B _4216_/B vssd1 vssd1 vccd1 vccd1 _4265_/S sky130_fd_sc_hd__a21o_1
X_4165_ _3886_/X _3961_/Y _4188_/C _3993_/A _4086_/A vssd1 vssd1 vccd1 vccd1 _4165_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _3041_/Y _3742_/B _3174_/A vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4096_ _4240_/A _4081_/Y _4095_/X _4270_/B input5/X vssd1 vssd1 vccd1 vccd1 _4096_/X
+ sky130_fd_sc_hd__a32o_1
X_3047_ _3770_/S _3739_/A _3046_/Y _3020_/S vssd1 vssd1 vccd1 vccd1 _3048_/C sky130_fd_sc_hd__o211a_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3949_ _4261_/B _4261_/C _4261_/A vssd1 vssd1 vccd1 vccd1 _4262_/B sky130_fd_sc_hd__a21oi_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout92 _2444_/X vssd1 vssd1 vccd1 vccd1 _3256_/S sky130_fd_sc_hd__buf_8
Xfanout70 _4330_/A vssd1 vssd1 vccd1 vccd1 _4310_/B sky130_fd_sc_hd__clkbuf_4
Xfanout81 _2353_/X vssd1 vssd1 vccd1 vccd1 _2847_/A1 sky130_fd_sc_hd__buf_8
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2280_ _2244_/X _2245_/X _3585_/B vssd1 vssd1 vccd1 vccd1 _2280_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3803_ _4692_/Q _4042_/C _4042_/A vssd1 vssd1 vccd1 vccd1 _3804_/B sky130_fd_sc_hd__or3b_4
X_3734_ _3739_/A _3068_/B _3760_/A vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__mux2_1
X_3665_ _4487_/Q _3762_/B _4013_/S _3664_/X vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__o31a_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2616_ _4061_/B _2617_/B _2617_/C _2617_/D vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__o31a_1
X_3596_ _2181_/Y _4606_/Q _4623_/Q _2186_/Y _3591_/Y vssd1 vssd1 vccd1 vccd1 _3598_/B
+ sky130_fd_sc_hd__o221a_1
X_2547_ _2544_/X _2545_/X _2546_/X _2829_/S1 _2549_/A vssd1 vssd1 vccd1 vccd1 _2547_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2478_ _4349_/Q _2798_/B _2798_/C vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__and3_1
X_4217_ _4217_/A _4233_/A vssd1 vssd1 vccd1 vccd1 _4217_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4148_ _3912_/X _3913_/Y _3916_/A _3921_/X vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__a211o_1
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4079_ _2995_/A _4078_/X _4224_/A vssd1 vssd1 vccd1 vccd1 _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout271 _4003_/B vssd1 vssd1 vccd1 vccd1 _2354_/A sky130_fd_sc_hd__clkbuf_4
Xfanout282 input14/X vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__clkbuf_16
Xfanout260 _2598_/S vssd1 vssd1 vccd1 vccd1 _2546_/S sky130_fd_sc_hd__buf_8
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _4471_/Q _3540_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4471_/D sky130_fd_sc_hd__mux2_1
X_3381_ _4434_/Q _3570_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4434_/D sky130_fd_sc_hd__mux2_1
X_2401_ _3572_/A _3563_/A _3563_/B vssd1 vssd1 vccd1 vccd1 _2857_/S sky130_fd_sc_hd__and3_4
X_2332_ _3930_/A _3990_/A _2384_/D vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__and3_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2263_ _2263_/A _2263_/B _2263_/C _2263_/D vssd1 vssd1 vccd1 vccd1 _2264_/B sky130_fd_sc_hd__or4_4
X_4002_ _2178_/Y _3992_/X _4001_/Y _3849_/A vssd1 vssd1 vccd1 vccd1 _4643_/D sky130_fd_sc_hd__a211oi_1
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2194_ _3689_/A vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3717_ _3716_/A _2995_/A _3716_/Y vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__o21ai_1
X_4697_ _4697_/CLK _4697_/D vssd1 vssd1 vccd1 vccd1 _4697_/Q sky130_fd_sc_hd__dfxtp_1
X_3648_ _2617_/B _3747_/B2 _3666_/B1 _3647_/X vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3579_ _4586_/Q _4317_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4586_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2950_ _4373_/Q _4677_/Q _2950_/S vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _3257_/A1 _2875_/X _2879_/X _2866_/X _2871_/X vssd1 vssd1 vccd1 vccd1 _2940_/A
+ sky130_fd_sc_hd__o32ai_4
X_4620_ _4674_/CLK _4620_/D vssd1 vssd1 vccd1 vccd1 _4620_/Q sky130_fd_sc_hd__dfxtp_2
X_4551_ _4551_/CLK _4551_/D vssd1 vssd1 vccd1 vccd1 _4551_/Q sky130_fd_sc_hd__dfxtp_1
X_3502_ _4517_/Q _3565_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4517_/D sky130_fd_sc_hd__mux2_1
X_4482_ _4490_/CLK _4482_/D vssd1 vssd1 vccd1 vccd1 _4482_/Q sky130_fd_sc_hd__dfxtp_1
X_3433_ _4456_/Q _3541_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4456_/D sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _4419_/Q _4338_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4419_/D sky130_fd_sc_hd__mux2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2366_/B _2261_/B _2230_/B vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__a21o_1
X_3295_ _4691_/Q _3239_/B _3294_/Y vssd1 vssd1 vccd1 vccd1 _3295_/X sky130_fd_sc_hd__o21a_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _3846_/A _4615_/Q vssd1 vssd1 vccd1 vccd1 _2384_/B sky130_fd_sc_hd__and2_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2177_ _4646_/Q vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput25 _4614_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_4
Xoutput36 _4674_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_4
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _4686_/Q _4687_/Q _3080_/C vssd1 vssd1 vccd1 vccd1 _3130_/B sky130_fd_sc_hd__or3_1
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3982_ _3927_/A _4086_/A _2366_/B vssd1 vssd1 vccd1 vccd1 _4228_/B sky130_fd_sc_hd__o21ai_4
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2933_ _2937_/A1 _2932_/X _2931_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2933_/X sky130_fd_sc_hd__o211a_2
X_2864_ _4356_/Q _2932_/S _2863_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__a211o_1
X_4603_ _4700_/CLK _4603_/D vssd1 vssd1 vccd1 vccd1 _4603_/Q sky130_fd_sc_hd__dfxtp_2
X_2795_ _4490_/Q _2794_/B _2571_/A vssd1 vssd1 vccd1 vccd1 _2795_/Y sky130_fd_sc_hd__a21oi_1
X_4534_ _4574_/CLK _4534_/D vssd1 vssd1 vccd1 vccd1 _4534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ _4481_/CLK _4465_/D vssd1 vssd1 vccd1 vccd1 _4465_/Q sky130_fd_sc_hd__dfxtp_1
X_3416_ _4671_/Q _4081_/A _3415_/Y vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__o21a_1
X_4396_ _4584_/CLK _4396_/D vssd1 vssd1 vccd1 vccd1 _4396_/Q sky130_fd_sc_hd__dfxtp_1
X_3347_ _4319_/A _4310_/B _3446_/C vssd1 vssd1 vccd1 vccd1 _3355_/S sky130_fd_sc_hd__and3_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3278_/A _3278_/B vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__nor2_1
X_2229_ _2373_/C _2230_/B vssd1 vssd1 vccd1 vccd1 _3581_/D sky130_fd_sc_hd__nor2_4
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2580_ _4519_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__and3_1
X_4250_ _4662_/Q _4267_/B1 _4221_/A _4249_/X vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__a211o_1
X_4181_ _4181_/A _4181_/B _4181_/C _4181_/D vssd1 vssd1 vccd1 vccd1 _4181_/X sky130_fd_sc_hd__or4_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3201_ _4699_/Q _4370_/Q _3201_/S vssd1 vssd1 vccd1 vccd1 _3201_/X sky130_fd_sc_hd__mux2_1
X_3132_ _3237_/C _3131_/Y _3129_/X vssd1 vssd1 vccd1 vccd1 _3132_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _4399_/Q _4407_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _3972_/A _4116_/A vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__or2_2
X_3896_ _3896_/A _3896_/B vssd1 vssd1 vccd1 vccd1 _4244_/B sky130_fd_sc_hd__nand2_2
X_2916_ _2916_/A _2916_/B vssd1 vssd1 vccd1 vccd1 _2916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ _2847_/A1 _2846_/X _3239_/A vssd1 vssd1 vccd1 vccd1 _2847_/Y sky130_fd_sc_hd__a21oi_1
X_2778_ _2898_/A _2777_/X _2774_/X vssd1 vssd1 vccd1 vccd1 _3689_/B sky130_fd_sc_hd__o21a_4
X_4517_ _4573_/CLK _4517_/D vssd1 vssd1 vccd1 vccd1 _4517_/Q sky130_fd_sc_hd__dfxtp_1
X_4448_ _4552_/CLK _4448_/D vssd1 vssd1 vccd1 vccd1 _4448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4379_ _4683_/CLK _4379_/D vssd1 vssd1 vccd1 vccd1 _4379_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3750_ _4603_/Q _3741_/S _3749_/X vssd1 vssd1 vccd1 vccd1 _4603_/D sky130_fd_sc_hd__a21bo_1
X_2701_ _4489_/Q _2699_/S _2700_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__a211o_1
X_3681_ _3689_/A _2848_/A _3680_/Y vssd1 vssd1 vccd1 vccd1 _3681_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2632_ _4424_/Q _4432_/Q _2636_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
X_2563_ _2846_/S _2555_/X _2561_/X _2562_/Y vssd1 vssd1 vccd1 vccd1 _2563_/Y sky130_fd_sc_hd__o22ai_4
X_4302_ _4646_/Q _2367_/Y _3629_/Y _4654_/Q vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__a22o_1
X_4233_ _4233_/A _4233_/B vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__nand2_1
X_2494_ _2541_/A _2540_/A vssd1 vssd1 vccd1 vccd1 _2517_/S sky130_fd_sc_hd__nand2b_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _3585_/Y _4205_/B _4161_/A _2371_/C vssd1 vssd1 vccd1 vccd1 _4167_/C sky130_fd_sc_hd__a2bb2o_1
X_4095_ _4123_/A _4095_/B _4095_/C _4095_/D vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__or4_1
X_3115_ _3109_/X _3111_/X _3114_/X _3270_/A vssd1 vssd1 vccd1 vccd1 _3742_/B sky130_fd_sc_hd__o22a_4
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3770_/S _3049_/B vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _4212_/B _3947_/X _4213_/B vssd1 vssd1 vccd1 vccd1 _4261_/C sky130_fd_sc_hd__a21o_1
X_3879_ _4063_/A _3941_/A vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout82 _2466_/X vssd1 vssd1 vccd1 vccd1 _4061_/B sky130_fd_sc_hd__buf_4
Xfanout60 _2688_/X vssd1 vssd1 vccd1 vccd1 _3568_/A1 sky130_fd_sc_hd__buf_6
Xfanout71 _2861_/X vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__clkbuf_4
Xfanout93 _3194_/C1 vssd1 vssd1 vccd1 vccd1 _2933_/C1 sky130_fd_sc_hd__buf_8
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3802_ _3802_/A _3802_/B vssd1 vssd1 vccd1 vccd1 _4042_/C sky130_fd_sc_hd__or2_1
X_3733_ _4601_/Q _3741_/S _3732_/Y vssd1 vssd1 vccd1 vccd1 _4601_/D sky130_fd_sc_hd__a21o_1
X_3664_ _3754_/A1 _3662_/X _3663_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _3664_/X sky130_fd_sc_hd__o22a_1
X_2615_ _2611_/X _2614_/X _2846_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
X_3595_ _4628_/Q _2184_/Y _2185_/Y _4599_/Q _3594_/Y vssd1 vssd1 vccd1 vccd1 _3595_/X
+ sky130_fd_sc_hd__o221a_1
X_2546_ _4430_/Q _4422_/Q _2546_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_2
X_2477_ _2805_/C1 _2476_/X _2475_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__o211a_2
X_4216_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__or2_1
X_4147_ _3872_/Y _3938_/Y _4114_/B _4146_/Y vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__a31o_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4248_/A _4092_/A _4103_/B _3585_/Y _4077_/Y vssd1 vssd1 vccd1 vccd1 _4078_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _3216_/S _4583_/Q _3266_/A1 vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__a21bo_1
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout250 _2776_/S1 vssd1 vssd1 vccd1 vccd1 _2775_/S1 sky130_fd_sc_hd__buf_4
Xfanout272 _4003_/B vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__buf_4
Xfanout261 _2598_/S vssd1 vssd1 vccd1 vccd1 _2775_/S0 sky130_fd_sc_hd__buf_6
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2400_ _3826_/A _2400_/B _2400_/C _2861_/B vssd1 vssd1 vccd1 vccd1 _2400_/X sky130_fd_sc_hd__or4_4
X_3380_ _4433_/Q _3569_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4433_/D sky130_fd_sc_hd__mux2_1
X_2331_ _2331_/A _2372_/C vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__or2_4
X_2262_ _3846_/B _3993_/B vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__nand2_4
X_4001_ _4238_/A _3993_/X _4000_/X _3986_/X _3992_/X vssd1 vssd1 vccd1 vccd1 _4001_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2193_ _4056_/B vssd1 vssd1 vccd1 vccd1 _3846_/B sky130_fd_sc_hd__clkinv_4
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3716_ _3716_/A _3716_/B vssd1 vssd1 vccd1 vccd1 _3716_/Y sky130_fd_sc_hd__nand2_1
X_4696_ _4696_/CLK _4696_/D vssd1 vssd1 vccd1 vccd1 _4696_/Q sky130_fd_sc_hd__dfxtp_1
X_3647_ _4485_/Q _3407_/B _4013_/S _3646_/X vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__o31a_1
X_3578_ _4585_/Q _4336_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4585_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2529_ _2814_/A1 _2526_/X _2528_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__o211a_2
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2880_ _3257_/A1 _2875_/X _2879_/X _2866_/X _2871_/X vssd1 vssd1 vccd1 vccd1 _2996_/A
+ sky130_fd_sc_hd__o32a_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4551_/CLK _4550_/D vssd1 vssd1 vccd1 vccd1 _4550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3501_ _4516_/Q _3564_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4516_/D sky130_fd_sc_hd__mux2_1
X_4481_ _4481_/CLK _4481_/D vssd1 vssd1 vccd1 vccd1 _4481_/Q sky130_fd_sc_hd__dfxtp_1
X_3432_ _4455_/Q _3567_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4455_/D sky130_fd_sc_hd__mux2_1
X_3363_ _4418_/Q _4337_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4418_/D sky130_fd_sc_hd__mux2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _4042_/A _2286_/C _3581_/D _2284_/X _2313_/X vssd1 vssd1 vccd1 vccd1 _2316_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3294_ _4691_/Q _3239_/B _2389_/A vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__a21oi_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _3917_/A _3941_/A _3936_/A _3938_/A vssd1 vssd1 vccd1 vccd1 _2245_/X sky130_fd_sc_hd__or4_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2176_ _4647_/Q vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4679_ _4679_/CLK _4679_/D vssd1 vssd1 vccd1 vccd1 _4679_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput15 _4708_/A vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_4
Xoutput26 _4637_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_4
Xoutput37 _4675_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3981_ _3927_/A _4086_/A _2366_/B vssd1 vssd1 vccd1 vccd1 _4084_/A sky130_fd_sc_hd__o21a_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ _4694_/Q _4365_/Q _2932_/S vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4584_/CLK sky130_fd_sc_hd__clkbuf_16
X_2863_ _4580_/Q _2863_/B _2863_/C vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__and3_1
X_4602_ _4691_/CLK _4602_/D vssd1 vssd1 vccd1 vccd1 _4602_/Q sky130_fd_sc_hd__dfxtp_1
X_2794_ _4490_/Q _2794_/B vssd1 vssd1 vccd1 vccd1 _2854_/B sky130_fd_sc_hd__or2_2
X_4533_ _4544_/CLK _4533_/D vssd1 vssd1 vccd1 vccd1 _4533_/Q sky130_fd_sc_hd__dfxtp_1
X_4464_ _4464_/CLK _4464_/D vssd1 vssd1 vccd1 vccd1 _4464_/Q sky130_fd_sc_hd__dfxtp_1
X_3415_ _3629_/A _4081_/A _3405_/A vssd1 vssd1 vccd1 vccd1 _3415_/Y sky130_fd_sc_hd__a21oi_1
X_4395_ _4587_/CLK _4395_/D vssd1 vssd1 vccd1 vccd1 _4395_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _4403_/Q _3580_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4403_/D sky130_fd_sc_hd__mux2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3041_/A _3274_/Y _3275_/X _3174_/A _3276_/X vssd1 vssd1 vccd1 vccd1 _3278_/B
+ sky130_fd_sc_hd__o221a_1
X_2228_ _3629_/A _2261_/B vssd1 vssd1 vccd1 vccd1 _2230_/B sky130_fd_sc_hd__nor2_4
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4700_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4643_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4180_ _3910_/X _4141_/Y _4202_/B _4264_/B vssd1 vssd1 vccd1 vccd1 _4181_/D sky130_fd_sc_hd__o211a_1
X_3200_ _4418_/Q _4690_/Q _3201_/S vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__mux2_1
X_3131_ _4688_/Q _3130_/B _2389_/A vssd1 vssd1 vccd1 vccd1 _3131_/Y sky130_fd_sc_hd__a21oi_1
X_3062_ _4391_/Q _4383_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _3964_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_15_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4464_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3895_ _3896_/A _3896_/B vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__and2_4
X_2915_ _3966_/B _2860_/C _3239_/A _2887_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _2916_/B
+ sky130_fd_sc_hd__a2111o_1
X_2846_ _2841_/X _2845_/X _2846_/S vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__mux2_1
X_2777_ _2775_/X _2776_/X _3036_/S vssd1 vssd1 vccd1 vccd1 _2777_/X sky130_fd_sc_hd__mux2_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4516_ _4572_/CLK _4516_/D vssd1 vssd1 vccd1 vccd1 _4516_/Q sky130_fd_sc_hd__dfxtp_1
X_4447_ _4667_/CLK _4447_/D vssd1 vssd1 vccd1 vccd1 _4447_/Q sky130_fd_sc_hd__dfxtp_1
X_4378_ _4682_/CLK _4378_/D vssd1 vssd1 vccd1 vccd1 _4378_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _4310_/B _3446_/C _4330_/C vssd1 vssd1 vccd1 vccd1 _3337_/S sky130_fd_sc_hd__and3_4
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2700_ _4481_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__and3_1
X_3680_ _3689_/A _3680_/B vssd1 vssd1 vccd1 vccd1 _3680_/Y sky130_fd_sc_hd__nand2_1
X_2631_ _4536_/Q _4544_/Q _2636_/S vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__mux2_1
X_2562_ _3938_/B _2345_/Y _3280_/B1 vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4301_ _4300_/X _4673_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4673_/D sky130_fd_sc_hd__mux2_1
X_4232_ _3927_/A _3927_/B _3925_/Y _4231_/X _4230_/X vssd1 vssd1 vccd1 vccd1 _4232_/X
+ sky130_fd_sc_hd__o41a_1
X_2493_ _4061_/B _2617_/B vssd1 vssd1 vccd1 vccd1 _2540_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_4_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4555_/CLK sky130_fd_sc_hd__clkbuf_16
X_4163_ _3934_/A _4267_/A2 _4267_/B1 _3936_/A vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__a22o_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4094_ _4084_/B _4235_/A _4092_/Y _4229_/A _4093_/X vssd1 vssd1 vccd1 vccd1 _4095_/D
+ sky130_fd_sc_hd__a221o_1
X_3114_ _3112_/X _3113_/X _3261_/A vssd1 vssd1 vccd1 vccd1 _3114_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3045_ _4671_/Q _3232_/S _3280_/B1 _3044_/Y vssd1 vssd1 vccd1 vccd1 _3048_/B sky130_fd_sc_hd__o211a_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3947_ _4205_/B _4205_/C _4205_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _3972_/A _4082_/A vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__nand2b_2
X_2829_ _4475_/Q _4467_/Q _4459_/Q _4451_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2829_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout61 _2688_/X vssd1 vssd1 vccd1 vccd1 _3541_/A1 sky130_fd_sc_hd__buf_2
Xfanout50 _4332_/A1 vssd1 vssd1 vccd1 vccd1 _4312_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout72 _2400_/X vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__buf_4
Xfanout83 _2365_/X vssd1 vssd1 vccd1 vccd1 _3160_/B1 sky130_fd_sc_hd__buf_6
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout94 _3194_/C1 vssd1 vssd1 vccd1 vccd1 _2814_/C1 sky130_fd_sc_hd__buf_6
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ _3619_/B _3799_/X _3800_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3732_ _3749_/A1 _3730_/X _3731_/X vssd1 vssd1 vccd1 vccd1 _3732_/Y sky130_fd_sc_hd__a21oi_2
X_3663_ _2669_/C _3662_/X _3771_/S vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__mux2_1
X_2614_ _4671_/Q _2613_/X _2614_/S vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__mux2_1
X_3594_ _4626_/Q _4602_/Q vssd1 vssd1 vccd1 vccd1 _3594_/Y sky130_fd_sc_hd__xnor2_1
X_2545_ _2546_/S _4534_/Q _2829_/S1 vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__a21bo_1
X_2476_ _4421_/Q _4429_/Q _2636_/S vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__mux2_1
X_4215_ _4215_/A _4215_/B _4247_/S vssd1 vssd1 vccd1 vccd1 _4221_/C sky130_fd_sc_hd__and3_1
X_4146_ _4229_/A _4177_/C vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4077_ _4104_/A _3883_/X _4072_/Y _4076_/X _4071_/X vssd1 vssd1 vccd1 vccd1 _4077_/Y
+ sky130_fd_sc_hd__a311oi_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3028_ _3216_/S _4359_/Q vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__and2b_1
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout240 _3270_/A vssd1 vssd1 vccd1 vccd1 _2668_/A1 sky130_fd_sc_hd__buf_8
Xfanout273 _4003_/B vssd1 vssd1 vccd1 vccd1 _3383_/B sky130_fd_sc_hd__buf_2
Xfanout251 _4441_/Q vssd1 vssd1 vccd1 vccd1 _2776_/S1 sky130_fd_sc_hd__buf_4
Xfanout262 _2823_/A1 vssd1 vssd1 vccd1 vccd1 _2598_/S sky130_fd_sc_hd__buf_6
XFILLER_75_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ _2331_/A _2372_/C vssd1 vssd1 vccd1 vccd1 _2330_/Y sky130_fd_sc_hd__nor2_2
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2261_ _2366_/B _2261_/B vssd1 vssd1 vccd1 vccd1 _2300_/A sky130_fd_sc_hd__nor2_2
X_4000_ _3855_/B _3857_/B _2261_/B _2373_/C _4246_/A vssd1 vssd1 vccd1 vccd1 _4000_/X
+ sky130_fd_sc_hd__a221o_1
X_2192_ _2373_/B vssd1 vssd1 vccd1 vccd1 _2368_/A sky130_fd_sc_hd__clkinv_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _3713_/Y _3714_/X _4599_/Q _3741_/S vssd1 vssd1 vccd1 vccd1 _4599_/D sky130_fd_sc_hd__a2bb2o_1
X_4695_ _4695_/CLK _4695_/D vssd1 vssd1 vccd1 vccd1 _4695_/Q sky130_fd_sc_hd__dfxtp_1
X_3646_ _3754_/A1 _3644_/Y _3645_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__o22a_1
X_3577_ _4584_/Q _3577_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4584_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2528_ _4542_/Q _2809_/S _2527_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2528_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2459_ _4484_/Q _2811_/S _2456_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__a211o_1
X_4129_ _3885_/Y _4140_/A _3886_/X _4104_/A vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__o211a_1
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3500_ _3563_/A _3563_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _3508_/S sky130_fd_sc_hd__and3_4
X_4480_ _4552_/CLK _4480_/D vssd1 vssd1 vccd1 vccd1 _4480_/Q sky130_fd_sc_hd__dfxtp_1
X_3431_ _4454_/Q _3539_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4454_/D sky130_fd_sc_hd__mux2_1
X_3362_ _4417_/Q _4336_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4417_/D sky130_fd_sc_hd__mux2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2233_/C _3601_/B _4050_/A vssd1 vssd1 vccd1 vccd1 _2313_/X sky130_fd_sc_hd__o21a_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _2385_/Y _3290_/X _3292_/X _2389_/A vssd1 vssd1 vccd1 vccd1 _3293_/X sky130_fd_sc_hd__o31a_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _3934_/A _3935_/A _3259_/A _4662_/Q vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__or4_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4678_ _4678_/CLK _4678_/D vssd1 vssd1 vccd1 vccd1 _4678_/Q sky130_fd_sc_hd__dfxtp_1
X_3629_ _3629_/A _3629_/B vssd1 vssd1 vccd1 vccd1 _3629_/Y sky130_fd_sc_hd__nor2_4
Xoutput27 _4635_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_4
Xoutput16 _4668_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ _3980_/A _4266_/A vssd1 vssd1 vccd1 vccd1 _3980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2931_ _4685_/Q _2932_/S _2930_/X _2931_/C1 vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2862_ _4319_/A _4310_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _3297_/S sky130_fd_sc_hd__and3_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4601_ _4691_/CLK _4601_/D vssd1 vssd1 vccd1 vccd1 _4601_/Q sky130_fd_sc_hd__dfxtp_2
X_2793_ _2793_/A _2793_/B vssd1 vssd1 vccd1 vccd1 _2793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4576_/CLK _4532_/D vssd1 vssd1 vccd1 vccd1 _4532_/Q sky130_fd_sc_hd__dfxtp_1
X_4463_ _4667_/CLK _4463_/D vssd1 vssd1 vccd1 vccd1 _4463_/Q sky130_fd_sc_hd__dfxtp_1
X_3414_ _4347_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _4442_/D sky130_fd_sc_hd__and2_1
X_4394_ _4587_/CLK _4394_/D vssd1 vssd1 vccd1 vccd1 _4394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _4402_/Q _4337_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4402_/D sky130_fd_sc_hd__mux2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _4618_/Q _3276_/B _3276_/C vssd1 vssd1 vccd1 vccd1 _3276_/X sky130_fd_sc_hd__or3_1
X_2227_ _3930_/A _4262_/A _3581_/C _2349_/B _2217_/B vssd1 vssd1 vccd1 vccd1 _2286_/C
+ sky130_fd_sc_hd__o2111a_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3130_ _4688_/Q _3130_/B vssd1 vssd1 vccd1 vccd1 _3237_/C sky130_fd_sc_hd__or2_2
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3061_ _3059_/X _3060_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _4127_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__and2_2
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3894_ _3894_/A _4072_/A _3894_/C vssd1 vssd1 vccd1 vccd1 _3899_/D sky130_fd_sc_hd__or3_1
X_2914_ _3183_/A _2912_/X _2913_/Y _3282_/A vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__o211a_1
X_2845_ _2422_/A _2843_/X _2844_/Y _2614_/S _3857_/B vssd1 vssd1 vccd1 vccd1 _2845_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4515_ _4579_/CLK _4515_/D vssd1 vssd1 vccd1 vccd1 _4515_/Q sky130_fd_sc_hd__dfxtp_1
X_2776_ _4554_/Q _4498_/Q _4490_/Q _4482_/Q _2598_/S _2776_/S1 vssd1 vssd1 vccd1 vccd1
+ _2776_/X sky130_fd_sc_hd__mux4_1
X_4446_ _4481_/CLK _4446_/D vssd1 vssd1 vccd1 vccd1 _4446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4377_ _4681_/CLK _4377_/D vssd1 vssd1 vccd1 vccd1 _4377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3328_/A _3328_/B vssd1 vssd1 vccd1 vccd1 _4330_/C sky130_fd_sc_hd__nor2_8
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3259_ _3259_/A _3259_/B vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _4351_/Q _3567_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4351_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2561_ _3041_/A _2554_/Y _2560_/X _2345_/Y vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__o211a_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4300_ input9/X _4299_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4300_/X sky130_fd_sc_hd__mux2_1
X_2492_ _4061_/B _2617_/B vssd1 vssd1 vccd1 vccd1 _2541_/A sky130_fd_sc_hd__nor2_1
X_4231_ _3904_/Y _3905_/X _3908_/A _3924_/X vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__o211a_1
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4162_ _4161_/A _4161_/B _3927_/B vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__a21o_1
X_4093_ _4260_/B _4264_/B _4093_/S vssd1 vssd1 vccd1 vccd1 _4093_/X sky130_fd_sc_hd__mux2_1
X_3113_ _4384_/Q _4392_/Q _4408_/Q _4400_/Q _3163_/S _3113_/S1 vssd1 vssd1 vccd1 vccd1
+ _3113_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _3232_/S _3044_/B vssd1 vssd1 vccd1 vccd1 _3044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ _4177_/B _4177_/C _4177_/A vssd1 vssd1 vccd1 vccd1 _4205_/C sky130_fd_sc_hd__a21o_1
X_3877_ _3964_/B _4132_/A vssd1 vssd1 vccd1 vccd1 _3877_/Y sky130_fd_sc_hd__nand2_1
X_2828_ _4555_/Q _4499_/Q _4491_/Q _4483_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2828_/X sky130_fd_sc_hd__mux4_1
X_2759_ _4490_/Q _2811_/S _2758_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__a211o_1
X_4429_ _4544_/CLK _4429_/D vssd1 vssd1 vccd1 vccd1 _4429_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout40 _4337_/A1 vssd1 vssd1 vccd1 vccd1 _4317_/A1 sky130_fd_sc_hd__buf_4
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout51 _2973_/Y vssd1 vssd1 vccd1 vccd1 _4332_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout62 _2629_/X vssd1 vssd1 vccd1 vccd1 _3567_/A1 sky130_fd_sc_hd__buf_4
Xfanout73 _2400_/X vssd1 vssd1 vccd1 vccd1 _3536_/A sky130_fd_sc_hd__clkbuf_2
Xfanout95 _2443_/X vssd1 vssd1 vccd1 vccd1 _3194_/C1 sky130_fd_sc_hd__clkbuf_16
Xfanout84 _2365_/X vssd1 vssd1 vccd1 vccd1 _2768_/B1 sky130_fd_sc_hd__buf_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3800_ _4614_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3800_/X sky130_fd_sc_hd__or2_1
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3731_ _3731_/A1 _3072_/B _3119_/B _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3731_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3662_ _2591_/X _2669_/C _3689_/A vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2613_ _2610_/Y _2612_/X _3041_/A vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__mux2_1
X_3593_ _4630_/Q _2182_/Y _2183_/Y _4604_/Q _3592_/Y vssd1 vssd1 vccd1 vccd1 _3593_/X
+ sky130_fd_sc_hd__o221a_1
X_2544_ _2546_/S _4542_/Q vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__and2b_1
X_2475_ _4541_/Q _2636_/S _2474_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__a211o_1
X_4214_ _4213_/B _4213_/A _3904_/Y vssd1 vssd1 vccd1 vccd1 _4247_/S sky130_fd_sc_hd__a21oi_1
X_4145_ _4266_/B _4139_/X _4140_/Y _4144_/X vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__o31a_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _4215_/A _3894_/C _4074_/Y _4075_/X vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__a31o_1
X_3027_ _4358_/Q _4313_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4358_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3929_ _3896_/A _3926_/X _3928_/Y vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout230 _4618_/Q vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__buf_8
Xfanout241 _4443_/Q vssd1 vssd1 vccd1 vccd1 _3270_/A sky130_fd_sc_hd__buf_12
Xfanout274 _3405_/A vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__buf_8
Xfanout263 _4440_/Q vssd1 vssd1 vccd1 vccd1 _2823_/A1 sky130_fd_sc_hd__buf_4
Xfanout252 _3165_/S1 vssd1 vssd1 vccd1 vccd1 _3113_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2260_ _4248_/A vssd1 vssd1 vccd1 vccd1 _2371_/C sky130_fd_sc_hd__inv_2
X_2191_ _2292_/B vssd1 vssd1 vccd1 vccd1 _2360_/A sky130_fd_sc_hd__inv_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4694_ _4694_/CLK _4694_/D vssd1 vssd1 vccd1 vccd1 _4694_/Q sky130_fd_sc_hd__dfxtp_1
X_3714_ _3731_/A1 _2940_/A _3013_/B _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3714_/X
+ sky130_fd_sc_hd__a221o_2
X_3645_ _3643_/B _3644_/Y _3771_/S vssd1 vssd1 vccd1 vccd1 _3645_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3576_ _4583_/Q _4314_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4583_/D sky130_fd_sc_hd__mux2_1
X_2527_ _4534_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__and3_1
X_2458_ _4548_/Q _2809_/S _2457_/X _2814_/A1 vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2389_ _2389_/A _2389_/B vssd1 vssd1 vccd1 vccd1 _2861_/B sky130_fd_sc_hd__nand2_1
X_4128_ _4229_/A _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__and3_1
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4059_ _4059_/A _4059_/B _4059_/C vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__or3_1
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3430_ _4453_/Q _3565_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4453_/D sky130_fd_sc_hd__mux2_1
X_3361_ _4416_/Q _4335_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4416_/D sky130_fd_sc_hd__mux2_1
X_2312_ _4631_/Q _3608_/A vssd1 vssd1 vccd1 vccd1 _3601_/B sky130_fd_sc_hd__or2_1
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3288_/B _3288_/C _2385_/B vssd1 vssd1 vccd1 vccd1 _3292_/X sky130_fd_sc_hd__o21a_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2243_/A _4238_/A vssd1 vssd1 vccd1 vccd1 _2243_/Y sky130_fd_sc_hd__nor2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4677_ _4678_/CLK _4677_/D vssd1 vssd1 vccd1 vccd1 _4677_/Q sky130_fd_sc_hd__dfxtp_1
X_3628_ _3628_/A _3628_/B vssd1 vssd1 vccd1 vccd1 _3851_/C sky130_fd_sc_hd__nor2_1
Xoutput28 _4708_/X vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_4
Xoutput17 _4607_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_4
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3559_ _4568_/Q _3577_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4568_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _4413_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__and3_1
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4600_ _4626_/CLK _4600_/D vssd1 vssd1 vccd1 vccd1 _4600_/Q sky130_fd_sc_hd__dfxtp_1
X_2861_ _2861_/A _2861_/B _2861_/C vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__or3_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2792_ _2353_/X _2789_/X _2791_/X vssd1 vssd1 vccd1 vccd1 _2793_/B sky130_fd_sc_hd__a21bo_1
X_4531_ _4683_/CLK _4531_/D vssd1 vssd1 vccd1 vccd1 _4531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4462_ _4481_/CLK _4462_/D vssd1 vssd1 vccd1 vccd1 _4462_/Q sky130_fd_sc_hd__dfxtp_1
X_3413_ _4666_/Q _3412_/X _3417_/S vssd1 vssd1 vccd1 vccd1 _4346_/B sky130_fd_sc_hd__mux2_1
X_4393_ _4698_/CLK _4393_/D vssd1 vssd1 vccd1 vccd1 _4393_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _4401_/Q _4336_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4401_/D sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3276_/C _3274_/Y _3275_/S vssd1 vssd1 vccd1 vccd1 _3275_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2226_ _2373_/C _3993_/B vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__nand2_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3060_ _4415_/Q _4687_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3060_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _4127_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _3962_/Y sky130_fd_sc_hd__nor2_8
X_3893_ _4074_/A _4074_/B vssd1 vssd1 vccd1 vccd1 _3894_/C sky130_fd_sc_hd__or2_2
X_2913_ _3183_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2913_/Y sky130_fd_sc_hd__nand2_1
X_2844_ _2844_/A _2844_/B vssd1 vssd1 vccd1 vccd1 _2844_/Y sky130_fd_sc_hd__nor2_1
X_4514_ _4579_/CLK _4514_/D vssd1 vssd1 vccd1 vccd1 _4514_/Q sky130_fd_sc_hd__dfxtp_1
X_2775_ _4474_/Q _4466_/Q _4458_/Q _4450_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2775_/X sky130_fd_sc_hd__mux4_1
X_4445_ _4552_/CLK _4445_/D vssd1 vssd1 vccd1 vccd1 _4445_/Q sky130_fd_sc_hd__dfxtp_1
X_4376_ _4570_/CLK _4376_/D vssd1 vssd1 vccd1 vccd1 _4376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _4387_/Q _3580_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4387_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3286_/B vssd1 vssd1 vccd1 vccd1 _3258_/Y sky130_fd_sc_hd__inv_2
X_2209_ _3623_/B _4619_/Q vssd1 vssd1 vccd1 vccd1 _2293_/A sky130_fd_sc_hd__nand2_8
X_3189_ _3160_/X _3184_/X _3186_/X _3188_/Y vssd1 vssd1 vccd1 vccd1 _3189_/X sky130_fd_sc_hd__o31a_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_8_clk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _2612_/S _2555_/X _2559_/Y _2904_/A vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__a211o_1
X_2491_ _2938_/A1 _2486_/X _2490_/X _2477_/X _2482_/X vssd1 vssd1 vccd1 vccd1 _2617_/B
+ sky130_fd_sc_hd__o32ai_4
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4213_/B _4212_/B _3947_/X _4229_/Y vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4161_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4092_ _4092_/A _4092_/B vssd1 vssd1 vccd1 vccd1 _4092_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _4368_/Q _4697_/Q _4688_/Q _4416_/Q _3163_/S _3165_/S1 vssd1 vssd1 vccd1 vccd1
+ _3112_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3043_ _3231_/S _3049_/B _3042_/Y _3176_/A _3041_/Y vssd1 vssd1 vccd1 vccd1 _3044_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3945_ _3938_/Y _4114_/B _3872_/Y vssd1 vssd1 vccd1 vccd1 _4177_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3876_ _3964_/B _4132_/A vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__and2_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2827_ _2953_/A _2826_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2758_ _4482_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__and3_1
X_4428_ _4576_/CLK _4428_/D vssd1 vssd1 vccd1 vccd1 _4428_/Q sky130_fd_sc_hd__dfxtp_1
X_2689_ _4352_/Q _3568_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4352_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4679_/CLK _4359_/D vssd1 vssd1 vccd1 vccd1 _4359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout63 _2629_/X vssd1 vssd1 vccd1 vccd1 _3540_/A1 sky130_fd_sc_hd__buf_2
Xfanout41 _3240_/Y vssd1 vssd1 vccd1 vccd1 _4337_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout52 _2919_/Y vssd1 vssd1 vccd1 vccd1 _4320_/A1 sky130_fd_sc_hd__buf_4
Xfanout74 _3775_/B1 vssd1 vssd1 vccd1 vccd1 _3741_/S sky130_fd_sc_hd__buf_4
Xfanout85 _3257_/A1 vssd1 vssd1 vccd1 vccd1 _2938_/A1 sky130_fd_sc_hd__buf_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout96 _2694_/S vssd1 vssd1 vccd1 vccd1 _2636_/S sky130_fd_sc_hd__buf_6
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3666_/B1 _3729_/X _3072_/B _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _4593_/Q _3775_/B1 _3660_/Y vssd1 vssd1 vccd1 vccd1 _4593_/D sky130_fd_sc_hd__a21o_1
X_2612_ _2608_/X _2611_/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3592_ _4624_/Q _4600_/Q vssd1 vssd1 vccd1 vccd1 _3592_/Y sky130_fd_sc_hd__xnor2_1
X_2543_ _2953_/A _2543_/B vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__nand2_2
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2474_ _4533_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__and3_1
X_4213_ _4213_/A _4213_/B _3905_/A vssd1 vssd1 vccd1 vccd1 _4215_/B sky130_fd_sc_hd__or3b_1
XFILLER_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4144_ _4141_/Y _4142_/X _4143_/X vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__o21ba_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _4229_/A _4103_/C _4073_/Y _4095_/B vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__a31o_1
X_3026_ _3239_/A _2975_/Y _3022_/X _3025_/X vssd1 vssd1 vccd1 vccd1 _3026_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ _3896_/A _3926_/X _4260_/B _4264_/A vssd1 vssd1 vccd1 vccd1 _3928_/Y sky130_fd_sc_hd__o211ai_1
X_3859_ _3860_/A _3933_/B vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout231 _2373_/C vssd1 vssd1 vccd1 vccd1 _2366_/B sky130_fd_sc_hd__buf_8
Xfanout220 _2292_/B vssd1 vssd1 vccd1 vccd1 _3623_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout264 _3163_/S vssd1 vssd1 vccd1 vccd1 _3108_/S sky130_fd_sc_hd__buf_6
Xfanout253 _3265_/A vssd1 vssd1 vccd1 vccd1 _3266_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout242 _2889_/A vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__buf_6
Xfanout275 _4436_/Q vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__buf_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2190_ _3623_/B vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4693_ _4694_/CLK _4693_/D vssd1 vssd1 vccd1 vccd1 _4693_/Q sky130_fd_sc_hd__dfxtp_1
X_3713_ _3713_/A _3713_/B vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__nor2_1
X_3644_ _3689_/A _2617_/B _3643_/Y vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__o21ai_1
X_3575_ _4582_/Q _4313_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4582_/D sky130_fd_sc_hd__mux2_1
X_2526_ _4422_/Q _4430_/Q _2809_/S vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__mux2_1
X_2457_ _4492_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__and3_1
X_2388_ _4664_/Q _2847_/A1 _2768_/B1 _2373_/B _2382_/X vssd1 vssd1 vccd1 vccd1 _2388_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4127_ _4127_/A _4127_/B _4127_/C vssd1 vssd1 vccd1 vccd1 _4128_/C sky130_fd_sc_hd__or3_1
XFILLER_83_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4058_ _4073_/B _4221_/A _3941_/X _3931_/A vssd1 vssd1 vccd1 vccd1 _4059_/C sky130_fd_sc_hd__o211a_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ _3007_/X _3008_/X _3261_/A vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3360_ _4415_/Q _4334_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4415_/D sky130_fd_sc_hd__mux2_1
X_2311_ _3581_/B _4437_/Q _4439_/Q _2289_/X _2308_/Y vssd1 vssd1 vccd1 vccd1 _2316_/B
+ sky130_fd_sc_hd__o32a_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _2364_/Y _3259_/Y _3289_/X _3282_/Y vssd1 vssd1 vccd1 vccd1 _3291_/X sky130_fd_sc_hd__o31a_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2293_/A _3387_/B vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__or2_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4694_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4676_ _4694_/CLK _4676_/D vssd1 vssd1 vccd1 vccd1 _4676_/Q sky130_fd_sc_hd__dfxtp_1
X_3627_ _3627_/A _3627_/B _2341_/B vssd1 vssd1 vccd1 vccd1 _3628_/B sky130_fd_sc_hd__or3b_1
Xoutput29 _4636_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_4
X_3558_ _4567_/Q _4314_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4567_/D sky130_fd_sc_hd__mux2_1
Xoutput18 _4608_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_4
X_2509_ _2507_/Y _2508_/X _4071_/A2 _2348_/B vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ _4506_/Q _4317_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4506_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4587_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4613_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2860_ _3826_/A _3278_/A _2860_/C _2860_/D vssd1 vssd1 vccd1 vccd1 _2861_/C sky130_fd_sc_hd__or4_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2791_ _2652_/A _2766_/Y _2790_/X _2655_/Y _2571_/A vssd1 vssd1 vccd1 vccd1 _2791_/X
+ sky130_fd_sc_hd__o221a_1
X_4530_ _4570_/CLK _4530_/D vssd1 vssd1 vccd1 vccd1 _4530_/Q sky130_fd_sc_hd__dfxtp_1
X_4461_ _4464_/CLK _4461_/D vssd1 vssd1 vccd1 vccd1 _4461_/Q sky130_fd_sc_hd__dfxtp_1
X_3412_ _3938_/B _4081_/A _3411_/Y vssd1 vssd1 vccd1 vccd1 _3412_/X sky130_fd_sc_hd__o21a_1
X_4392_ _4683_/CLK _4392_/D vssd1 vssd1 vccd1 vccd1 _4392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3343_ _4400_/Q _3577_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4400_/D sky130_fd_sc_hd__mux2_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3276_/C _3274_/B vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__xnor2_2
X_2225_ _3993_/A _2261_/B vssd1 vssd1 vccd1 vccd1 _2225_/Y sky130_fd_sc_hd__nor2_4
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _4390_/Q _4382_/Q _3089_/S vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__mux2_1
X_4659_ _4671_/CLK _4659_/D vssd1 vssd1 vccd1 vccd1 _4659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _3961_/Y sky130_fd_sc_hd__inv_2
X_2912_ _3280_/B1 _2910_/Y _2911_/Y _2909_/X vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__o31a_1
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3892_ _3941_/A _4063_/A vssd1 vssd1 vccd1 vccd1 _4074_/B sky130_fd_sc_hd__and2b_1
X_2843_ _3041_/A _2840_/X _2842_/X _2844_/A vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__o211a_1
X_2774_ _2953_/A _2769_/X _2773_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__a211o_4
X_4513_ _4545_/CLK _4513_/D vssd1 vssd1 vccd1 vccd1 _4513_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_7_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4543_/CLK sky130_fd_sc_hd__clkbuf_16
X_4444_ _4548_/CLK _4444_/D vssd1 vssd1 vccd1 vccd1 _4444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4375_ _4679_/CLK _4375_/D vssd1 vssd1 vccd1 vccd1 _4375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _4386_/Q _4317_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4386_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3257_/A1 _3256_/X _3249_/X vssd1 vssd1 vccd1 vccd1 _3286_/B sky130_fd_sc_hd__o21a_4
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2208_ _2292_/B _2360_/B vssd1 vssd1 vccd1 vccd1 _2473_/A sky130_fd_sc_hd__or2_4
X_3188_ _4689_/Q _3237_/C _3187_/Y vssd1 vssd1 vccd1 vccd1 _3188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2490_ _2644_/S _2487_/X _2489_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__o211a_1
X_4160_ _3872_/Y _4132_/Y _3910_/B vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3111_ _3261_/A _3110_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__a21o_1
X_4091_ _4091_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__or2_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3042_ _3231_/S _3739_/A vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3944_ _4116_/A _4113_/B vssd1 vssd1 vccd1 vccd1 _4114_/B sky130_fd_sc_hd__nand2_1
X_3875_ _3938_/B _3938_/A vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__nand2b_4
X_2826_ _4579_/Q _4523_/Q _4515_/Q _4355_/Q _2824_/S _2404_/A vssd1 vssd1 vccd1 vccd1
+ _2826_/X sky130_fd_sc_hd__mux4_1
X_2757_ _4498_/Q _4554_/Q _2811_/S vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__mux2_1
X_2688_ _2571_/A _2686_/X _2687_/Y _2685_/X vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__o31a_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4427_ _4573_/CLK _4427_/D vssd1 vssd1 vccd1 vccd1 _4427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4358_ _4582_/CLK _4358_/D vssd1 vssd1 vccd1 vccd1 _4358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4289_ _4288_/X _3938_/B _4309_/S vssd1 vssd1 vccd1 vccd1 _4670_/D sky130_fd_sc_hd__mux2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _4310_/A _4310_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3317_/S sky130_fd_sc_hd__and3_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout42 _3189_/X vssd1 vssd1 vccd1 vccd1 _4316_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout53 _2919_/Y vssd1 vssd1 vccd1 vccd1 _4331_/A1 sky130_fd_sc_hd__buf_2
Xfanout64 _3539_/A1 vssd1 vssd1 vccd1 vccd1 _3566_/A1 sky130_fd_sc_hd__buf_4
Xfanout86 _2454_/X vssd1 vssd1 vccd1 vccd1 _3257_/A1 sky130_fd_sc_hd__buf_12
Xfanout75 _4329_/S vssd1 vssd1 vccd1 vccd1 _3775_/B1 sky130_fd_sc_hd__buf_2
Xfanout97 _2800_/S vssd1 vssd1 vccd1 vccd1 _2694_/S sky130_fd_sc_hd__buf_6
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _3739_/B _3658_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__a21oi_2
X_2611_ _2669_/C _2610_/Y _2841_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
X_3591_ _4627_/Q _4603_/Q vssd1 vssd1 vccd1 vccd1 _3591_/Y sky130_fd_sc_hd__xnor2_1
X_2542_ _4574_/Q _4518_/Q _4510_/Q _4350_/Q _2824_/S _2825_/B2 vssd1 vssd1 vccd1 vccd1
+ _2543_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4212_ _4213_/B _4212_/B _4212_/C vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand3_1
X_2473_ _2473_/A _2473_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__or3_4
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4143_ _3935_/A _4267_/A2 _4267_/B1 _4658_/Q _4228_/B vssd1 vssd1 vccd1 vccd1 _4143_/X
+ sky130_fd_sc_hd__a221o_1
X_4074_ _4074_/A _4074_/B vssd1 vssd1 vccd1 vccd1 _4074_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3160_/B1 _2999_/X _3000_/X _3024_/X _2382_/X vssd1 vssd1 vccd1 vccd1 _3025_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3927_ _3927_/A _3927_/B vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__nor2_4
X_3858_ _3860_/A _3933_/B vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__and2_2
X_3789_ _3619_/B _3787_/X _3788_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4610_/D sky130_fd_sc_hd__o211a_1
X_2809_ _4467_/Q _4475_/Q _2809_/S vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout232 _4056_/B vssd1 vssd1 vccd1 vccd1 _2373_/C sky130_fd_sc_hd__buf_8
Xfanout221 _4622_/Q vssd1 vssd1 vccd1 vccd1 _2292_/B sky130_fd_sc_hd__buf_6
Xfanout210 _3259_/A vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout243 _4442_/Q vssd1 vssd1 vccd1 vccd1 _2889_/A sky130_fd_sc_hd__buf_12
Xfanout265 _4440_/Q vssd1 vssd1 vccd1 vccd1 _3163_/S sky130_fd_sc_hd__buf_4
Xfanout254 _3165_/S1 vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__buf_4
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout276 _4347_/A vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4692_ _4692_/CLK _4692_/D vssd1 vssd1 vccd1 vccd1 _4692_/Q sky130_fd_sc_hd__dfxtp_2
X_3712_ _2996_/A _3631_/X _3989_/B _3711_/X vssd1 vssd1 vccd1 vccd1 _3713_/B sky130_fd_sc_hd__o22a_1
X_3643_ _3689_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _3643_/Y sky130_fd_sc_hd__nand2_1
X_3574_ _4581_/Q _4312_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4581_/D sky130_fd_sc_hd__mux2_1
X_2525_ _4510_/Q _2636_/S _2524_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__a211o_1
X_2456_ _4476_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__and3_1
XFILLER_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _3938_/A _4125_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4658_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2387_ _4665_/Q _2847_/A1 _2383_/X vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__a21o_4
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4057_/A _4057_/B vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__or2_4
X_3008_ _4382_/Q _4390_/Q _4406_/Q _4398_/Q _3108_/S _3113_/S1 vssd1 vssd1 vccd1 vccd1
+ _3008_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2310_ _3623_/B _2360_/B _2292_/B _4619_/Q vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__or4bb_4
X_3290_ _3290_/A _3290_/B vssd1 vssd1 vccd1 vccd1 _3290_/X sky130_fd_sc_hd__and2_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2241_ _2293_/A _3387_/B vssd1 vssd1 vccd1 vccd1 _2241_/Y sky130_fd_sc_hd__nor2_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4675_ _4691_/CLK _4675_/D vssd1 vssd1 vccd1 vccd1 _4675_/Q sky130_fd_sc_hd__dfxtp_4
X_3626_ _3987_/B _3990_/B _3625_/X vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__o21ai_1
X_3557_ _4566_/Q _4313_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4566_/D sky130_fd_sc_hd__mux2_1
Xoutput19 _4609_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_4
X_2508_ _3275_/S _2513_/B _2348_/B vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__a21o_1
X_3488_ _4505_/Q _4316_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4505_/D sky130_fd_sc_hd__mux2_1
X_2439_ _2440_/B _2440_/C _4615_/Q vssd1 vssd1 vccd1 vccd1 _2439_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4109_ _4059_/A _4108_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4109_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2790_ _2790_/A _2848_/B vssd1 vssd1 vccd1 vccd1 _2790_/X sky130_fd_sc_hd__xor2_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4548_/CLK _4460_/D vssd1 vssd1 vccd1 vccd1 _4460_/Q sky130_fd_sc_hd__dfxtp_1
X_3411_ _3993_/A _4081_/A _3405_/A vssd1 vssd1 vccd1 vccd1 _3411_/Y sky130_fd_sc_hd__a21oi_1
X_4391_ _4679_/CLK _4391_/D vssd1 vssd1 vccd1 vccd1 _4391_/Q sky130_fd_sc_hd__dfxtp_1
X_3342_ _4399_/Q _4334_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4399_/D sky130_fd_sc_hd__mux2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3273_/A _3273_/B _3273_/C _3761_/B vssd1 vssd1 vccd1 vccd1 _3274_/B sky130_fd_sc_hd__or4_2
X_2224_ _3846_/A _2373_/B vssd1 vssd1 vccd1 vccd1 _2261_/B sky130_fd_sc_hd__or2_4
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2988_ _3086_/A _2985_/X _2987_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__o211a_1
X_4658_ _4671_/CLK _4658_/D vssd1 vssd1 vccd1 vccd1 _4658_/Q sky130_fd_sc_hd__dfxtp_4
X_3609_ _2217_/Y _3987_/B _3990_/B _3604_/Y _3605_/X vssd1 vssd1 vccd1 vccd1 _3613_/C
+ sky130_fd_sc_hd__o311a_1
X_4589_ _4692_/CLK _4589_/D vssd1 vssd1 vccd1 vccd1 _4589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _4177_/A _3960_/B vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__or2_4
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2911_ _3742_/A _3013_/B vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__nor2_1
X_3891_ _3896_/A _4244_/A _3980_/A vssd1 vssd1 vccd1 vccd1 _3891_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2842_ _2837_/Y _2838_/X _2841_/X _2612_/S _2904_/A vssd1 vssd1 vccd1 vccd1 _2842_/X
+ sky130_fd_sc_hd__a221o_1
X_2773_ _2770_/X _2771_/X _2772_/X _2893_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2773_/X
+ sky130_fd_sc_hd__o221a_1
X_4512_ _4537_/CLK _4512_/D vssd1 vssd1 vccd1 vccd1 _4512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4443_ _4549_/CLK _4443_/D vssd1 vssd1 vccd1 vccd1 _4443_/Q sky130_fd_sc_hd__dfxtp_1
X_4374_ _4678_/CLK _4374_/D vssd1 vssd1 vccd1 vccd1 _4374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _4385_/Q _4316_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4385_/D sky130_fd_sc_hd__mux2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3252_/X _3255_/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2207_ _3623_/C _2360_/B vssd1 vssd1 vccd1 vccd1 _4046_/A sky130_fd_sc_hd__nor2_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3187_ _4689_/Q _3237_/C _2389_/A vssd1 vssd1 vccd1 vccd1 _3187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3110_ _4528_/Q _4568_/Q _4560_/Q _4504_/Q _3108_/S _3113_/S1 vssd1 vssd1 vccd1 vccd1
+ _3110_/X sky130_fd_sc_hd__mux4_1
X_4090_ _4091_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4264_/B sky130_fd_sc_hd__nor2_2
XFILLER_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3041_ _3041_/A _3273_/A _3739_/A vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3943_ _4074_/A _4092_/B _4103_/B vssd1 vssd1 vccd1 vccd1 _4113_/B sky130_fd_sc_hd__a21bo_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3964_/B sky130_fd_sc_hd__nand2b_4
X_2825_ _2822_/X _2823_/X _2824_/X _2825_/B2 _2549_/A vssd1 vssd1 vccd1 vccd1 _2825_/X
+ sky130_fd_sc_hd__o221a_1
X_2756_ _2645_/S _2753_/X _2755_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__a31o_2
X_2687_ _4488_/Q _2745_/C vssd1 vssd1 vccd1 vccd1 _2687_/Y sky130_fd_sc_hd__nor2_1
X_4426_ _4572_/CLK _4426_/D vssd1 vssd1 vccd1 vccd1 _4426_/Q sky130_fd_sc_hd__dfxtp_1
X_4357_ _4581_/CLK _4357_/D vssd1 vssd1 vccd1 vccd1 _4357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4288_ input6/X _4287_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__mux2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _4371_/Q _4338_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4371_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3239_ _3239_/A _3239_/B _3239_/C vssd1 vssd1 vccd1 vccd1 _3239_/X sky130_fd_sc_hd__and3_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout65 _2572_/X vssd1 vssd1 vccd1 vccd1 _3539_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout54 _2856_/Y vssd1 vssd1 vccd1 vccd1 _3571_/A1 sky130_fd_sc_hd__buf_4
Xfanout43 _3189_/X vssd1 vssd1 vccd1 vccd1 _4336_/A1 sky130_fd_sc_hd__buf_2
Xfanout76 _3630_/X vssd1 vssd1 vccd1 vccd1 _4329_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout98 _2932_/S vssd1 vssd1 vccd1 vccd1 _2934_/S sky130_fd_sc_hd__buf_6
Xfanout87 _2453_/X vssd1 vssd1 vccd1 vccd1 _2984_/B1 sky130_fd_sc_hd__buf_8
XFILLER_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ _4629_/Q _4605_/Q vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__xnor2_1
X_2610_ _2670_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2610_/Y sky130_fd_sc_hd__nor2_1
X_2541_ _2541_/A _2617_/C vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__xnor2_1
X_2472_ _2473_/A _2473_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__nor3_4
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _3934_/A _4210_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4661_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4142_ _3964_/A _4132_/A _4115_/X _4117_/B vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4073_ _4092_/A _4073_/B vssd1 vssd1 vccd1 vccd1 _4073_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3024_ _3183_/A _3020_/X _3023_/X _3282_/A vssd1 vssd1 vccd1 vccd1 _3024_/X sky130_fd_sc_hd__o211a_1
X_3926_ _3904_/Y _3925_/Y _4264_/A _3903_/X vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__o211a_1
X_3857_ _3855_/B _3857_/B vssd1 vssd1 vccd1 vccd1 _3896_/B sky130_fd_sc_hd__nand2b_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2808_ _4459_/Q _2809_/S _2807_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__a211o_1
X_3788_ _4610_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__or2_1
X_2739_ _4673_/Q _2345_/Y _2846_/S _2738_/X vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__o211a_1
Xfanout222 _4621_/Q vssd1 vssd1 vccd1 vccd1 _2360_/B sky130_fd_sc_hd__buf_6
Xfanout211 _4663_/Q vssd1 vssd1 vccd1 vccd1 _3259_/A sky130_fd_sc_hd__clkbuf_4
Xfanout200 _2194_/Y vssd1 vssd1 vccd1 vccd1 _3760_/A sky130_fd_sc_hd__clkbuf_16
X_4409_ _4681_/CLK _4409_/D vssd1 vssd1 vccd1 vccd1 _4409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout233 _4057_/B vssd1 vssd1 vccd1 vccd1 _4056_/B sky130_fd_sc_hd__buf_6
Xfanout255 _4441_/Q vssd1 vssd1 vccd1 vccd1 _3165_/S1 sky130_fd_sc_hd__buf_4
Xfanout244 _4442_/Q vssd1 vssd1 vccd1 vccd1 _3261_/A sky130_fd_sc_hd__buf_6
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout277 _2195_/Y vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout266 _3264_/S vssd1 vssd1 vccd1 vccd1 _3216_/S sky130_fd_sc_hd__buf_6
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3711_ _3709_/X _3710_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__mux2_1
X_4691_ _4691_/CLK _4691_/D vssd1 vssd1 vccd1 vccd1 _4691_/Q sky130_fd_sc_hd__dfxtp_2
X_3642_ _3640_/Y _3641_/X _4591_/Q _3775_/B1 vssd1 vssd1 vccd1 vccd1 _4591_/D sky130_fd_sc_hd__a2bb2o_1
X_3573_ _4580_/Q _4320_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4580_/D sky130_fd_sc_hd__mux2_1
X_2524_ _4350_/Q _2798_/B _2798_/C vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__and3_1
X_2455_ _2937_/C1 _2450_/X _2452_/X _2938_/A1 vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__o31ai_4
X_2386_ _4665_/Q _2847_/A1 _2383_/X vssd1 vssd1 vccd1 vccd1 _2858_/A sky130_fd_sc_hd__a21oi_4
X_4125_ _4240_/A _4111_/Y _4124_/X _4270_/B input6/X vssd1 vssd1 vccd1 vccd1 _4125_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4056_ _4057_/A _4056_/B vssd1 vssd1 vccd1 vccd1 _4221_/A sky130_fd_sc_hd__nor2_4
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3007_ _4366_/Q _4695_/Q _4686_/Q _4414_/Q _3108_/S _3113_/S1 vssd1 vssd1 vccd1 vccd1
+ _3007_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3909_ _4177_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _4204_/B sky130_fd_sc_hd__nand2_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2240_ _2360_/A _3622_/B vssd1 vssd1 vccd1 vccd1 _3387_/B sky130_fd_sc_hd__nand2_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4674_ _4674_/CLK _4674_/D vssd1 vssd1 vccd1 vccd1 _4674_/Q sky130_fd_sc_hd__dfxtp_4
X_3625_ _3581_/D _2351_/C _3399_/X _2233_/Y _3608_/B vssd1 vssd1 vccd1 vccd1 _3625_/X
+ sky130_fd_sc_hd__o221a_1
X_3556_ _4565_/Q _4332_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4565_/D sky130_fd_sc_hd__mux2_1
X_2507_ _3275_/S _3643_/B vssd1 vssd1 vccd1 vccd1 _2507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3487_ _4504_/Q _3577_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4504_/D sky130_fd_sc_hd__mux2_1
X_2438_ _4057_/A _2454_/S _2436_/X vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2369_ _2372_/C _4013_/S vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__nor2_2
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _3938_/A _3938_/B _4057_/X _4107_/X vssd1 vssd1 vccd1 vccd1 _4108_/X sky130_fd_sc_hd__o31a_1
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4039_ _4062_/B _2373_/Y _4038_/Y _3987_/A _2373_/C vssd1 vssd1 vccd1 vccd1 _4040_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3410_ _4665_/Q _3417_/S _3409_/Y vssd1 vssd1 vccd1 vccd1 _4441_/D sky130_fd_sc_hd__o21a_1
X_4390_ _4582_/CLK _4390_/D vssd1 vssd1 vccd1 vccd1 _4390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3341_ _4398_/Q _4313_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4398_/D sky130_fd_sc_hd__mux2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3276_/C vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__inv_2
X_2223_ _4057_/A _2373_/B vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__nor2_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2987_ _4686_/Q _3089_/S _2986_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _2987_/X sky130_fd_sc_hd__a211o_1
X_4657_ _4671_/CLK _4657_/D vssd1 vssd1 vccd1 vccd1 _4657_/Q sky130_fd_sc_hd__dfxtp_4
X_3608_ _3608_/A _3608_/B vssd1 vssd1 vccd1 vccd1 _3608_/Y sky130_fd_sc_hd__nor2_1
X_4588_ _4692_/CLK _4588_/D vssd1 vssd1 vccd1 vccd1 _4588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3539_ _4550_/Q _3539_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4550_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2910_ _3760_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2910_/Y sky130_fd_sc_hd__nor2_1
X_3890_ _3951_/A _4216_/A _3903_/A vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__a21oi_2
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2841_ _3699_/B _2840_/X _2841_/S vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2772_ _4434_/Q _4426_/Q _2892_/S vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__mux2_1
X_4511_ _4543_/CLK _4511_/D vssd1 vssd1 vccd1 vccd1 _4511_/Q sky130_fd_sc_hd__dfxtp_1
X_4442_ _4549_/CLK _4442_/D vssd1 vssd1 vccd1 vccd1 _4442_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4373_ _4678_/CLK _4373_/D vssd1 vssd1 vccd1 vccd1 _4373_/Q sky130_fd_sc_hd__dfxtp_1
X_3324_ _4384_/Q _3577_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4384_/D sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3253_/X _3254_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__mux2_1
X_2206_ _2274_/A _4439_/Q _3989_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__and3_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3186_ _3185_/A _3158_/X _3185_/Y _2382_/X vssd1 vssd1 vccd1 vccd1 _3186_/X sky130_fd_sc_hd__o211a_1
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3040_ _3040_/A _3040_/B vssd1 vssd1 vccd1 vccd1 _3049_/B sky130_fd_sc_hd__or2_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3942_ _4643_/Q _3941_/X _4073_/B vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__a21bo_1
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3873_ _3960_/B _3910_/B vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__or2_4
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2824_ _4435_/Q _4427_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2755_ _4578_/Q _2934_/S _2754_/X _2937_/A1 vssd1 vssd1 vccd1 vccd1 _2755_/X sky130_fd_sc_hd__a211o_1
X_2686_ _4488_/Q _2745_/C vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__and2_1
X_4425_ _4537_/CLK _4425_/D vssd1 vssd1 vccd1 vccd1 _4425_/Q sky130_fd_sc_hd__dfxtp_1
X_4356_ _4580_/CLK _4356_/D vssd1 vssd1 vccd1 vccd1 _4356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _4370_/Q _4337_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4370_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4287_ _3938_/A _4278_/Y _4286_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__a22o_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _4689_/Q _3237_/C _4690_/Q vssd1 vssd1 vccd1 vccd1 _3239_/C sky130_fd_sc_hd__o21ai_1
X_3169_ _3167_/X _3168_/X _4442_/Q vssd1 vssd1 vccd1 vccd1 _3169_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout44 _4335_/A1 vssd1 vssd1 vccd1 vccd1 _3577_/A1 sky130_fd_sc_hd__buf_4
Xfanout55 _2856_/Y vssd1 vssd1 vccd1 vccd1 _3544_/A1 sky130_fd_sc_hd__buf_2
Xfanout66 _2520_/X vssd1 vssd1 vccd1 vccd1 _3565_/A1 sky130_fd_sc_hd__buf_4
Xfanout77 _3630_/X vssd1 vssd1 vccd1 vccd1 _3749_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout99 _2800_/S vssd1 vssd1 vccd1 vccd1 _2932_/S sky130_fd_sc_hd__buf_6
Xfanout88 _2453_/X vssd1 vssd1 vccd1 vccd1 _3249_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2540_ _2540_/A _2617_/C vssd1 vssd1 vccd1 vccd1 _2566_/B sky130_fd_sc_hd__xnor2_1
X_2471_ _3623_/C _2473_/B vssd1 vssd1 vccd1 vccd1 _3391_/B sky130_fd_sc_hd__or2_4
X_4210_ _4240_/A _4197_/Y _4209_/X _4270_/B input9/X vssd1 vssd1 vccd1 vccd1 _4210_/X
+ sky130_fd_sc_hd__a32o_1
X_4141_ _4132_/A _4115_/X _3964_/A vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _4072_/A _4074_/A vssd1 vssd1 vccd1 vccd1 _4072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3023_ _3230_/A _3023_/B vssd1 vssd1 vccd1 vccd1 _3023_/X sky130_fd_sc_hd__or2_1
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3925_ _3908_/A _3924_/X _3904_/Y _3905_/X vssd1 vssd1 vccd1 vccd1 _3925_/Y sky130_fd_sc_hd__a211oi_4
X_3856_ _3855_/B _3857_/B vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__and2b_2
X_3787_ _4602_/Q _4594_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__mux2_1
X_2807_ _4451_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__and3_1
X_2738_ _2735_/X _2736_/X _2737_/X vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__a21o_1
X_4408_ _4584_/CLK _4408_/D vssd1 vssd1 vccd1 vccd1 _4408_/Q sky130_fd_sc_hd__dfxtp_1
X_2669_ _3643_/B _3652_/B _2669_/C _3670_/B vssd1 vssd1 vccd1 vccd1 _2834_/A sky130_fd_sc_hd__and4_4
Xfanout223 _4621_/Q vssd1 vssd1 vccd1 vccd1 _3622_/B sky130_fd_sc_hd__buf_2
Xfanout212 _4661_/Q vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__buf_6
Xfanout201 _2194_/Y vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__buf_12
Xfanout234 _4617_/Q vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__buf_4
X_4339_ _4632_/Q _3602_/B _4300_/S _3383_/B vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__o211a_1
Xfanout245 _2954_/S1 vssd1 vssd1 vccd1 vccd1 _2404_/A sky130_fd_sc_hd__clkbuf_8
Xfanout256 _2824_/S vssd1 vssd1 vccd1 vccd1 _2661_/S sky130_fd_sc_hd__buf_6
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout278 _2274_/A vssd1 vssd1 vccd1 vccd1 _3828_/A sky130_fd_sc_hd__buf_4
Xfanout267 _4440_/Q vssd1 vssd1 vccd1 vccd1 _3264_/S sky130_fd_sc_hd__buf_8
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3710_ _4684_/Q _3691_/C _3708_/X _2331_/A vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__o22a_1
X_4690_ _4696_/CLK _4690_/D vssd1 vssd1 vccd1 vccd1 _4690_/Q sky130_fd_sc_hd__dfxtp_2
X_3641_ _3731_/A1 _4061_/B _3640_/A _2413_/X _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3641_/X
+ sky130_fd_sc_hd__a221o_1
X_3572_ _3572_/A _4310_/A _4330_/A vssd1 vssd1 vccd1 vccd1 _3580_/S sky130_fd_sc_hd__and3_4
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2523_ _4574_/Q _2800_/S _2522_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__a211o_1
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2454_ _4647_/Q _3689_/A _2454_/S vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__mux2_2
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2385_ _2385_/A _2385_/B vssd1 vssd1 vccd1 vccd1 _2385_/Y sky130_fd_sc_hd__nor2_8
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4124_ _3974_/Y _4228_/B _4112_/X _4123_/X vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__a31o_1
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4055_ _3941_/A _4063_/A _3584_/Y _4267_/A2 _3917_/A vssd1 vssd1 vccd1 vccd1 _4059_/B
+ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_48_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3006_ _3261_/A _3005_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _3006_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ _3908_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__nand2_1
X_3839_ _3802_/A _3618_/A _4708_/A vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/CLK _4673_/D vssd1 vssd1 vccd1 vccd1 _4673_/Q sky130_fd_sc_hd__dfxtp_4
X_3624_ _3836_/A _3989_/A _3624_/C _3624_/D vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__or4_1
X_3555_ _4564_/Q _4320_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4564_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3486_ _4503_/Q _4314_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4503_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2506_ _2500_/X _2502_/X _2505_/X _2668_/A1 vssd1 vssd1 vccd1 vccd1 _2513_/B sky130_fd_sc_hd__o22a_4
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2437_ _4057_/A _2454_/S _2436_/X vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__a21o_1
X_2368_ _2368_/A _2368_/B vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__or2_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4107_ _4107_/A _4123_/B _4102_/X _4106_/X vssd1 vssd1 vccd1 vccd1 _4107_/X sky130_fd_sc_hd__or4bb_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2299_ _3629_/B _2300_/C vssd1 vssd1 vccd1 vccd1 _2425_/A sky130_fd_sc_hd__or2_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4038_ _3629_/A _2432_/B _2300_/A vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ _4397_/Q _4332_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4397_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3270_/A _3261_/Y _3266_/X _3270_/Y vssd1 vssd1 vccd1 vccd1 _3276_/C sky130_fd_sc_hd__a31o_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2302_/A _4003_/A vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__or2_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2986_ _4414_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__and3_1
X_4656_ _4667_/CLK _4656_/D vssd1 vssd1 vccd1 vccd1 _4656_/Q sky130_fd_sc_hd__dfxtp_2
X_3607_ _3633_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3608_/B sky130_fd_sc_hd__nand2_1
X_4587_ _4587_/CLK _4587_/D vssd1 vssd1 vccd1 vccd1 _4587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _4549_/Q _3538_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4549_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3469_ _4488_/Q _3568_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4488_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _3013_/A _2840_/B vssd1 vssd1 vccd1 vccd1 _2840_/X sky130_fd_sc_hd__and2_1
X_2771_ _2950_/S _4538_/Q _2893_/A vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__a21bo_1
X_4510_ _4574_/CLK _4510_/D vssd1 vssd1 vccd1 vccd1 _4510_/Q sky130_fd_sc_hd__dfxtp_1
X_4441_ _4551_/CLK _4441_/D vssd1 vssd1 vccd1 vccd1 _4441_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4580_/CLK _4372_/D vssd1 vssd1 vccd1 vccd1 _4372_/Q sky130_fd_sc_hd__dfxtp_1
X_3323_ _4383_/Q _4314_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4383_/D sky130_fd_sc_hd__mux2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _4403_/Q _4411_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__mux2_1
X_2205_ _4590_/Q _3618_/A _4588_/Q vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__or3_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _3185_/A _3212_/A _3185_/C vssd1 vssd1 vccd1 vccd1 _3185_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2969_ _2652_/A _2942_/X _2945_/X _2655_/Y _2968_/Y vssd1 vssd1 vccd1 vccd1 _2969_/X
+ sky130_fd_sc_hd__o221a_1
X_4708_ _4708_/A vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__clkbuf_2
X_4639_ _4643_/CLK _4639_/D vssd1 vssd1 vccd1 vccd1 _4639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _3941_/A _4063_/A vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__or2_1
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _3960_/B _3910_/B vssd1 vssd1 vccd1 vccd1 _3872_/Y sky130_fd_sc_hd__nor2_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2823_ _2823_/A1 _4539_/Q _2404_/A vssd1 vssd1 vccd1 vccd1 _2823_/X sky130_fd_sc_hd__a21bo_1
X_2754_ _4522_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__and3_1
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2685_ _2685_/A _2685_/B vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__or2_1
X_4424_ _4544_/CLK _4424_/D vssd1 vssd1 vccd1 vccd1 _4424_/Q sky130_fd_sc_hd__dfxtp_1
X_4355_ _4545_/CLK _4355_/D vssd1 vssd1 vccd1 vccd1 _4355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _4369_/Q _4336_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4369_/D sky130_fd_sc_hd__mux2_1
X_4286_ _4666_/Q _2367_/Y _3629_/Y _4650_/Q vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__a22o_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _4689_/Q _4690_/Q _3237_/C vssd1 vssd1 vccd1 vccd1 _3239_/B sky130_fd_sc_hd__or3_2
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3168_ _4385_/Q _4393_/Q _4409_/Q _4401_/Q _3264_/S _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3168_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3099_ _3086_/A _3096_/X _3098_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3099_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout45 _3132_/Y vssd1 vssd1 vccd1 vccd1 _4335_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout56 _2796_/Y vssd1 vssd1 vccd1 vccd1 _3570_/A1 sky130_fd_sc_hd__buf_4
Xfanout78 _2708_/B vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__clkbuf_4
Xfanout67 _2520_/X vssd1 vssd1 vccd1 vccd1 _3538_/A1 sky130_fd_sc_hd__buf_2
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout89 _2645_/S vssd1 vssd1 vccd1 vccd1 _2937_/C1 sky130_fd_sc_hd__buf_8
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2470_ _4348_/Q _3564_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4348_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4140_ _4140_/A _4140_/B vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4071_ _3917_/A _4071_/A2 _4221_/A vssd1 vssd1 vccd1 vccd1 _4071_/X sky130_fd_sc_hd__o21a_1
X_3022_ _3290_/A _2994_/Y _3021_/Y _2389_/B vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__a211o_1
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3924_ _4204_/B _4204_/C _4204_/A vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__a21o_2
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3855_ _3857_/B _3855_/B vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__nand2b_4
X_2806_ _2937_/C1 _2803_/X _2805_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__a31o_2
X_3786_ _3619_/B _3784_/X _3785_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4609_/D sky130_fd_sc_hd__o211a_1
X_2737_ _2337_/C _2729_/X _2422_/A vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__a21o_1
X_2668_ _2668_/A1 _2658_/Y _2662_/Y _2664_/Y _2666_/Y vssd1 vssd1 vccd1 vccd1 _3671_/B
+ sky130_fd_sc_hd__a32o_4
X_4407_ _4679_/CLK _4407_/D vssd1 vssd1 vccd1 vccd1 _4407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout213 _4660_/Q vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__buf_6
Xfanout202 _3846_/B vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__buf_12
X_2599_ _2596_/X _2597_/X _2598_/X _2776_/S1 _3036_/S vssd1 vssd1 vccd1 vccd1 _2599_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout235 _4057_/A vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__buf_8
Xfanout224 _4620_/Q vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__buf_8
Xfanout246 _2954_/S1 vssd1 vssd1 vccd1 vccd1 _2825_/B2 sky130_fd_sc_hd__buf_4
X_4338_ _4700_/Q _4338_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4700_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout279 _2195_/Y vssd1 vssd1 vccd1 vccd1 _2274_/A sky130_fd_sc_hd__clkbuf_4
X_4269_ _4269_/A _4269_/B _4269_/C _4262_/X vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__or4b_2
Xfanout268 _4042_/A vssd1 vssd1 vccd1 vccd1 _3581_/B sky130_fd_sc_hd__buf_6
Xfanout257 _2823_/A1 vssd1 vssd1 vccd1 vccd1 _2824_/S sky130_fd_sc_hd__buf_6
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3640_ _3640_/A _3640_/B vssd1 vssd1 vccd1 vccd1 _3640_/Y sky130_fd_sc_hd__nor2_1
X_3571_ _4579_/Q _3571_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4579_/D sky130_fd_sc_hd__mux2_1
X_2522_ _4518_/Q _2863_/B _2863_/C vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__and3_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2453_ _2176_/Y _3760_/A _2454_/S vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__mux2_8
X_2384_ _3832_/B _2384_/B _2384_/C _2384_/D vssd1 vssd1 vccd1 vccd1 _2385_/B sky130_fd_sc_hd__and4_4
X_4123_ _4123_/A _4123_/B _4123_/C _4122_/X vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__or4b_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_4054_ _3610_/Y _4054_/B _4054_/C vssd1 vssd1 vccd1 vccd1 _4272_/S sky130_fd_sc_hd__and3b_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3005_ _4526_/Q _4566_/Q _4558_/Q _4502_/Q _3108_/S _3113_/S1 vssd1 vssd1 vccd1 vccd1
+ _3005_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3907_ _4205_/A _3907_/B vssd1 vssd1 vccd1 vccd1 _3908_/B sky130_fd_sc_hd__or2_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3838_ _4633_/Q _3608_/Y _3837_/Y _2274_/A vssd1 vssd1 vccd1 vccd1 _4633_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3769_ _4605_/Q _3741_/S _3768_/X vssd1 vssd1 vccd1 vccd1 _4605_/D sky130_fd_sc_hd__a21o_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _4672_/CLK _4672_/D vssd1 vssd1 vccd1 vccd1 _4672_/Q sky130_fd_sc_hd__dfxtp_4
X_3623_ _3623_/A _3623_/B _3623_/C _3988_/C vssd1 vssd1 vccd1 vccd1 _3624_/D sky130_fd_sc_hd__and4_1
X_3554_ _3563_/A _4310_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _3562_/S sky130_fd_sc_hd__and3_4
X_2505_ _2503_/X _2504_/X _2889_/A vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__mux2_1
X_3485_ _4502_/Q _4333_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4502_/D sky130_fd_sc_hd__mux2_1
X_2436_ _4645_/Q _2440_/B _2440_/C vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__and3_1
X_2367_ _2368_/A _2368_/B vssd1 vssd1 vccd1 vccd1 _2367_/Y sky130_fd_sc_hd__nor2_8
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4106_ _4262_/A _4127_/C _4103_/X _4105_/X vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2298_ _3987_/A _4062_/B vssd1 vssd1 vccd1 vccd1 _2306_/A sky130_fd_sc_hd__and2_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _4037_/A _4037_/B vssd1 vssd1 vccd1 vccd1 _4655_/D sky130_fd_sc_hd__and2_1
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3270_ _3270_/A _3270_/B vssd1 vssd1 vccd1 vccd1 _3270_/Y sky130_fd_sc_hd__nor2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2302_/A _4003_/A vssd1 vssd1 vccd1 vccd1 _3581_/C sky130_fd_sc_hd__nor2_8
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2985_ _4695_/Q _4366_/Q _3089_/S vssd1 vssd1 vccd1 vccd1 _2985_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4655_ _4673_/CLK _4655_/D vssd1 vssd1 vccd1 vccd1 _4655_/Q sky130_fd_sc_hd__dfxtp_1
X_3606_ _4050_/A _4050_/C vssd1 vssd1 vccd1 vccd1 _3607_/B sky130_fd_sc_hd__nor2_1
X_4586_ _4683_/CLK _4586_/D vssd1 vssd1 vccd1 vccd1 _4586_/Q sky130_fd_sc_hd__dfxtp_1
X_3537_ _4548_/Q _3537_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4548_/D sky130_fd_sc_hd__mux2_1
X_3468_ _4487_/Q _3540_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4487_/D sky130_fd_sc_hd__mux2_1
X_3399_ _4011_/A _3399_/B vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__and2_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2419_ _4063_/A _2961_/A _2837_/A vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2770_ _2950_/S _4546_/Q vssd1 vssd1 vccd1 vccd1 _2770_/X sky130_fd_sc_hd__and2b_1
X_4440_ _4549_/CLK _4440_/D vssd1 vssd1 vccd1 vccd1 _4440_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _4700_/CLK _4371_/D vssd1 vssd1 vccd1 vccd1 _4371_/Q sky130_fd_sc_hd__dfxtp_1
X_3322_ _4382_/Q _4313_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4382_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _4395_/Q _4387_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3253_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2204_ _4590_/Q _3618_/A _4588_/Q vssd1 vssd1 vccd1 vccd1 _2204_/Y sky130_fd_sc_hd__nor3_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3282_/A _3182_/X _3183_/Y _3239_/A vssd1 vssd1 vccd1 vccd1 _3184_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2968_ _3282_/A _2967_/X _3239_/A vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__a21oi_1
X_4638_ _4643_/CLK _4638_/D vssd1 vssd1 vccd1 vccd1 _4638_/Q sky130_fd_sc_hd__dfxtp_1
X_2899_ _2898_/A _2889_/Y _2894_/X _2898_/Y vssd1 vssd1 vccd1 vccd1 _3013_/B sky130_fd_sc_hd__a31o_4
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4569_ _4584_/CLK _4569_/D vssd1 vssd1 vccd1 vccd1 _4569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _4092_/A _4073_/B vssd1 vssd1 vccd1 vccd1 _4103_/C sky130_fd_sc_hd__or2_2
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3871_ _4671_/Q _3936_/A vssd1 vssd1 vccd1 vccd1 _3910_/B sky130_fd_sc_hd__and2b_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2822_ _2661_/S _4547_/Q vssd1 vssd1 vccd1 vccd1 _2822_/X sky130_fd_sc_hd__and2b_1
X_2753_ _4514_/Q _2934_/S _2752_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2684_ _2682_/X _2683_/X _3239_/A _2652_/Y _2656_/Y vssd1 vssd1 vccd1 vccd1 _2685_/B
+ sky130_fd_sc_hd__a2111o_1
X_4423_ _4543_/CLK _4423_/D vssd1 vssd1 vccd1 vccd1 _4423_/Q sky130_fd_sc_hd__dfxtp_1
X_4354_ _4579_/CLK _4354_/D vssd1 vssd1 vccd1 vccd1 _4354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _4368_/Q _4335_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4368_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4285_ _4284_/X _4082_/A _4309_/S vssd1 vssd1 vccd1 vccd1 _4669_/D sky130_fd_sc_hd__mux2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3227_/Y _3228_/Y _3230_/Y _3235_/Y _2389_/A vssd1 vssd1 vccd1 vccd1 _3236_/X
+ sky130_fd_sc_hd__o221a_1
X_3167_ _4369_/Q _4698_/Q _4689_/Q _4417_/Q _3264_/S _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3167_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3098_ _4408_/Q _3140_/S _3097_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _3098_/X sky130_fd_sc_hd__a211o_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout46 _4334_/A1 vssd1 vssd1 vccd1 vccd1 _4314_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout79 _2646_/Y vssd1 vssd1 vccd1 vccd1 _2708_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout57 _2796_/Y vssd1 vssd1 vccd1 vccd1 _3543_/A1 sky130_fd_sc_hd__buf_2
Xfanout68 _2469_/X vssd1 vssd1 vccd1 vccd1 _3564_/A1 sky130_fd_sc_hd__buf_4
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _3938_/A _4267_/A2 _4267_/B1 _3941_/A vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__a22o_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3021_ _2996_/X _2997_/X _3290_/A vssd1 vssd1 vccd1 vccd1 _3021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3923_ _3911_/Y _3922_/X _4204_/B _3910_/X vssd1 vssd1 vccd1 vccd1 _4204_/C sky130_fd_sc_hd__o211ai_4
X_3854_ _4642_/Q _3853_/Y _3854_/S vssd1 vssd1 vccd1 vccd1 _4642_/D sky130_fd_sc_hd__mux2_1
X_2805_ _4579_/Q _2694_/S _2804_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__a211o_1
X_3785_ _4609_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3785_/X sky130_fd_sc_hd__or2_1
X_2736_ _3041_/A _2733_/X _2844_/A vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__o21a_1
X_2667_ _2668_/A1 _2658_/Y _2662_/Y _2664_/Y _2666_/Y vssd1 vssd1 vccd1 vccd1 _3670_/B
+ sky130_fd_sc_hd__a32oi_4
X_4406_ _4695_/CLK _4406_/D vssd1 vssd1 vccd1 vccd1 _4406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout203 _3623_/A vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__clkbuf_16
Xfanout214 _4659_/Q vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__buf_6
X_2598_ _4431_/Q _4423_/Q _2598_/S vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout236 _4616_/Q vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__buf_12
Xfanout225 _3689_/A vssd1 vssd1 vccd1 vccd1 _3716_/A sky130_fd_sc_hd__buf_4
Xfanout247 _2954_/S1 vssd1 vssd1 vccd1 vccd1 _2893_/A sky130_fd_sc_hd__buf_6
X_4337_ _4699_/Q _4337_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4699_/D sky130_fd_sc_hd__mux2_1
X_4268_ _4268_/A _4268_/B _4266_/X vssd1 vssd1 vccd1 vccd1 _4269_/C sky130_fd_sc_hd__or3b_1
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout269 _4438_/Q vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__buf_4
Xfanout258 _2823_/A1 vssd1 vssd1 vccd1 vccd1 _2950_/S sky130_fd_sc_hd__buf_6
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3219_ _4386_/Q _4394_/Q _4410_/Q _4402_/Q _3264_/S _3266_/A1 vssd1 vssd1 vccd1 vccd1
+ _3219_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4199_ _3894_/A _4200_/B _3958_/A vssd1 vssd1 vccd1 vccd1 _4233_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _4578_/Q _3570_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4578_/D sky130_fd_sc_hd__mux2_1
X_2521_ _4349_/Q _3565_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4349_/D sky130_fd_sc_hd__mux2_1
X_2452_ _4532_/Q _2636_/S _2451_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__o211a_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2383_ _4057_/A _3160_/B1 _2382_/X _4645_/Q _2746_/A1 vssd1 vssd1 vccd1 vccd1 _2383_/X
+ sky130_fd_sc_hd__a221o_4
X_4122_ _3921_/X _4118_/Y _4121_/X _4117_/X vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__o211a_1
X_4053_ _2217_/Y _4049_/X _4052_/X _4045_/X vssd1 vssd1 vccd1 vccd1 _4054_/C sky130_fd_sc_hd__o211a_1
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3004_ _3001_/X _3002_/X _3003_/X _3113_/S1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3004_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _4205_/A _3907_/B vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3837_ _4632_/Q _3837_/B vssd1 vssd1 vccd1 vccd1 _3837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3768_ _2432_/X _3283_/A _3713_/A _3766_/X _3767_/Y vssd1 vssd1 vccd1 vccd1 _3768_/X
+ sky130_fd_sc_hd__o221a_1
X_2719_ _2716_/X _2717_/X _2718_/X _2404_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2719_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3699_ _3716_/A _3699_/B vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671_ _4671_/CLK _4671_/D vssd1 vssd1 vccd1 vccd1 _4671_/Q sky130_fd_sc_hd__dfxtp_4
X_3622_ _4619_/Q _3622_/B vssd1 vssd1 vccd1 vccd1 _3988_/C sky130_fd_sc_hd__nand2_1
XFILLER_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3553_ _4563_/Q _4338_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4563_/D sky130_fd_sc_hd__mux2_1
X_2504_ _4469_/Q _4461_/Q _4453_/Q _4445_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2504_/X sky130_fd_sc_hd__mux4_1
X_3484_ _4501_/Q _4312_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4501_/D sky130_fd_sc_hd__mux2_1
X_2435_ _2440_/B _2440_/C vssd1 vssd1 vccd1 vccd1 _2454_/S sky130_fd_sc_hd__nand2_8
XFILLER_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4105_ _3899_/C _3881_/A _3883_/X _4104_/Y vssd1 vssd1 vccd1 vccd1 _4105_/X sky130_fd_sc_hd__a31o_1
X_2366_ _4057_/A _2366_/B _3629_/A vssd1 vssd1 vccd1 vccd1 _2368_/B sky130_fd_sc_hd__or3_4
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2297_ _2473_/B _3387_/B vssd1 vssd1 vccd1 vccd1 _4062_/B sky130_fd_sc_hd__or2_4
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4036_ _4647_/Q _4655_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4037_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2220_ _2292_/B _2360_/B vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__nand2_8
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2984_ _3065_/S _2977_/X _2979_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__a31o_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654_ _4673_/CLK _4654_/D vssd1 vssd1 vccd1 vccd1 _4654_/Q sky130_fd_sc_hd__dfxtp_1
X_3605_ _3608_/A _3633_/A _3624_/C vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__or3b_1
X_4585_ _4689_/CLK _4585_/D vssd1 vssd1 vccd1 vccd1 _4585_/Q sky130_fd_sc_hd__dfxtp_1
X_3536_ _3536_/A _3563_/C _4330_/B vssd1 vssd1 vccd1 vccd1 _3544_/S sky130_fd_sc_hd__and3_4
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3467_ _4486_/Q _3566_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4486_/D sky130_fd_sc_hd__mux2_1
X_3398_ _4046_/B _4003_/A vssd1 vssd1 vccd1 vccd1 _3399_/B sky130_fd_sc_hd__or2_1
X_2418_ _2841_/S _2418_/B vssd1 vssd1 vccd1 vccd1 _2418_/Y sky130_fd_sc_hd__nor2_1
X_2349_ _4437_/Q _2349_/B vssd1 vssd1 vccd1 vccd1 _2352_/B sky130_fd_sc_hd__nand2_4
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4019_ _4647_/Q _4018_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4370_ _4700_/CLK _4370_/D vssd1 vssd1 vccd1 vccd1 _4370_/Q sky130_fd_sc_hd__dfxtp_1
X_3321_ _4381_/Q _4312_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4381_/D sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3252_ _3250_/X _3251_/X _3252_/S vssd1 vssd1 vccd1 vccd1 _3252_/X sky130_fd_sc_hd__mux2_1
X_2203_ input4/X vssd1 vssd1 vccd1 vccd1 _4641_/D sky130_fd_sc_hd__inv_2
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3183_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2967_ _3280_/B1 _2966_/X _2965_/X vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__o21a_1
X_2898_ _2898_/A _2898_/B vssd1 vssd1 vccd1 vccd1 _2898_/Y sky130_fd_sc_hd__nor2_1
X_4637_ _4643_/CLK _4637_/D vssd1 vssd1 vccd1 vccd1 _4637_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ _4570_/CLK _4568_/D vssd1 vssd1 vccd1 vccd1 _4568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _4532_/Q _3564_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4532_/D sky130_fd_sc_hd__mux2_1
X_4499_ _4555_/CLK _4499_/D vssd1 vssd1 vccd1 vccd1 _4499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4673_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3870_ _4177_/A _3960_/B vssd1 vssd1 vccd1 vccd1 _3870_/Y sky130_fd_sc_hd__nand2_4
X_2821_ _3259_/A _2712_/B _3160_/B1 vssd1 vssd1 vccd1 vccd1 _2821_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4549_/CLK sky130_fd_sc_hd__clkbuf_16
X_2752_ _4354_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__and3_1
XFILLER_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4422_ _4574_/CLK _4422_/D vssd1 vssd1 vccd1 vccd1 _4422_/Q sky130_fd_sc_hd__dfxtp_1
X_2683_ _3183_/A _2674_/X _2400_/B _2907_/A vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__o2bb2a_1
X_4353_ _4545_/CLK _4353_/D vssd1 vssd1 vccd1 vccd1 _4353_/Q sky130_fd_sc_hd__dfxtp_1
X_4284_ input5/X _4283_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4284_/X sky130_fd_sc_hd__mux2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _4367_/Q _4334_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4367_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3183_/A _3234_/X _3282_/A vssd1 vssd1 vccd1 vccd1 _3235_/Y sky130_fd_sc_hd__o21ai_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3261_/A _3165_/X _2199_/Y vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3097_ _4400_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _3097_/X sky130_fd_sc_hd__and3_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout47 _3083_/Y vssd1 vssd1 vccd1 vccd1 _4334_/A1 sky130_fd_sc_hd__clkbuf_4
X_3999_ _4261_/B _4245_/C _4261_/A vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__a21oi_2
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout58 _2746_/Y vssd1 vssd1 vccd1 vccd1 _3569_/A1 sky130_fd_sc_hd__buf_4
Xfanout69 _2469_/X vssd1 vssd1 vccd1 vccd1 _3537_/A1 sky130_fd_sc_hd__buf_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4537_/CLK sky130_fd_sc_hd__clkbuf_16
X_3020_ _3018_/X _3019_/X _3020_/S vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3916_/A _3921_/X _3912_/X _3913_/Y vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__o211a_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3853_ _3987_/A _3852_/X _3713_/A vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__a21oi_1
X_2804_ _4523_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2804_/X sky130_fd_sc_hd__and3_1
X_3784_ _4601_/Q _4593_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3784_/X sky130_fd_sc_hd__mux2_1
X_2735_ _2612_/S _2734_/X _2731_/X _2904_/A vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__a211o_1
X_2666_ _2889_/A _2665_/X _2668_/A1 vssd1 vssd1 vccd1 vccd1 _2666_/Y sky130_fd_sc_hd__a21oi_4
X_4405_ _4678_/CLK _4405_/D vssd1 vssd1 vccd1 vccd1 _4405_/Q sky130_fd_sc_hd__dfxtp_1
X_4336_ _4698_/Q _4336_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4698_/D sky130_fd_sc_hd__mux2_1
X_2597_ _2598_/S _4535_/Q _2776_/S1 vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__a21bo_1
Xfanout204 _4675_/Q vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__buf_4
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout237 _4615_/Q vssd1 vssd1 vccd1 vccd1 _2373_/B sky130_fd_sc_hd__buf_12
Xfanout226 _4618_/Q vssd1 vssd1 vccd1 vccd1 _3689_/A sky130_fd_sc_hd__buf_6
Xfanout215 _4658_/Q vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__buf_6
X_4267_ _4643_/Q _4267_/A2 _4267_/B1 _4662_/Q _4238_/A vssd1 vssd1 vccd1 vccd1 _4268_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout248 _4441_/Q vssd1 vssd1 vccd1 vccd1 _2954_/S1 sky130_fd_sc_hd__buf_4
Xfanout259 _2823_/A1 vssd1 vssd1 vccd1 vccd1 _2892_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4198_ _3958_/Y _4200_/A _4172_/A _3870_/Y vssd1 vssd1 vccd1 vccd1 _4198_/Y sky130_fd_sc_hd__o211ai_1
X_3218_ _3261_/A _3213_/X _3217_/X _2199_/Y vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__a211o_2
XFILLER_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _2443_/X _3144_/X _3148_/X _3257_/A1 vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2520_ _2516_/X _2518_/X _2519_/Y _2571_/A vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__o22a_4
X_2451_ _2804_/B _2804_/C _4540_/Q vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__a21o_1
X_2382_ _3185_/A _2385_/A vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__or2_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4121_ _4116_/A _3881_/A _4119_/Y _4140_/B _4266_/B vssd1 vssd1 vccd1 vccd1 _4121_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4052_ _4642_/Q _4042_/X _4048_/X _4051_/X vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__o211a_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _4374_/Q _4678_/Q _3108_/S vssd1 vssd1 vccd1 vccd1 _3003_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_101_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3905_ _3905_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _3905_/X sky130_fd_sc_hd__and2_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3836_ _3836_/A _3836_/B vssd1 vssd1 vccd1 vccd1 _4632_/D sky130_fd_sc_hd__or2_1
X_3767_ _3761_/B _3713_/A _3775_/B1 vssd1 vssd1 vccd1 vccd1 _3767_/Y sky130_fd_sc_hd__a21oi_1
X_2718_ _4433_/Q _4425_/Q _2824_/S vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__mux2_1
X_3698_ _4597_/Q _4329_/S _3697_/Y vssd1 vssd1 vccd1 vccd1 _4597_/D sky130_fd_sc_hd__a21o_1
X_2649_ _2709_/A _2649_/B vssd1 vssd1 vccd1 vccd1 _2652_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _4319_/A _4330_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _4327_/S sky130_fd_sc_hd__and3_4
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670_ _4671_/CLK _4670_/D vssd1 vssd1 vccd1 vccd1 _4670_/Q sky130_fd_sc_hd__dfxtp_4
X_3621_ _3802_/A _3617_/B _3836_/A _3600_/Y vssd1 vssd1 vccd1 vccd1 _4590_/D sky130_fd_sc_hd__a211oi_1
X_3552_ _4562_/Q _4317_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4562_/D sky130_fd_sc_hd__mux2_1
X_2503_ _4549_/Q _4493_/Q _4485_/Q _4477_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2503_/X sky130_fd_sc_hd__mux4_1
X_3483_ _4500_/Q _4320_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4500_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2434_ _3384_/A _2243_/A _2307_/D _2428_/X _2433_/X vssd1 vssd1 vccd1 vccd1 _2440_/C
+ sky130_fd_sc_hd__o311a_4
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2365_ _2860_/C _2400_/C vssd1 vssd1 vccd1 vccd1 _2365_/X sky130_fd_sc_hd__or2_2
X_4104_ _4104_/A _4104_/B vssd1 vssd1 vccd1 vccd1 _4104_/Y sky130_fd_sc_hd__nand2_1
X_2296_ _3832_/B _2331_/A vssd1 vssd1 vccd1 vccd1 _3987_/A sky130_fd_sc_hd__nand2_8
XFILLER_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ _4037_/A _4035_/B vssd1 vssd1 vccd1 vccd1 _4654_/D sky130_fd_sc_hd__and2_1
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3819_ _4626_/Q _4602_/Q _3827_/S vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2983_ _3086_/A _2980_/X _2982_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__o211a_1
X_4653_ _4672_/CLK _4653_/D vssd1 vssd1 vccd1 vccd1 _4653_/Q sky130_fd_sc_hd__dfxtp_1
X_3604_ _3604_/A _3837_/B _4341_/A vssd1 vssd1 vccd1 vccd1 _3604_/Y sky130_fd_sc_hd__nor3b_1
X_4584_ _4584_/CLK _4584_/D vssd1 vssd1 vccd1 vccd1 _4584_/Q sky130_fd_sc_hd__dfxtp_1
X_3535_ _4547_/Q _3571_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4547_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3466_ _4485_/Q _3538_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4485_/D sky130_fd_sc_hd__mux2_1
X_2417_ _3742_/A _3275_/S vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__nor2_1
X_3397_ _3630_/B _3397_/B _3833_/C vssd1 vssd1 vccd1 vccd1 _3397_/Y sky130_fd_sc_hd__nor3_2
X_2348_ _2861_/A _2348_/B _2422_/A vssd1 vssd1 vccd1 vccd1 _2400_/B sky130_fd_sc_hd__or3_2
XFILLER_96_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2279_ _2248_/Y _2250_/X _2277_/X _4091_/B vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__a22o_2
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4018_ _4081_/A _4017_/X _3415_/Y vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3320_ _4380_/Q _4320_/A1 _3327_/S vssd1 vssd1 vccd1 vccd1 _4380_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _4700_/Q _4371_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__mux2_1
X_2202_ input3/X vssd1 vssd1 vccd1 vccd1 _4640_/D sky130_fd_sc_hd__inv_2
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3183_/A _3182_/B _3182_/C vssd1 vssd1 vccd1 vccd1 _3182_/X sky130_fd_sc_hd__or3_1
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2966_ _3716_/B _2963_/B _3770_/S vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__mux2_1
X_2897_ _2895_/X _2896_/X _3261_/A vssd1 vssd1 vccd1 vccd1 _2898_/B sky130_fd_sc_hd__mux2_1
X_4636_ _4692_/CLK _4636_/D vssd1 vssd1 vccd1 vccd1 _4636_/Q sky130_fd_sc_hd__dfxtp_1
X_4567_ _4682_/CLK _4567_/D vssd1 vssd1 vccd1 vccd1 _4567_/Q sky130_fd_sc_hd__dfxtp_1
X_3518_ _3572_/A _3563_/B _4310_/A vssd1 vssd1 vccd1 vccd1 _3526_/S sky130_fd_sc_hd__and3_4
X_4498_ _4684_/CLK _4498_/D vssd1 vssd1 vccd1 vccd1 _4498_/Q sky130_fd_sc_hd__dfxtp_1
X_3449_ _4470_/Q _3539_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4470_/D sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _2655_/B _2819_/Y _2618_/B vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__o21a_1
X_2751_ _2937_/A1 _2748_/X _2750_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2751_/X sky130_fd_sc_hd__o211a_2
X_2682_ _3183_/A _2682_/B _2682_/C vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__or3_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4421_ _4544_/CLK _4421_/D vssd1 vssd1 vccd1 vccd1 _4421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4352_ _4537_/CLK _4352_/D vssd1 vssd1 vccd1 vccd1 _4352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4283_ _3917_/A _4278_/Y _4282_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__a22o_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _4366_/Q _4333_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4366_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3020_/S _3232_/X _3233_/X vssd1 vssd1 vccd1 vccd1 _3234_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3165_ _4529_/Q _4569_/Q _4561_/Q _4505_/Q _3163_/S _3165_/S1 vssd1 vssd1 vccd1 vccd1
+ _3165_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096_ _4392_/Q _4384_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3096_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3998_ _4212_/B _4212_/C _4213_/B vssd1 vssd1 vccd1 vccd1 _4245_/C sky130_fd_sc_hd__a21o_1
Xfanout48 _4333_/A1 vssd1 vssd1 vccd1 vccd1 _4313_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout59 _2746_/Y vssd1 vssd1 vccd1 vccd1 _3542_/A1 sky130_fd_sc_hd__buf_2
X_2949_ _2950_/S _4581_/Q _2893_/A vssd1 vssd1 vccd1 vccd1 _2949_/X sky130_fd_sc_hd__a21bo_1
X_4619_ _4672_/CLK _4619_/D vssd1 vssd1 vccd1 vccd1 _4619_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3921_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3921_/X sky130_fd_sc_hd__and2_1
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3852_ _3581_/C _3832_/B _3629_/B _2302_/A _3623_/C vssd1 vssd1 vccd1 vccd1 _3852_/X
+ sky130_fd_sc_hd__o32a_1
X_2803_ _4515_/Q _2694_/S _2802_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__a211o_1
X_3783_ _3619_/B _3781_/X _3782_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4608_/D sky130_fd_sc_hd__o211a_1
X_2734_ _2725_/X _2733_/X _2841_/S vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__mux2_1
X_2665_ _4472_/Q _4464_/Q _4456_/Q _4448_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2665_/X sky130_fd_sc_hd__mux4_2
X_4404_ _4697_/CLK _4404_/D vssd1 vssd1 vccd1 vccd1 _4404_/Q sky130_fd_sc_hd__dfxtp_1
X_2596_ _2598_/S _4543_/Q vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__and2b_1
Xfanout205 _4674_/Q vssd1 vssd1 vccd1 vccd1 _3933_/B sky130_fd_sc_hd__buf_6
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4335_ _4697_/Q _4335_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4697_/D sky130_fd_sc_hd__mux2_1
Xfanout216 _3917_/A vssd1 vssd1 vccd1 vccd1 _3972_/A sky130_fd_sc_hd__buf_8
Xfanout238 _4589_/Q vssd1 vssd1 vccd1 vccd1 _3618_/A sky130_fd_sc_hd__buf_6
Xfanout227 _3742_/A vssd1 vssd1 vccd1 vccd1 _3770_/S sky130_fd_sc_hd__buf_4
X_4266_ _4266_/A _4266_/B _4266_/C vssd1 vssd1 vccd1 vccd1 _4266_/X sky130_fd_sc_hd__or3_1
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout249 _2776_/S1 vssd1 vssd1 vccd1 vccd1 _2829_/S1 sky130_fd_sc_hd__buf_6
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4197_ _4080_/S _2848_/A _4196_/Y _4081_/A vssd1 vssd1 vccd1 vccd1 _4197_/Y sky130_fd_sc_hd__o211ai_1
X_3217_ _3214_/X _3215_/X _3216_/X _3266_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3217_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _3144_/S _3145_/X _3147_/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__o211a_1
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _3290_/A _3070_/Y _3074_/Y _2652_/A _2389_/A vssd1 vssd1 vccd1 vccd1 _3079_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2450_ _4420_/Q _2636_/S _2449_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__o211a_1
X_2381_ _3185_/A _2385_/A vssd1 vssd1 vccd1 vccd1 _2389_/B sky130_fd_sc_hd__nor2_1
X_4120_ _3881_/A _4119_/Y _4116_/A vssd1 vssd1 vccd1 vccd1 _4140_/B sky130_fd_sc_hd__a21oi_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ _3989_/A _3633_/A _4050_/X _2424_/B _2243_/A vssd1 vssd1 vccd1 vccd1 _4051_/X
+ sky130_fd_sc_hd__o32a_1
Xinput5 io_in[1] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_3002_ _3108_/S _4582_/Q _3113_/S1 vssd1 vssd1 vccd1 vccd1 _3002_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3904_ _3905_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _3904_/Y sky130_fd_sc_hd__nor2_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3835_ _4632_/Q _3607_/B _3835_/S vssd1 vssd1 vccd1 vccd1 _3836_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3766_ _3283_/A _3631_/X _3989_/B _3765_/X vssd1 vssd1 vccd1 vccd1 _3766_/X sky130_fd_sc_hd__o22a_1
X_2717_ _2824_/S _4537_/Q _2404_/A vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__a21bo_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _3739_/B _3695_/X _3696_/X vssd1 vssd1 vccd1 vccd1 _3697_/Y sky130_fd_sc_hd__a21oi_4
X_2648_ _2817_/A _2708_/B vssd1 vssd1 vccd1 vccd1 _2649_/B sky130_fd_sc_hd__nand2_1
X_2579_ _4511_/Q _2932_/S _2578_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__a211o_1
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4318_ _4683_/Q _4338_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4683_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4249_ _3855_/B _3857_/B _3584_/Y _4248_/Y vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3620_ _3614_/Y _3619_/X _3836_/A vssd1 vssd1 vccd1 vccd1 _4589_/D sky130_fd_sc_hd__a21oi_1
X_3551_ _4561_/Q _4316_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4561_/D sky130_fd_sc_hd__mux2_1
X_2502_ _2953_/A _2501_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__a21o_1
X_3482_ _3572_/A _3563_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _3490_/S sky130_fd_sc_hd__and3_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2433_ _3384_/A _2432_/B _2373_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2364_ _2860_/C _2400_/C vssd1 vssd1 vccd1 vccd1 _2364_/Y sky130_fd_sc_hd__nor2_2
X_4103_ _4103_/A _4103_/B _4103_/C vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__and3_1
X_2295_ _3581_/B _2295_/B vssd1 vssd1 vccd1 vccd1 _2331_/A sky130_fd_sc_hd__nand2_8
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _4646_/Q _4654_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4035_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3818_ _3826_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _4625_/D sky130_fd_sc_hd__or2_1
X_3749_ _3749_/A1 _3747_/X _3748_/X _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__a211o_1
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2982_ _4358_/Q _3089_/S _2981_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4652_ _4667_/CLK _4652_/D vssd1 vssd1 vccd1 vccd1 _4652_/Q sky130_fd_sc_hd__dfxtp_1
X_3603_ _4588_/Q _4692_/Q _3836_/A vssd1 vssd1 vccd1 vccd1 _3604_/A sky130_fd_sc_hd__a21o_1
X_4583_ _4679_/CLK _4583_/D vssd1 vssd1 vccd1 vccd1 _4583_/Q sky130_fd_sc_hd__dfxtp_1
X_3534_ _4546_/Q _3570_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4546_/D sky130_fd_sc_hd__mux2_1
X_3465_ _4484_/Q _3564_/A1 _3472_/S vssd1 vssd1 vccd1 vccd1 _4484_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2416_ _3742_/A _3275_/S vssd1 vssd1 vccd1 vccd1 _2511_/A sky130_fd_sc_hd__nand2_4
X_3396_ _3396_/A _3396_/B vssd1 vssd1 vccd1 vccd1 _3833_/C sky130_fd_sc_hd__nand2_1
X_2347_ _4437_/Q _2424_/A _2352_/A vssd1 vssd1 vccd1 vccd1 _2614_/S sky130_fd_sc_hd__or3_4
X_2278_ _2366_/B _3930_/A vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__nand2_8
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4017_ _4667_/Q _3857_/B _4017_/S vssd1 vssd1 vccd1 vccd1 _4017_/X sky130_fd_sc_hd__mux2_2
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _4419_/Q _4691_/Q _3251_/S vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__mux2_1
X_2201_ input2/X vssd1 vssd1 vccd1 vccd1 _4639_/D sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3770_/S _3751_/B _3180_/Y _3020_/S vssd1 vssd1 vccd1 vccd1 _3182_/C sky130_fd_sc_hd__o211a_1
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2965_ _4669_/Q _3278_/A _2425_/Y _2964_/X vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__a211o_1
X_2896_ _4380_/Q _4388_/Q _4404_/Q _4396_/Q _3163_/S _3165_/S1 vssd1 vssd1 vccd1 vccd1
+ _2896_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ _4692_/CLK _4635_/D vssd1 vssd1 vccd1 vccd1 _4635_/Q sky130_fd_sc_hd__dfxtp_1
X_4566_ _4678_/CLK _4566_/D vssd1 vssd1 vccd1 vccd1 _4566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3517_ _4531_/Q _4338_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4531_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4497_ _4553_/CLK _4497_/D vssd1 vssd1 vccd1 vccd1 _4497_/Q sky130_fd_sc_hd__dfxtp_1
X_3448_ _4469_/Q _3538_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4469_/D sky130_fd_sc_hd__mux2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _4432_/Q _3568_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4432_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2750_ _4546_/Q _2934_/S _2749_/X _2931_/C1 vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__a211o_1
X_2681_ _2846_/S _2681_/B vssd1 vssd1 vccd1 vccd1 _2682_/C sky130_fd_sc_hd__nor2_1
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4420_ _4573_/CLK _4420_/D vssd1 vssd1 vccd1 vccd1 _4420_/Q sky130_fd_sc_hd__dfxtp_1
X_4351_ _4543_/CLK _4351_/D vssd1 vssd1 vccd1 vccd1 _4351_/Q sky130_fd_sc_hd__dfxtp_1
X_4282_ _4665_/Q _2367_/Y _3629_/Y _4649_/Q vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__a22o_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _4365_/Q _4332_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4365_/D sky130_fd_sc_hd__mux2_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3770_/S _3230_/B _3224_/Y _3280_/B1 vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__a211o_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3164_ _3161_/X _3162_/X _3163_/X _3165_/S1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3164_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3095_ _3093_/X _3094_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _3095_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout38 _3296_/Y vssd1 vssd1 vccd1 vccd1 _4338_/A1 sky130_fd_sc_hd__buf_4
X_3997_ _4205_/B _4185_/C _4205_/A vssd1 vssd1 vccd1 vccd1 _4212_/C sky130_fd_sc_hd__a21o_1
Xfanout49 _3026_/X vssd1 vssd1 vccd1 vccd1 _4333_/A1 sky130_fd_sc_hd__clkbuf_4
X_2948_ _2950_/S _4357_/Q vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__and2b_1
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4618_ _4671_/CLK _4618_/D vssd1 vssd1 vccd1 vccd1 _4618_/Q sky130_fd_sc_hd__dfxtp_4
X_2879_ _3086_/A _2876_/X _2878_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__o211a_2
X_4549_ _4549_/CLK _4549_/D vssd1 vssd1 vccd1 vccd1 _4549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3920_ _4103_/B _3920_/B vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3851_ _3630_/B _3851_/B _3851_/C _3851_/D vssd1 vssd1 vccd1 vccd1 _3854_/S sky130_fd_sc_hd__and4b_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2802_ _4355_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2802_/X sky130_fd_sc_hd__and3_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3782_ _4608_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__or2_1
X_2733_ _2783_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__and2_1
X_2664_ _3036_/S _2664_/B vssd1 vssd1 vccd1 vccd1 _2664_/Y sky130_fd_sc_hd__nand2_2
X_2595_ _2885_/A _2595_/B vssd1 vssd1 vccd1 vccd1 _2595_/Y sky130_fd_sc_hd__nand2b_1
X_4403_ _4587_/CLK _4403_/D vssd1 vssd1 vccd1 vccd1 _4403_/Q sky130_fd_sc_hd__dfxtp_1
X_4334_ _4696_/Q _4334_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4696_/D sky130_fd_sc_hd__mux2_1
Xfanout217 _4657_/Q vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__buf_4
Xfanout206 _4670_/Q vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout228 _4618_/Q vssd1 vssd1 vccd1 vccd1 _3742_/A sky130_fd_sc_hd__buf_6
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4265_ _4261_/A _3953_/B _4265_/S vssd1 vssd1 vccd1 vccd1 _4266_/C sky130_fd_sc_hd__mux2_1
Xfanout239 _3270_/A vssd1 vssd1 vccd1 vccd1 _2898_/A sky130_fd_sc_hd__buf_12
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4196_ _4184_/Y _4195_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__o21ai_1
X_3216_ _4378_/Q _4682_/Q _3216_/S vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3147_ _4409_/Q _3254_/S _3146_/X _3252_/S vssd1 vssd1 vccd1 vccd1 _3147_/X sky130_fd_sc_hd__a211o_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3078_ _3076_/X _3077_/Y _3050_/X vssd1 vssd1 vccd1 vccd1 _3078_/X sky130_fd_sc_hd__a21bo_1
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ _2380_/A _2380_/B vssd1 vssd1 vccd1 vccd1 _2385_/A sky130_fd_sc_hd__nor2_8
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A _4062_/B _4050_/C vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__or3_1
Xinput6 io_in[2] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3108_/S _4358_/Q vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__and2b_1
XFILLER_49_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _3903_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__or2_2
X_3834_ _3833_/X _3834_/B vssd1 vssd1 vccd1 vccd1 _3835_/S sky130_fd_sc_hd__and2b_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3765_ _3634_/Y _3763_/X _3764_/X _3762_/X vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__o211a_1
X_2716_ _2824_/S _4545_/Q vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__and2b_1
X_3696_ _3731_/A1 _2848_/B _3690_/B _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3696_/X
+ sky130_fd_sc_hd__a221o_2
X_2647_ _2817_/A _2708_/B vssd1 vssd1 vccd1 vccd1 _2709_/A sky130_fd_sc_hd__or2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2578_ _4351_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__and3_1
XFILLER_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4317_ _4682_/Q _4317_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4682_/D sky130_fd_sc_hd__mux2_1
X_4248_ _4248_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _4248_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4179_ _3910_/B _4141_/Y _4177_/A vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__o21ai_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3550_ _4560_/Q _3577_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4560_/D sky130_fd_sc_hd__mux2_1
X_2501_ _4573_/Q _4517_/Q _4509_/Q _4349_/Q _2661_/S _2825_/B2 vssd1 vssd1 vccd1 vccd1
+ _2501_/X sky130_fd_sc_hd__mux4_1
X_3481_ _4499_/Q _3544_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4499_/D sky130_fd_sc_hd__mux2_1
X_2432_ _3384_/A _2432_/B vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__or2_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2363_ _2860_/D _2363_/B vssd1 vssd1 vccd1 vccd1 _2400_/C sky130_fd_sc_hd__or2_2
X_4102_ _4248_/A _4103_/A _3938_/Y _3585_/Y _4057_/X vssd1 vssd1 vccd1 vccd1 _4102_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4033_ _4037_/A _4033_/B vssd1 vssd1 vccd1 vccd1 _4653_/D sky130_fd_sc_hd__and2_1
X_2294_ _3581_/B _2295_/B vssd1 vssd1 vccd1 vccd1 _3634_/B sky130_fd_sc_hd__and2_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3817_ _4625_/Q _4601_/Q _3827_/S vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3748_ _3742_/B _3749_/A1 _2431_/Y _4157_/B vssd1 vssd1 vccd1 vccd1 _3748_/X sky130_fd_sc_hd__a2bb2o_1
X_3679_ _4595_/Q _4329_/S _3678_/Y vssd1 vssd1 vccd1 vccd1 _4595_/D sky130_fd_sc_hd__a21o_1
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4572_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2981_ _4582_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__and3_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4582_/CLK sky130_fd_sc_hd__clkbuf_16
X_4651_ _4651_/CLK _4651_/D vssd1 vssd1 vccd1 vccd1 _4651_/Q sky130_fd_sc_hd__dfxtp_1
X_3602_ _3608_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3837_/B sky130_fd_sc_hd__nor2_1
X_4582_ _4582_/CLK _4582_/D vssd1 vssd1 vccd1 vccd1 _4582_/Q sky130_fd_sc_hd__dfxtp_1
X_3533_ _4545_/Q _3569_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4545_/D sky130_fd_sc_hd__mux2_1
X_3464_ _3536_/A _4319_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _3472_/S sky130_fd_sc_hd__and3_4
X_2415_ _3760_/A _2961_/A vssd1 vssd1 vccd1 vccd1 _2841_/S sky130_fd_sc_hd__nor2_4
X_3395_ _3833_/A _3395_/B _3394_/X vssd1 vssd1 vccd1 vccd1 _3397_/B sky130_fd_sc_hd__or3b_1
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2346_ _4042_/A _2351_/B _2351_/C vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__or3_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2277_ _2366_/B _3930_/A vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__or2_4
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4016_ _4347_/A _4016_/B vssd1 vssd1 vccd1 vccd1 _4646_/D sky130_fd_sc_hd__and2_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4691_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2200_/A vssd1 vssd1 vccd1 vccd1 _4638_/D sky130_fd_sc_hd__inv_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3180_ _3770_/S _3183_/B vssd1 vssd1 vccd1 vccd1 _3180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2964_ _3278_/A _2964_/B _2964_/C _2964_/D vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_14_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4552_/CLK sky130_fd_sc_hd__clkbuf_16
X_2895_ _4364_/Q _4693_/Q _4684_/Q _4412_/Q _2950_/S _2893_/A vssd1 vssd1 vccd1 vccd1
+ _2895_/X sky130_fd_sc_hd__mux4_1
X_4634_ _4702_/CLK _4634_/D vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__dfxtp_1
X_4565_ _4581_/CLK _4565_/D vssd1 vssd1 vccd1 vccd1 _4565_/Q sky130_fd_sc_hd__dfxtp_1
X_3516_ _4530_/Q _4317_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4530_/D sky130_fd_sc_hd__mux2_1
X_4496_ _4552_/CLK _4496_/D vssd1 vssd1 vccd1 vccd1 _4496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3447_ _4468_/Q _3537_/A1 _3454_/S vssd1 vssd1 vccd1 vccd1 _4468_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _4431_/Q _3567_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4431_/D sky130_fd_sc_hd__mux2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _3832_/B _2384_/D vssd1 vssd1 vccd1 vccd1 _2372_/C sky130_fd_sc_hd__nand2_2
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2680_ _4672_/Q _2345_/Y _2846_/S _2679_/Y vssd1 vssd1 vccd1 vccd1 _2682_/B sky130_fd_sc_hd__o211a_1
X_4350_ _4574_/CLK _4350_/D vssd1 vssd1 vccd1 vccd1 _4350_/Q sky130_fd_sc_hd__dfxtp_1
X_3301_ _4364_/Q _4331_/A1 _3308_/S vssd1 vssd1 vccd1 vccd1 _4364_/D sky130_fd_sc_hd__mux2_1
X_4281_ _4280_/X _4063_/A _4309_/S vssd1 vssd1 vccd1 vccd1 _4668_/D sky130_fd_sc_hd__mux2_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4544_/CLK sky130_fd_sc_hd__clkbuf_16
X_3232_ _3933_/B _3231_/X _3232_/S vssd1 vssd1 vccd1 vccd1 _3232_/X sky130_fd_sc_hd__mux2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _4377_/Q _4681_/Q _3163_/S vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3094_ _4697_/Q _4368_/Q _3201_/S vssd1 vssd1 vccd1 vccd1 _3094_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3996_ _4177_/B _4128_/B _4177_/A vssd1 vssd1 vccd1 vccd1 _4185_/C sky130_fd_sc_hd__a21o_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout39 _3296_/Y vssd1 vssd1 vccd1 vccd1 _3580_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2947_ _2953_/A _2947_/B vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__and2_1
X_4617_ _4671_/CLK _4617_/D vssd1 vssd1 vccd1 vccd1 _4617_/Q sky130_fd_sc_hd__dfxtp_1
X_2878_ _4404_/Q _3140_/S _2877_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__a211o_1
X_4548_ _4548_/CLK _4548_/D vssd1 vssd1 vccd1 vccd1 _4548_/Q sky130_fd_sc_hd__dfxtp_1
X_4479_ _4549_/CLK _4479_/D vssd1 vssd1 vccd1 vccd1 _4479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3850_ _2354_/A _4303_/B2 _2350_/A vssd1 vssd1 vccd1 vccd1 _3851_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2801_ _2805_/C1 _2800_/X _2799_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2801_/X sky130_fd_sc_hd__o211a_2
X_3781_ _4600_/Q _4592_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2732_ _2834_/A _3680_/B vssd1 vssd1 vccd1 vccd1 _2733_/B sky130_fd_sc_hd__or2_1
X_2663_ _4552_/Q _4496_/Q _4488_/Q _4480_/Q _2775_/S0 _2775_/S1 vssd1 vssd1 vccd1
+ vccd1 _2664_/B sky130_fd_sc_hd__mux4_2
X_2594_ _4061_/B _2617_/B _2617_/C _2617_/D vssd1 vssd1 vccd1 vccd1 _2595_/B sky130_fd_sc_hd__a31o_1
X_4402_ _4587_/CLK _4402_/D vssd1 vssd1 vccd1 vccd1 _4402_/Q sky130_fd_sc_hd__dfxtp_1
X_4333_ _4695_/Q _4333_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4695_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout229 _3927_/A vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__buf_8
X_4264_ _4264_/A _4264_/B _4264_/C vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__and3_1
Xfanout207 _4071_/A2 vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__buf_6
Xfanout218 _4656_/Q vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__buf_6
X_3215_ _3216_/S _4586_/Q _3266_/A1 vssd1 vssd1 vccd1 vccd1 _3215_/X sky130_fd_sc_hd__a21bo_1
X_4195_ _3934_/A _4673_/Q _4057_/X _4194_/X _4224_/A vssd1 vssd1 vccd1 vccd1 _4195_/X
+ sky130_fd_sc_hd__o311a_1
X_3146_ _4401_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__and3_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3077_ _3936_/A _2860_/C _2364_/Y vssd1 vssd1 vccd1 vccd1 _3077_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3979_ _3955_/X _4228_/A _3953_/X vssd1 vssd1 vccd1 vccd1 _4258_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 io_in[3] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ _4658_/Q _3259_/B vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__or2_1
XFILLER_49_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3902_ _3903_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__nand2_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3833_ _3833_/A _3833_/B _3833_/C _3832_/X vssd1 vssd1 vccd1 vccd1 _3833_/X sky130_fd_sc_hd__or4b_2
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3764_ _3761_/A _3763_/X _3761_/Y _3773_/S vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__a211o_1
X_3695_ _3666_/B1 _3694_/X _2848_/B _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__a2bb2o_2
X_2715_ _2790_/A _2715_/B vssd1 vssd1 vccd1 vccd1 _2715_/Y sky130_fd_sc_hd__nor2_1
X_2646_ _2938_/A1 _2645_/X _2638_/X vssd1 vssd1 vccd1 vccd1 _2646_/Y sky130_fd_sc_hd__o21ai_2
X_2577_ _2937_/A1 _2574_/X _2576_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__o211a_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4316_ _4681_/Q _4316_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4681_/D sky130_fd_sc_hd__mux2_1
X_4247_ _4244_/B _3903_/X _4247_/S vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4178_ _4229_/A _4205_/C _4177_/Y _4176_/X vssd1 vssd1 vccd1 vccd1 _4181_/C sky130_fd_sc_hd__a31o_1
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3103_/X _3104_/Y _3128_/X vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2500_ _2497_/X _2498_/X _2499_/X _2404_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2500_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ _4498_/Q _3543_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4498_/D sky130_fd_sc_hd__mux2_1
X_2431_ _4003_/B _2432_/B vssd1 vssd1 vccd1 vccd1 _2431_/Y sky130_fd_sc_hd__nor2_4
X_2362_ _2473_/B _3991_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _2618_/B sky130_fd_sc_hd__or3_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ _3936_/A _4267_/A2 _4267_/B1 _3972_/A vssd1 vssd1 vccd1 vccd1 _4123_/B sky130_fd_sc_hd__a22o_1
X_2293_ _2293_/A _2293_/B _3991_/B vssd1 vssd1 vccd1 vccd1 _2354_/B sky130_fd_sc_hd__or3_1
X_4032_ _4645_/Q _4653_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4033_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3816_ _3826_/A _3816_/B vssd1 vssd1 vccd1 vccd1 _4624_/D sky130_fd_sc_hd__or2_1
X_3747_ _3989_/B _3746_/X _4157_/B _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3678_ _3739_/B _3676_/X _3677_/X vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__a21oi_4
X_2629_ _2571_/A _2626_/X _2628_/Y _2625_/Y vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__o31a_2
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2980_ _4678_/Q _4374_/Q _3089_/S vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4667_/CLK _4650_/D vssd1 vssd1 vccd1 vccd1 _4650_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 io_in[6] vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__clkbuf_2
X_3601_ _4011_/A _3601_/B _2233_/C vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__or3b_1
X_4581_ _4581_/CLK _4581_/D vssd1 vssd1 vccd1 vccd1 _4581_/Q sky130_fd_sc_hd__dfxtp_1
X_3532_ _4544_/Q _3568_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4544_/D sky130_fd_sc_hd__mux2_1
X_3463_ _4483_/Q _3544_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4483_/D sky130_fd_sc_hd__mux2_1
X_2414_ _2414_/A _2414_/B vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__nand2_4
X_3394_ _4050_/A _2190_/Y _3991_/B _2351_/C vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2345_ _2349_/B _3630_/A vssd1 vssd1 vccd1 vccd1 _2345_/Y sky130_fd_sc_hd__nand2_4
X_2276_ _2373_/C _3930_/A vssd1 vssd1 vccd1 vccd1 _2384_/C sky130_fd_sc_hd__nor2_2
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4015_ _4646_/Q _4014_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2963_ _3174_/A _2963_/B vssd1 vssd1 vccd1 vccd1 _2964_/D sky130_fd_sc_hd__or2_1
X_4702_ _4702_/CLK _4702_/D vssd1 vssd1 vccd1 vccd1 _4702_/Q sky130_fd_sc_hd__dfxtp_1
X_2894_ _2954_/S1 _2891_/Y _2893_/Y _2889_/A vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__a211o_1
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4633_ _4702_/CLK _4633_/D vssd1 vssd1 vccd1 vccd1 _4633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _4580_/CLK _4564_/D vssd1 vssd1 vccd1 vccd1 _4564_/Q sky130_fd_sc_hd__dfxtp_1
X_3515_ _4529_/Q _4316_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4529_/D sky130_fd_sc_hd__mux2_1
X_4495_ _4549_/CLK _4495_/D vssd1 vssd1 vccd1 vccd1 _4495_/Q sky130_fd_sc_hd__dfxtp_1
X_3446_ _3536_/A _3563_/C _3446_/C vssd1 vssd1 vccd1 vccd1 _3454_/S sky130_fd_sc_hd__and3_4
XFILLER_69_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _4430_/Q _3566_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4430_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2328_ _4003_/B _4238_/A vssd1 vssd1 vccd1 vccd1 _3390_/B sky130_fd_sc_hd__nor2_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2259_ _3993_/A _2384_/B vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__nand2_8
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ _4330_/A _3563_/C _4330_/B vssd1 vssd1 vccd1 vccd1 _3308_/S sky130_fd_sc_hd__and3_4
X_4280_ input1/X _4279_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4280_/X sky130_fd_sc_hd__mux2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3223_/X _3230_/B _3231_/S vssd1 vssd1 vccd1 vccd1 _3231_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3264_/S _4585_/Q _3113_/S1 vssd1 vssd1 vccd1 vccd1 _3162_/X sky130_fd_sc_hd__a21bo_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _4416_/Q _4688_/Q _3201_/S vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3995_ _4127_/B _4127_/C _4127_/A vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__o21ai_2
X_2946_ _4525_/Q _4565_/Q _4557_/Q _4501_/Q _2950_/S _2893_/A vssd1 vssd1 vccd1 vccd1
+ _2947_/B sky130_fd_sc_hd__mux4_1
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2877_ _4396_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__and3_1
X_4616_ _4671_/CLK _4616_/D vssd1 vssd1 vccd1 vccd1 _4616_/Q sky130_fd_sc_hd__dfxtp_1
X_4547_ _4573_/CLK _4547_/D vssd1 vssd1 vccd1 vccd1 _4547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4478_ _4549_/CLK _4478_/D vssd1 vssd1 vccd1 vccd1 _4478_/Q sky130_fd_sc_hd__dfxtp_1
X_3429_ _4452_/Q _3537_/A1 _3436_/S vssd1 vssd1 vccd1 vccd1 _4452_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2800_ _4427_/Q _4435_/Q _2800_/S vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _3619_/B _3778_/X _3779_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4607_/D sky130_fd_sc_hd__o211a_1
X_2731_ _2348_/B _2729_/X _2730_/X _3276_/B vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__o211a_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ _4681_/CLK _4401_/D vssd1 vssd1 vccd1 vccd1 _4401_/Q sky130_fd_sc_hd__dfxtp_1
X_2662_ _2659_/X _2660_/X _2661_/X _2825_/B2 _2549_/A vssd1 vssd1 vccd1 vccd1 _2662_/Y
+ sky130_fd_sc_hd__o221ai_4
X_2593_ _4061_/B _2617_/B _2617_/C _2617_/D vssd1 vssd1 vccd1 vccd1 _2885_/A sky130_fd_sc_hd__and4_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _4694_/Q _4332_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4694_/D sky130_fd_sc_hd__mux2_1
X_4263_ _3903_/X _4244_/B _4263_/S vssd1 vssd1 vccd1 vccd1 _4264_/C sky130_fd_sc_hd__mux2_1
Xfanout208 _4669_/Q vssd1 vssd1 vccd1 vccd1 _4071_/A2 sky130_fd_sc_hd__buf_4
Xfanout219 _4656_/Q vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__buf_4
XFILLER_101_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3214_ _3216_/S _4362_/Q vssd1 vssd1 vccd1 vccd1 _3214_/X sky130_fd_sc_hd__and2b_1
X_4194_ _2225_/Y _4212_/C _4185_/Y _4193_/X vssd1 vssd1 vccd1 vccd1 _4194_/X sky130_fd_sc_hd__a31o_1
X_3145_ _4393_/Q _4385_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _2655_/B _3070_/Y _3075_/Y _2860_/C vssd1 vssd1 vccd1 vccd1 _3076_/X sky130_fd_sc_hd__a211o_1
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _3958_/A _3977_/X _3954_/Y _4233_/A vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__a211o_1
X_2929_ _2937_/C1 _2926_/X _2928_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput8 io_in[4] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3901_ _3927_/B _3900_/X _3891_/X _4104_/A vssd1 vssd1 vccd1 vccd1 _3993_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3832_ _4050_/A _3832_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _3832_/X sky130_fd_sc_hd__or3_2
X_3763_ _3760_/A _3283_/A _3760_/Y vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__a21o_1
X_3694_ _3754_/A1 _3692_/Y _3693_/X _3691_/X vssd1 vssd1 vccd1 vccd1 _3694_/X sky130_fd_sc_hd__o211a_1
X_2714_ _2885_/A _2885_/B _2848_/A vssd1 vssd1 vccd1 vccd1 _2715_/B sky130_fd_sc_hd__a21oi_1
X_2645_ _2641_/X _2644_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4315_ _4680_/Q _4335_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4680_/D sky130_fd_sc_hd__mux2_1
X_2576_ _4543_/Q _2811_/S _2575_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4246_ _4246_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4177_/A _4177_/B _4177_/C vssd1 vssd1 vccd1 vccd1 _4177_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _2652_/A _3102_/Y _3105_/Y _2655_/Y _3127_/Y vssd1 vssd1 vccd1 vccd1 _3128_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _4696_/Q _4367_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3059_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _3384_/A _4620_/Q _3623_/C _3622_/B vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__or4b_1
X_2361_ _2473_/B _3991_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _2363_/B sky130_fd_sc_hd__nor3_4
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4100_ _4099_/X _4132_/B vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__and2b_1
X_2292_ _2360_/B _2292_/B vssd1 vssd1 vccd1 vccd1 _3991_/B sky130_fd_sc_hd__nand2b_4
X_4031_ _4037_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _4652_/D sky130_fd_sc_hd__and2_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3815_ _4624_/Q _4600_/Q _3827_/S vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__mux2_1
X_3746_ _4688_/Q _3762_/B _3691_/C _3745_/X vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__o31a_1
X_3677_ _3731_/A1 _2885_/B _3671_/B _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3677_/X
+ sky130_fd_sc_hd__a221o_2
X_2628_ _2745_/C vssd1 vssd1 vccd1 vccd1 _2628_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2559_ _3938_/B _2348_/B _2558_/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2559_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _4229_/A _4261_/C vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput11 io_in[7] vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__clkbuf_2
X_3600_ _3802_/A _3799_/S _3617_/B vssd1 vssd1 vccd1 vccd1 _3600_/Y sky130_fd_sc_hd__a21oi_1
X_4580_ _4580_/CLK _4580_/D vssd1 vssd1 vccd1 vccd1 _4580_/Q sky130_fd_sc_hd__dfxtp_1
X_3531_ _4543_/Q _3567_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4543_/D sky130_fd_sc_hd__mux2_1
X_3462_ _4482_/Q _3543_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4482_/D sky130_fd_sc_hd__mux2_1
X_3393_ _4632_/Q _3602_/B vssd1 vssd1 vccd1 vccd1 _3395_/B sky130_fd_sc_hd__nor2_1
X_2413_ _2414_/A _2414_/B vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__and2_4
X_2344_ _2349_/B _3630_/A vssd1 vssd1 vccd1 vccd1 _2422_/A sky130_fd_sc_hd__and2_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2275_ _2217_/B _2349_/B _3990_/A _2274_/X vssd1 vssd1 vccd1 vccd1 _2275_/X sky130_fd_sc_hd__a31o_1
X_4014_ _4081_/A _4013_/X _3411_/Y vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _4686_/Q _3762_/B _3691_/C _3728_/X vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__o31a_1
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2962_ _2962_/A _3119_/A vssd1 vssd1 vccd1 vccd1 _2963_/B sky130_fd_sc_hd__and2_1
X_4701_ _4702_/CLK _4701_/D vssd1 vssd1 vccd1 vccd1 _4701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ _4702_/CLK _4632_/D vssd1 vssd1 vccd1 vccd1 _4632_/Q sky130_fd_sc_hd__dfxtp_4
X_2893_ _2893_/A _2893_/B vssd1 vssd1 vccd1 vccd1 _2893_/Y sky130_fd_sc_hd__nor2_1
X_4563_ _4683_/CLK _4563_/D vssd1 vssd1 vccd1 vccd1 _4563_/Q sky130_fd_sc_hd__dfxtp_1
X_4494_ _4549_/CLK _4494_/D vssd1 vssd1 vccd1 vccd1 _4494_/Q sky130_fd_sc_hd__dfxtp_1
X_3514_ _4528_/Q _3577_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4528_/D sky130_fd_sc_hd__mux2_1
X_3445_ _4467_/Q _3544_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4467_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _4429_/Q _3565_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4429_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2233_/Y _2424_/B _2327_/C vssd1 vssd1 vccd1 vccd1 _2327_/Y sky130_fd_sc_hd__nand3b_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2258_ _3993_/A _4638_/Q _3993_/B vssd1 vssd1 vccd1 vccd1 _2263_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2189_ _4642_/Q vssd1 vssd1 vccd1 vccd1 _2189_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3230_ _3230_/A _3230_/B vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__nor2_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3163_/S _4361_/Q vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__and2b_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _3086_/A _3089_/X _3091_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _3092_/X sky130_fd_sc_hd__o211a_1
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3994_ _4103_/B _4103_/C _4103_/A vssd1 vssd1 vccd1 vccd1 _4127_/C sky130_fd_sc_hd__a21oi_2
XFILLER_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _3287_/A _2995_/A vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__xor2_1
X_2876_ _4388_/Q _4380_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__mux2_1
X_4615_ _4671_/CLK _4615_/D vssd1 vssd1 vccd1 vccd1 _4615_/Q sky130_fd_sc_hd__dfxtp_4
X_4546_ _4572_/CLK _4546_/D vssd1 vssd1 vccd1 vccd1 _4546_/Q sky130_fd_sc_hd__dfxtp_1
X_4477_ _4549_/CLK _4477_/D vssd1 vssd1 vccd1 vccd1 _4477_/Q sky130_fd_sc_hd__dfxtp_1
X_3428_ _3563_/B _4319_/A _3446_/C vssd1 vssd1 vccd1 vccd1 _3436_/S sky130_fd_sc_hd__and3_4
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3359_ _4414_/Q _4333_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4414_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _4673_/Q _2837_/A vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__or2_1
X_2661_ _4432_/Q _4424_/Q _2661_/S vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__mux2_2
X_4400_ _4582_/CLK _4400_/D vssd1 vssd1 vccd1 vccd1 _4400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2592_ _3257_/A1 _2586_/X _2590_/X _2577_/X _2582_/X vssd1 vssd1 vccd1 vccd1 _2617_/D
+ sky130_fd_sc_hd__o32ai_4
X_4331_ _4693_/Q _4331_/A1 _4338_/S vssd1 vssd1 vccd1 vccd1 _4693_/D sky130_fd_sc_hd__mux2_1
Xfanout209 _4668_/Q vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__buf_6
X_4262_ _4262_/A _4262_/B _4262_/C vssd1 vssd1 vccd1 vccd1 _4262_/X sky130_fd_sc_hd__or3_1
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _4530_/Q _4570_/Q _4562_/Q _4506_/Q _3216_/S _3266_/A1 vssd1 vssd1 vccd1 vccd1
+ _3213_/X sky130_fd_sc_hd__mux4_1
X_4193_ _4215_/A _4187_/X _4192_/X vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3142_/X _3143_/X _3144_/S vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3075_ _3074_/A _3102_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3075_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3977_ _3870_/Y _4172_/A _4200_/A _3958_/Y vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _4525_/Q _2934_/S _2927_/X _2937_/A1 vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__a211o_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2859_/A _3299_/B vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__nor2_4
X_4529_ _4683_/CLK _4529_/D vssd1 vssd1 vccd1 vccd1 _4529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_in[5] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _4244_/B _4216_/B _3899_/X _3891_/X vssd1 vssd1 vccd1 vccd1 _3900_/X sky130_fd_sc_hd__o31a_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3831_ _2360_/B _2290_/B _3384_/B _2357_/Y vssd1 vssd1 vccd1 vccd1 _3990_/C sky130_fd_sc_hd__a211o_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3762_ _4690_/Q _3762_/B _4017_/S vssd1 vssd1 vccd1 vccd1 _3762_/X sky130_fd_sc_hd__or3_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3693_ _3727_/S _3692_/Y _3690_/Y _3720_/S vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__a211o_1
X_2713_ _2885_/A _2885_/B _2848_/A vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__and3_1
X_2644_ _2642_/X _2643_/X _2644_/S vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__mux2_1
X_2575_ _4535_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__and3_1
X_4314_ _4679_/Q _4314_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4679_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4245_ _4261_/A _4261_/B _4245_/C vssd1 vssd1 vccd1 vccd1 _4246_/B sky130_fd_sc_hd__and3_1
X_4176_ _3961_/A _4139_/X _4200_/B _4235_/A vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__o211a_1
X_3127_ _3239_/A _3127_/B vssd1 vssd1 vccd1 vccd1 _3127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _3194_/C1 _3053_/X _3055_/X _3057_/X _3249_/C1 vssd1 vssd1 vccd1 vccd1 _3058_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2360_ _2360_/A _2360_/B _2473_/B _2473_/C vssd1 vssd1 vccd1 vccd1 _2712_/B sky130_fd_sc_hd__or4_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2291_ _3608_/A _4046_/A _2290_/Y vssd1 vssd1 vccd1 vccd1 _2293_/B sky130_fd_sc_hd__or3b_1
X_4030_ _4644_/Q _4652_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4031_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3814_ _3828_/A _3814_/B vssd1 vssd1 vccd1 vccd1 _4623_/D sky130_fd_sc_hd__nand2_1
X_3745_ _3634_/Y _3743_/Y _3744_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3745_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _3666_/B1 _3675_/X _2885_/B _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3676_/X sky130_fd_sc_hd__a2bb2o_2
X_2627_ _4484_/Q _4485_/Q _4486_/Q _4487_/Q vssd1 vssd1 vccd1 vccd1 _2745_/C sky130_fd_sc_hd__or4_4
X_2558_ _2837_/A _2607_/A _2558_/C vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__and3_1
X_2489_ _4453_/Q _2699_/S _2488_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__a211o_1
X_4228_ _4228_/A _4228_/B _4228_/C vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__and3_1
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4159_ _4177_/A _4177_/B _4128_/B _4158_/Y vssd1 vssd1 vccd1 vccd1 _4159_/X sky130_fd_sc_hd__a31o_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 io_in[8] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
X_3530_ _4542_/Q _3566_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4542_/D sky130_fd_sc_hd__mux2_1
X_3461_ _4481_/Q _3542_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4481_/D sky130_fd_sc_hd__mux2_1
X_3392_ _2307_/D _2310_/X _3391_/B _2354_/A vssd1 vssd1 vccd1 vccd1 _3630_/B sky130_fd_sc_hd__a31oi_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2412_ _2412_/A _2412_/B vssd1 vssd1 vccd1 vccd1 _2414_/B sky130_fd_sc_hd__nand2_2
XFILLER_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2343_ _4437_/Q _2350_/A vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__nor2_4
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2274_ _2274_/A _4437_/Q _3989_/A vssd1 vssd1 vccd1 vccd1 _2274_/X sky130_fd_sc_hd__and3_1
X_4013_ _4666_/Q _3933_/B _4013_/S vssd1 vssd1 vccd1 vccd1 _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4651_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3728_ _3754_/A1 _3726_/Y _3727_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__o22a_1
X_3659_ _3731_/A1 _2617_/C _3653_/B _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3659_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2961_ _2961_/A _3013_/A _3013_/B _3013_/C vssd1 vssd1 vccd1 vccd1 _3119_/A sky130_fd_sc_hd__or4_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4700_/CLK _4700_/D vssd1 vssd1 vccd1 vccd1 _4700_/Q sky130_fd_sc_hd__dfxtp_1
X_4631_ _4702_/CLK _4631_/D vssd1 vssd1 vccd1 vccd1 _4631_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2892_ _4372_/Q _4676_/Q _2892_/S vssd1 vssd1 vccd1 vccd1 _2893_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4562_ _4570_/CLK _4562_/D vssd1 vssd1 vccd1 vccd1 _4562_/Q sky130_fd_sc_hd__dfxtp_1
X_4493_ _4552_/CLK _4493_/D vssd1 vssd1 vccd1 vccd1 _4493_/Q sky130_fd_sc_hd__dfxtp_1
X_3513_ _4527_/Q _4314_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4527_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4574_/CLK sky130_fd_sc_hd__clkbuf_16
X_3444_ _4466_/Q _3543_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4466_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _4428_/Q _3564_/A1 _3382_/S vssd1 vssd1 vccd1 vccd1 _4428_/D sky130_fd_sc_hd__mux2_1
X_2326_ _3385_/B _2354_/A _3581_/B vssd1 vssd1 vccd1 vccd1 _2327_/C sky130_fd_sc_hd__or3b_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _2366_/B _4640_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _2263_/C sky130_fd_sc_hd__and3_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2188_ _4588_/Q vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__inv_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3934_/A _3259_/B _3160_/B1 _3159_/X vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__o211a_1
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3091_ _4360_/Q _3089_/S _3090_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__a211o_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3993_ _3993_/A _3993_/B _3993_/C _3993_/D vssd1 vssd1 vccd1 vccd1 _3993_/X sky130_fd_sc_hd__or4_1
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2944_ _4657_/Q _3259_/B _3160_/B1 vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__o21ai_1
X_2875_ _3144_/S _2874_/X _2873_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__o211a_2
X_4614_ _4692_/CLK _4614_/D vssd1 vssd1 vccd1 vccd1 _4614_/Q sky130_fd_sc_hd__dfxtp_1
X_4545_ _4545_/CLK _4545_/D vssd1 vssd1 vccd1 vccd1 _4545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4476_ _4553_/CLK _4476_/D vssd1 vssd1 vccd1 vccd1 _4476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3427_ _4451_/Q _3571_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4451_/D sky130_fd_sc_hd__mux2_1
X_3358_ _4413_/Q _4332_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4413_/D sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _4046_/B _3991_/B vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__nor2_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3289_ _2655_/B _3290_/B _3288_/X _3259_/B vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__o211a_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2660_ _2661_/S _4536_/Q _2825_/B2 vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__a21bo_1
X_2591_ _2938_/A1 _2586_/X _2590_/X _2577_/X _2582_/X vssd1 vssd1 vccd1 vccd1 _2591_/X
+ sky130_fd_sc_hd__o32a_4
X_4330_ _4330_/A _4330_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _4338_/S sky130_fd_sc_hd__and3_4
X_4261_ _4261_/A _4261_/B _4261_/C vssd1 vssd1 vccd1 vccd1 _4262_/C sky130_fd_sc_hd__and3_1
X_3212_ _3212_/A _3283_/A vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__xnor2_1
X_4192_ _4104_/A _4217_/A _4188_/X _4191_/X vssd1 vssd1 vccd1 vccd1 _4192_/X sky130_fd_sc_hd__a31o_1
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3143_ _4417_/Q _4689_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3074_ _3074_/A _3102_/A vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3976_ _3962_/Y _3975_/Y _3870_/Y _3961_/A vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__o211ai_4
X_2927_ _4565_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__and3_1
X_2858_ _2858_/A _3298_/B vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__nor2_8
X_2789_ _3020_/S _2784_/X _2787_/X _2788_/X vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__a22o_1
X_4528_ _4570_/CLK _4528_/D vssd1 vssd1 vccd1 vccd1 _4528_/Q sky130_fd_sc_hd__dfxtp_1
X_4459_ _4555_/CLK _4459_/D vssd1 vssd1 vccd1 vccd1 _4459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3608_/A _3602_/B _3829_/X _2274_/A vssd1 vssd1 vccd1 vccd1 _4631_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3761_ _3761_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__nor2_1
X_2712_ _3934_/A _2712_/B vssd1 vssd1 vccd1 vccd1 _2712_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3692_ _3716_/A _2848_/B _3689_/Y vssd1 vssd1 vccd1 vccd1 _3692_/Y sky130_fd_sc_hd__o21ai_1
X_2643_ _4448_/Q _4456_/Q _2761_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2574_ _4423_/Q _4431_/Q _2811_/S vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4313_ _4678_/Q _4313_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4678_/D sky130_fd_sc_hd__mux2_1
X_4244_ _4244_/A _4244_/B vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4175_ _3960_/B _4139_/X _4177_/A vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__o21ai_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3126_ _3282_/A _3126_/B _3126_/C vssd1 vssd1 vccd1 vccd1 _3127_/B sky130_fd_sc_hd__and3_1
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3057_ _3255_/S _3056_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3057_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _3959_/A _4188_/B vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2290_ _3622_/B _2290_/B vssd1 vssd1 vccd1 vccd1 _2290_/Y sky130_fd_sc_hd__nand2_2
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _2185_/Y _2186_/Y _3827_/S vssd1 vssd1 vccd1 vccd1 _3814_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _3742_/B _3743_/Y _3771_/S vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__mux2_1
X_3675_ _3754_/A1 _3673_/Y _3674_/X _3672_/X vssd1 vssd1 vccd1 vccd1 _3675_/X sky130_fd_sc_hd__o211a_1
X_2626_ _4484_/Q _4485_/Q _4486_/Q _4487_/Q vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__o31a_1
XFILLER_99_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2557_ _3275_/S _3643_/B _3652_/B vssd1 vssd1 vccd1 vccd1 _2558_/C sky130_fd_sc_hd__a21o_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _4445_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__and3_1
X_4227_ _3954_/Y _4233_/A _3958_/A _3977_/X vssd1 vssd1 vccd1 vccd1 _4228_/C sky130_fd_sc_hd__o211ai_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _4229_/A _4185_/C vssd1 vssd1 vccd1 vccd1 _4158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _4116_/C _4089_/B vssd1 vssd1 vccd1 vccd1 _4093_/S sky130_fd_sc_hd__and2_1
X_3109_ _3106_/X _3107_/X _3108_/X _3113_/S1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3109_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 io_in[9] vssd1 vssd1 vccd1 vccd1 _2200_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3460_ _4480_/Q _3541_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4480_/D sky130_fd_sc_hd__mux2_1
X_3391_ _4050_/A _3391_/B vssd1 vssd1 vccd1 vccd1 _3833_/B sky130_fd_sc_hd__nor2_1
X_2411_ _2409_/X _2410_/X _2549_/A vssd1 vssd1 vccd1 vccd1 _2412_/B sky130_fd_sc_hd__mux2_1
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2342_ _3581_/B _2351_/B _2351_/C vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__or3_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4012_ _4645_/Q _4019_/S _4011_/Y _4347_/A vssd1 vssd1 vccd1 vccd1 _4645_/D sky130_fd_sc_hd__o211a_1
X_2273_ _3990_/A vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__inv_2
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3727_ _3725_/B _3726_/Y _3727_/S vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__mux2_1
X_3658_ _3666_/B1 _3657_/X _2617_/C _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__a2bb2o_1
X_3589_ _3628_/A _3630_/C _3588_/X _4062_/A vssd1 vssd1 vccd1 vccd1 _3589_/X sky130_fd_sc_hd__o31a_1
X_2609_ _3643_/B _3652_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _2610_/B sky130_fd_sc_hd__a21oi_1
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout190 _3761_/A vssd1 vssd1 vccd1 vccd1 _3771_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2960_ _2414_/Y _2904_/B _2901_/B _3716_/B vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__a31o_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _2891_/A vssd1 vssd1 vccd1 vccd1 _2891_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ _4630_/CLK _4630_/D vssd1 vssd1 vccd1 vccd1 _4630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4561_ _4584_/CLK _4561_/D vssd1 vssd1 vccd1 vccd1 _4561_/Q sky130_fd_sc_hd__dfxtp_1
X_3512_ _4526_/Q _4313_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4526_/D sky130_fd_sc_hd__mux2_1
X_4492_ _4553_/CLK _4492_/D vssd1 vssd1 vccd1 vccd1 _4492_/Q sky130_fd_sc_hd__dfxtp_1
X_3443_ _4465_/Q _3542_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4465_/D sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3563_/B _4310_/A _3563_/C vssd1 vssd1 vccd1 vccd1 _3382_/S sky130_fd_sc_hd__and3_4
X_2325_ _2354_/A _2425_/A vssd1 vssd1 vccd1 vccd1 _2424_/B sky130_fd_sc_hd__or2_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _2373_/C _3585_/B vssd1 vssd1 vccd1 vccd1 _3930_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2187_ _4590_/Q vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__clkinv_4
XFILLER_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ _4584_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _3090_/X sky130_fd_sc_hd__and3_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3992_ _3846_/B _3987_/Y _3991_/Y _3987_/A _3990_/X vssd1 vssd1 vccd1 vccd1 _3992_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2943_ _2655_/B _2942_/X _3259_/B vssd1 vssd1 vccd1 vccd1 _2943_/X sky130_fd_sc_hd__o21a_1
X_2874_ _4693_/Q _4364_/Q _2932_/S vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4613_ _4613_/CLK _4613_/D vssd1 vssd1 vccd1 vccd1 _4613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4544_ _4544_/CLK _4544_/D vssd1 vssd1 vccd1 vccd1 _4544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4475_ _4555_/CLK _4475_/D vssd1 vssd1 vccd1 vccd1 _4475_/Q sky130_fd_sc_hd__dfxtp_1
X_3426_ _4450_/Q _3570_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4450_/D sky130_fd_sc_hd__mux2_1
X_3357_ _4412_/Q _4331_/A1 _3364_/S vssd1 vssd1 vccd1 vccd1 _4412_/D sky130_fd_sc_hd__mux2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _3989_/A _2307_/X _2354_/B vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__o21ai_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3288_ _3288_/A _3288_/B _3288_/C vssd1 vssd1 vccd1 vccd1 _3288_/X sky130_fd_sc_hd__or3_1
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2239_ _2190_/Y _4046_/A _3989_/A vssd1 vssd1 vccd1 vccd1 _2243_/A sky130_fd_sc_hd__a21o_2
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2814_/A1 _2587_/X _2589_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__o211a_2
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _3926_/X _4260_/B _4260_/C vssd1 vssd1 vccd1 vccd1 _4269_/B sky130_fd_sc_hd__and3b_1
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4221_/A _4191_/B _4190_/X vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__or3b_1
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3211_ _3288_/A _3211_/B vssd1 vssd1 vccd1 vccd1 _3211_/Y sky130_fd_sc_hd__nand2_1
X_3142_ _4698_/Q _4369_/Q _3254_/S vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3073_ _3209_/A _3209_/B vssd1 vssd1 vccd1 vccd1 _3102_/A sky130_fd_sc_hd__or2_2
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3975_ _3973_/A _3974_/Y _3962_/Y _3963_/X vssd1 vssd1 vccd1 vccd1 _3975_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2926_ _4557_/Q _2934_/S _2925_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2926_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2857_ _4355_/Q _3571_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4355_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2788_ _3933_/B _2614_/S _2846_/S vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4527_ _4682_/CLK _4527_/D vssd1 vssd1 vccd1 vccd1 _4527_/Q sky130_fd_sc_hd__dfxtp_1
X_4458_ _4553_/CLK _4458_/D vssd1 vssd1 vccd1 vccd1 _4458_/Q sky130_fd_sc_hd__dfxtp_1
X_3409_ _3417_/S _3408_/X _3849_/A vssd1 vssd1 vccd1 vccd1 _3409_/Y sky130_fd_sc_hd__a21oi_4
X_4389_ _4678_/CLK _4389_/D vssd1 vssd1 vccd1 vccd1 _4389_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3760_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3760_/Y sky130_fd_sc_hd__nor2_1
X_2711_ _2472_/Y _2710_/Y _2618_/B vssd1 vssd1 vccd1 vccd1 _2711_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3691_ _4490_/Q _3762_/B _3691_/C vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__or3_1
X_2642_ _4464_/Q _4472_/Q _2761_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2573_ _4350_/Q _3566_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4350_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _4677_/Q _4312_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4677_/D sky130_fd_sc_hd__mux2_1
X_4243_ _4662_/Q _4242_/Y _4272_/S vssd1 vssd1 vccd1 vccd1 _4662_/D sky130_fd_sc_hd__mux2_1
X_4174_ _4204_/C _4260_/B _4173_/X _4167_/B _4123_/A vssd1 vssd1 vccd1 vccd1 _4181_/B
+ sky130_fd_sc_hd__a311o_1
X_3125_ _3760_/A _3742_/B _3124_/Y _3280_/B1 vssd1 vssd1 vccd1 vccd1 _3126_/C sky130_fd_sc_hd__a211o_1
X_3056_ _4567_/Q _4527_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3056_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _3958_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3889_ _3956_/A _4217_/A vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__and2_1
X_2909_ _4668_/Q _2907_/A _3020_/S _2908_/Y vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__a211o_1
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3812_ _2292_/B _4270_/A _3812_/S vssd1 vssd1 vccd1 vccd1 _4622_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3743_ _3742_/A _4157_/B _3742_/Y vssd1 vssd1 vccd1 vccd1 _3743_/Y sky130_fd_sc_hd__o21ai_1
X_3674_ _3771_/S _3673_/Y _3671_/Y _3720_/S vssd1 vssd1 vccd1 vccd1 _3674_/X sky130_fd_sc_hd__a211o_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2625_ _2618_/Y _2621_/Y _2624_/X vssd1 vssd1 vccd1 vccd1 _2625_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2556_ _3653_/B _2961_/A _2513_/B vssd1 vssd1 vccd1 vccd1 _2607_/A sky130_fd_sc_hd__or3b_2
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2487_ _4461_/Q _4469_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4226_ _4256_/A1 _2848_/B _4225_/Y _4081_/A vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__o211a_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4157_ _4224_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _4376_/Q _4680_/Q _3108_/S vssd1 vssd1 vccd1 vccd1 _3108_/X sky130_fd_sc_hd__mux2_1
X_4088_ _4092_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4089_/B sky130_fd_sc_hd__or2_1
XFILLER_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3039_ _3119_/A _3725_/B _3739_/A vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__and3b_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 rst vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2410_ _4548_/Q _4492_/Q _4484_/Q _4476_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2410_/X sky130_fd_sc_hd__mux4_1
X_3390_ _3634_/B _3390_/B vssd1 vssd1 vccd1 vccd1 _3396_/B sky130_fd_sc_hd__nand2_2
X_2341_ _2424_/A _2341_/B vssd1 vssd1 vccd1 vccd1 _2837_/A sky130_fd_sc_hd__or2_4
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2272_ _2300_/C _3629_/B _2300_/B vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__and3b_2
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _4011_/A _4011_/B _4019_/S _4011_/D vssd1 vssd1 vccd1 vccd1 _4011_/Y sky130_fd_sc_hd__nand4_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3726_ _3742_/A _3072_/B _3725_/Y vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__o21ai_1
X_3657_ _3754_/A1 _3655_/Y _3656_/X _3654_/X vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__o211a_1
X_3588_ _2351_/B _2288_/Y _2351_/C vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__o21ba_1
X_2608_ _4671_/Q _2607_/Y _2837_/A vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2539_ _2938_/A1 _2534_/X _2538_/X _2529_/X _2530_/X vssd1 vssd1 vccd1 vccd1 _2617_/C
+ sky130_fd_sc_hd__o32ai_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4209_ _3977_/X _4228_/B _4198_/Y _4208_/X vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout180 _3877_/Y vssd1 vssd1 vccd1 vccd1 _3899_/C sky130_fd_sc_hd__clkbuf_2
Xfanout191 _2310_/X vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__buf_6
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ _4356_/Q _4580_/Q _2892_/S vssd1 vssd1 vccd1 vccd1 _2891_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4582_/CLK _4560_/D vssd1 vssd1 vccd1 vccd1 _4560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3511_ _4525_/Q _4312_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4525_/D sky130_fd_sc_hd__mux2_1
X_4491_ _4684_/CLK _4491_/D vssd1 vssd1 vccd1 vccd1 _4491_/Q sky130_fd_sc_hd__dfxtp_2
X_3442_ _4464_/Q _3541_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4464_/D sky130_fd_sc_hd__mux2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _4427_/Q _3571_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4427_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2324_ _2284_/X _2285_/Y _2335_/C _2322_/Y vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__a211o_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _4641_/Q _4215_/A _4104_/A _4639_/Q vssd1 vssd1 vccd1 vccd1 _2263_/B sky130_fd_sc_hd__a22o_1
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2186_ _4599_/Q vssd1 vssd1 vccd1 vccd1 _2186_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4689_ _4689_/CLK _4689_/D vssd1 vssd1 vccd1 vccd1 _4689_/Q sky130_fd_sc_hd__dfxtp_2
X_3709_ _2901_/B _3708_/X _3771_/S vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3991_ _4238_/A _3991_/B vssd1 vssd1 vccd1 vccd1 _3991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2942_ _2942_/A _2994_/A vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__or2_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _4684_/Q _2932_/S _2872_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__a211o_1
X_4612_ _4629_/CLK _4612_/D vssd1 vssd1 vccd1 vccd1 _4612_/Q sky130_fd_sc_hd__dfxtp_1
X_4543_ _4543_/CLK _4543_/D vssd1 vssd1 vccd1 vccd1 _4543_/Q sky130_fd_sc_hd__dfxtp_1
X_4474_ _4553_/CLK _4474_/D vssd1 vssd1 vccd1 vccd1 _4474_/Q sky130_fd_sc_hd__dfxtp_1
X_3425_ _4449_/Q _3569_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4449_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3356_ _3572_/A _4330_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _3364_/S sky130_fd_sc_hd__and3_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2307_ _3633_/B _2307_/B _2307_/C _2307_/D vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__and4b_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3287_/A _3287_/B _3287_/C _3287_/D vssd1 vssd1 vccd1 vccd1 _3288_/C sky130_fd_sc_hd__and4_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2238_ _3846_/A _3930_/A _3931_/A _2373_/C vssd1 vssd1 vccd1 vccd1 _2295_/B sky130_fd_sc_hd__a2bb2o_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4190_ _4248_/A _4205_/A _4212_/B _3585_/Y vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3210_ _3210_/A _3283_/A vssd1 vssd1 vccd1 vccd1 _3211_/B sky130_fd_sc_hd__xnor2_1
X_3141_ _3086_/A _3140_/X _3139_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3141_/X sky130_fd_sc_hd__o211a_1
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3072_ _3072_/A _3072_/B _3068_/B vssd1 vssd1 vccd1 vccd1 _3209_/B sky130_fd_sc_hd__or3b_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3974_ _4112_/A _4112_/B vssd1 vssd1 vccd1 vccd1 _3974_/Y sky130_fd_sc_hd__nand2_2
X_2925_ _4501_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2925_/X sky130_fd_sc_hd__and3_1
X_2856_ _2917_/B _2855_/Y _2853_/X vssd1 vssd1 vccd1 vccd1 _2856_/Y sky130_fd_sc_hd__a21oi_4
X_2787_ _2337_/C _2780_/Y _2786_/X _2422_/A vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__a211o_1
X_4526_ _4582_/CLK _4526_/D vssd1 vssd1 vccd1 vccd1 _4526_/Q sky130_fd_sc_hd__dfxtp_1
X_4457_ _4555_/CLK _4457_/D vssd1 vssd1 vccd1 vccd1 _4457_/Q sky130_fd_sc_hd__dfxtp_1
X_3408_ _4071_/A2 _3390_/B _4011_/B _3405_/A vssd1 vssd1 vccd1 vccd1 _3408_/X sky130_fd_sc_hd__o2bb2a_2
X_4388_ _4584_/CLK _4388_/D vssd1 vssd1 vccd1 vccd1 _4388_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3339_ _4396_/Q _4331_/A1 _3346_/S vssd1 vssd1 vccd1 vccd1 _4396_/D sky130_fd_sc_hd__mux2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _2766_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__nand2_1
X_3690_ _3727_/S _3690_/B vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__nor2_1
X_2641_ _2639_/X _2640_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2572_ _2565_/Y _2568_/X _2571_/X vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4311_ _4676_/Q _4320_/A1 _4318_/S vssd1 vssd1 vccd1 vccd1 _4676_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4242_ _4226_/X _4240_/Y _4241_/Y vssd1 vssd1 vccd1 vccd1 _4242_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _4204_/B _3910_/X _3911_/Y _3922_/X vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__a211o_1
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3124_ _3760_/A _3124_/B vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3055_ _3252_/S _3055_/B vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__or2_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ _3959_/A _4188_/B vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _2913_/B _3231_/S _2907_/X vssd1 vssd1 vccd1 vccd1 _2908_/Y sky130_fd_sc_hd__a21oi_1
X_3888_ _4188_/B _4188_/C _4205_/A vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__o21ai_2
X_2839_ _2834_/A _3680_/B _3689_/B _3699_/B vssd1 vssd1 vccd1 vccd1 _2840_/B sky130_fd_sc_hd__a31o_1
X_4509_ _4544_/CLK _4509_/D vssd1 vssd1 vccd1 vccd1 _4509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_38_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4682_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4630_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3811_ _2360_/B _4241_/A _3812_/S vssd1 vssd1 vccd1 vccd1 _4621_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3742_ _3742_/A _3742_/B vssd1 vssd1 vccd1 vccd1 _3742_/Y sky130_fd_sc_hd__nand2_1
X_3673_ _3716_/A _2885_/B _3670_/Y vssd1 vssd1 vccd1 vccd1 _3673_/Y sky130_fd_sc_hd__o21ai_1
X_2624_ _2847_/A1 _2615_/X _2623_/X _2746_/A1 vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2555_ _3653_/B _2554_/Y _2555_/S vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__mux2_2
X_2486_ _2644_/S _2483_/X _2485_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__o211a_1
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4225_ _4223_/X _4224_/Y _4256_/A1 vssd1 vssd1 vccd1 vccd1 _4225_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4156_ _3936_/A _4155_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4659_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3107_ _3108_/S _4584_/Q _3113_/S1 vssd1 vssd1 vccd1 vccd1 _3107_/X sky130_fd_sc_hd__a21bo_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4087_ _4092_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4116_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3038_ _2961_/A _3273_/A _3739_/A vssd1 vssd1 vccd1 vccd1 _3040_/A sky130_fd_sc_hd__o21ba_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2424_/A _2341_/B vssd1 vssd1 vccd1 vccd1 _2348_/B sky130_fd_sc_hd__nor2_4
X_2271_ _2293_/A _4003_/A vssd1 vssd1 vccd1 vccd1 _2300_/C sky130_fd_sc_hd__or2_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4010_ _4010_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4011_/D sky130_fd_sc_hd__nand2_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3725_ _3742_/A _3725_/B vssd1 vssd1 vccd1 vccd1 _3725_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4490_/CLK sky130_fd_sc_hd__clkbuf_16
X_3656_ _3727_/S _3655_/Y _3653_/Y _3720_/S vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__a211o_1
X_3587_ _3587_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _3630_/C sky130_fd_sc_hd__nor2_1
X_2607_ _2607_/A _2669_/C vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2538_ _2814_/A1 _2535_/X _2537_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__o211a_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4208_ _4235_/A _4233_/B _4200_/Y _4207_/X vssd1 vssd1 vccd1 vccd1 _4208_/X sky130_fd_sc_hd__a31o_1
X_2469_ _2197_/Y _2746_/A1 _2427_/X _2468_/X vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__a211o_2
XFILLER_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _3872_/Y _4140_/B _3962_/Y vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout181 _3964_/A vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__buf_6
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout192 _4270_/B vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__buf_6
Xfanout170 _4123_/A vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__buf_4
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ _4524_/Q _4320_/A1 _3517_/S vssd1 vssd1 vccd1 vccd1 _4524_/D sky130_fd_sc_hd__mux2_1
X_4490_ _4490_/CLK _4490_/D vssd1 vssd1 vccd1 vccd1 _4490_/Q sky130_fd_sc_hd__dfxtp_1
X_3441_ _4463_/Q _3540_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4463_/D sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _4426_/Q _3570_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4426_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2323_ _2284_/X _2285_/Y _2335_/C _2322_/Y vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _3993_/A _4086_/A vssd1 vssd1 vccd1 vccd1 _4104_/A sky130_fd_sc_hd__nor2_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2185_ _4623_/Q vssd1 vssd1 vccd1 vccd1 _2185_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4688_ _4697_/CLK _4688_/D vssd1 vssd1 vccd1 vccd1 _4688_/Q sky130_fd_sc_hd__dfxtp_2
X_3708_ _2996_/A _2901_/B _3742_/A vssd1 vssd1 vccd1 vccd1 _3708_/X sky130_fd_sc_hd__mux2_1
X_3639_ _4061_/B _3747_/B2 _3666_/B1 _3638_/X vssd1 vssd1 vccd1 vccd1 _3640_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _3990_/A _3990_/B _3990_/C _3990_/D vssd1 vssd1 vccd1 vccd1 _3990_/X sky130_fd_sc_hd__or4_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2941_ _3209_/A _3072_/A vssd1 vssd1 vccd1 vccd1 _2994_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611_ _4629_/CLK _4611_/D vssd1 vssd1 vccd1 vccd1 _4611_/Q sky130_fd_sc_hd__dfxtp_1
X_2872_ _4412_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__and3_1
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4542_ _4574_/CLK _4542_/D vssd1 vssd1 vccd1 vccd1 _4542_/Q sky130_fd_sc_hd__dfxtp_1
X_4473_ _4481_/CLK _4473_/D vssd1 vssd1 vccd1 vccd1 _4473_/Q sky130_fd_sc_hd__dfxtp_1
X_3424_ _4448_/Q _3568_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4448_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3355_ _4411_/Q _3580_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4411_/D sky130_fd_sc_hd__mux2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2306_ _2306_/A _2425_/A _3987_/B _2306_/D vssd1 vssd1 vccd1 vccd1 _2307_/B sky130_fd_sc_hd__and4_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3283_/A _3286_/B vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__and2b_1
X_2237_ _2373_/B _3846_/A vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__nand2b_4
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _4569_/Q _4529_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3071_ _3209_/A _3072_/A _3072_/B _3067_/Y vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__o31ai_2
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3973_ _3973_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _4112_/B sky130_fd_sc_hd__and2_1
X_2924_ _2937_/A1 _2923_/X _2922_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2855_ _4491_/Q _2854_/B _2389_/A vssd1 vssd1 vccd1 vccd1 _2855_/Y sky130_fd_sc_hd__a21oi_2
X_4525_ _4581_/CLK _4525_/D vssd1 vssd1 vccd1 vccd1 _4525_/Q sky130_fd_sc_hd__dfxtp_1
X_2786_ _3041_/A _2783_/Y _2785_/X _2844_/A vssd1 vssd1 vccd1 vccd1 _2786_/X sky130_fd_sc_hd__o211a_1
X_4456_ _4552_/CLK _4456_/D vssd1 vssd1 vccd1 vccd1 _4456_/Q sky130_fd_sc_hd__dfxtp_1
X_3407_ _4057_/A _3407_/B vssd1 vssd1 vccd1 vccd1 _4011_/B sky130_fd_sc_hd__nand2_1
X_4387_ _4587_/CLK _4387_/D vssd1 vssd1 vccd1 vccd1 _4387_/Q sky130_fd_sc_hd__dfxtp_1
X_3338_ _3572_/A _4330_/A _3446_/C vssd1 vssd1 vccd1 vccd1 _3346_/S sky130_fd_sc_hd__and3_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3267_/X _3268_/X _3269_/S vssd1 vssd1 vccd1 vccd1 _3270_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2640_ _4496_/Q _4552_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__mux2_1
X_2571_ _2571_/A _2571_/B _2570_/X vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__or3b_1
X_4310_ _4310_/A _4310_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _4318_/S sky130_fd_sc_hd__and3_4
X_4241_ _4241_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4241_/Y sky130_fd_sc_hd__nand2_1
X_4172_ _4172_/A _4228_/B _4172_/C vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__and3_1
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3123_ _3232_/S _3121_/X _3122_/X vssd1 vssd1 vccd1 vccd1 _3126_/B sky130_fd_sc_hd__a21o_1
X_3054_ _4503_/Q _4559_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3055_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _3956_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4233_/A sky130_fd_sc_hd__and2_2
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2907_ _2907_/A _2907_/B _2959_/B vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__or3_1
X_3887_ _4161_/A _3886_/X _3870_/Y vssd1 vssd1 vccd1 vccd1 _4188_/C sky130_fd_sc_hd__o21ai_2
X_2838_ _3857_/B _2837_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__o21a_1
X_2769_ _4578_/Q _4522_/Q _4514_/Q _4354_/Q _2950_/S _2404_/A vssd1 vssd1 vccd1 vccd1
+ _2769_/X sky130_fd_sc_hd__mux4_2
X_4508_ _4576_/CLK _4508_/D vssd1 vssd1 vccd1 vccd1 _4508_/Q sky130_fd_sc_hd__dfxtp_1
X_4439_ _4692_/CLK _4439_/D vssd1 vssd1 vccd1 vccd1 _4439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3810_ _3623_/B input9/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4620_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3741_ _3740_/X _4602_/Q _3741_/S vssd1 vssd1 vccd1 vccd1 _4602_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3672_ _4488_/Q _3762_/B _4013_/S vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__or3_1
X_2623_ _3290_/A _2595_/Y _2622_/X _2382_/X vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__o211a_1
X_2554_ _3643_/B _3652_/B vssd1 vssd1 vccd1 vccd1 _2554_/Y sky130_fd_sc_hd__xnor2_1
X_2485_ _4485_/Q _2699_/S _2484_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__a211o_1
X_4224_ _4224_/A _4224_/B vssd1 vssd1 vccd1 vccd1 _4224_/Y sky130_fd_sc_hd__nor2_1
X_4155_ _4240_/A _4153_/Y _4154_/Y _4270_/B input7/X vssd1 vssd1 vccd1 vccd1 _4155_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3106_ _3108_/S _4360_/Q vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4086_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4266_/B sky130_fd_sc_hd__or2_2
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3037_ _3031_/X _3033_/X _3036_/X _3270_/A vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__o22a_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _3941_/A _4063_/A vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__nand2_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2270_ _4042_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _2300_/B sky130_fd_sc_hd__and2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3724_ _4600_/Q _3741_/S _3723_/Y vssd1 vssd1 vccd1 vccd1 _4600_/D sky130_fd_sc_hd__a21o_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3655_ _3716_/A _2617_/C _3652_/Y vssd1 vssd1 vccd1 vccd1 _3655_/Y sky130_fd_sc_hd__o21ai_1
X_2606_ _3643_/B _3652_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__and3_1
X_3586_ _3930_/A _3585_/Y _3401_/Y vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__o21ai_2
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2537_ _4454_/Q _2699_/S _2536_/X _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__a211o_1
X_2468_ _3185_/A _2377_/Y _2467_/X _2466_/X _2363_/B vssd1 vssd1 vccd1 vccd1 _2468_/X
+ sky130_fd_sc_hd__o32a_1
X_4207_ _3924_/X _4260_/B _4204_/Y _4206_/X vssd1 vssd1 vccd1 vccd1 _4207_/X sky130_fd_sc_hd__a31o_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2399_ _2859_/A _3318_/B vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__nor2_4
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4224_/A _3068_/B _4137_/X vssd1 vssd1 vccd1 vccd1 _4138_/Y sky130_fd_sc_hd__o21ai_2
X_4069_ _3941_/A _4272_/S _4067_/X _4068_/X vssd1 vssd1 vccd1 vccd1 _4656_/D sky130_fd_sc_hd__o22a_1
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout182 _3959_/A vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__buf_4
Xfanout160 _3385_/Y vssd1 vssd1 vccd1 vccd1 _3713_/A sky130_fd_sc_hd__buf_4
Xfanout171 _4123_/A vssd1 vssd1 vccd1 vccd1 _3407_/B sky130_fd_sc_hd__buf_4
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout193 _4270_/B vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__buf_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _4462_/Q _3539_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4462_/D sky130_fd_sc_hd__mux2_1
X_3371_ _4425_/Q _3569_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4425_/D sky130_fd_sc_hd__mux2_1
X_2322_ _3581_/C _2384_/D vssd1 vssd1 vccd1 vccd1 _2322_/Y sky130_fd_sc_hd__nand2_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2366_/B _2384_/B vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__nand2_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2184_ _4604_/Q vssd1 vssd1 vccd1 vccd1 _2184_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4687_ _4698_/CLK _4687_/D vssd1 vssd1 vccd1 vccd1 _4687_/Q sky130_fd_sc_hd__dfxtp_2
X_3707_ _4598_/Q _3741_/S _3706_/X vssd1 vssd1 vccd1 vccd1 _4598_/D sky130_fd_sc_hd__a21bo_1
X_3638_ _4484_/Q _3987_/A _4013_/S _3637_/X vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__o31a_1
X_3569_ _4577_/Q _3569_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4577_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2940_ _2940_/A _2995_/A vssd1 vssd1 vccd1 vccd1 _3072_/A sky130_fd_sc_hd__or2_2
X_2871_ _2937_/C1 _2868_/X _2870_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__a31o_2
X_4610_ _4629_/CLK _4610_/D vssd1 vssd1 vccd1 vccd1 _4610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4541_ _4544_/CLK _4541_/D vssd1 vssd1 vccd1 vccd1 _4541_/Q sky130_fd_sc_hd__dfxtp_1
X_4472_ _4651_/CLK _4472_/D vssd1 vssd1 vccd1 vccd1 _4472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3423_ _4447_/Q _3567_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4447_/D sky130_fd_sc_hd__mux2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _4410_/Q _4317_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4410_/D sky130_fd_sc_hd__mux2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _3771_/S _3581_/D _2288_/Y _2301_/X _2217_/B vssd1 vssd1 vccd1 vccd1 _2306_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3287_/A _3287_/B _3287_/C _4224_/B _3286_/B vssd1 vssd1 vccd1 vccd1 _3288_/B
+ sky130_fd_sc_hd__a41oi_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2373_/B _3846_/A vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__and2b_2
XFILLER_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ _2996_/X _3068_/B _3105_/A vssd1 vssd1 vccd1 vccd1 _3070_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _3972_/A _4116_/A vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2923_ _4677_/Q _4373_/Q _2934_/S vssd1 vssd1 vccd1 vccd1 _2923_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2854_ _4491_/Q _2854_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__or2_2
X_2785_ _2612_/S _2784_/X _2782_/X _2904_/A vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__a211o_1
X_4524_ _4695_/CLK _4524_/D vssd1 vssd1 vccd1 vccd1 _4524_/Q sky130_fd_sc_hd__dfxtp_1
X_4455_ _4667_/CLK _4455_/D vssd1 vssd1 vccd1 vccd1 _4455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3406_ _4664_/Q _3417_/S _3405_/X _4037_/A vssd1 vssd1 vccd1 vccd1 _4440_/D sky130_fd_sc_hd__o211a_1
X_4386_ _4587_/CLK _4386_/D vssd1 vssd1 vccd1 vccd1 _4386_/Q sky130_fd_sc_hd__dfxtp_1
X_3337_ _4395_/Q _3580_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4395_/D sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _4371_/Q _4700_/Q _4691_/Q _4419_/Q _4440_/Q _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3268_/X sky130_fd_sc_hd__mux4_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2219_ _4590_/Q _3618_/A _4588_/Q _3836_/A vssd1 vssd1 vccd1 vccd1 _2424_/A sky130_fd_sc_hd__or4_4
X_3199_ _3065_/S _3196_/X _3198_/X _3249_/C1 vssd1 vssd1 vccd1 vccd1 _3199_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _4484_/Q _4485_/Q _4486_/Q vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__or3_1
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4240_ _4240_/A _4240_/B vssd1 vssd1 vccd1 vccd1 _4240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4171_ _3870_/Y _3961_/A _3962_/Y _3975_/Y vssd1 vssd1 vccd1 vccd1 _4172_/C sky130_fd_sc_hd__a211o_1
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3122_ _4672_/Q _2907_/A _3020_/S vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ _3051_/X _3052_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _3956_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__or2_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2906_ _3013_/B _2906_/B vssd1 vssd1 vccd1 vccd1 _2959_/B sky130_fd_sc_hd__nor2_1
X_3886_ _3964_/B _4104_/B _3964_/A vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__a21o_1
X_2837_ _2837_/A _2844_/B vssd1 vssd1 vccd1 vccd1 _2837_/Y sky130_fd_sc_hd__nand2_1
X_2768_ _4662_/Q _2712_/B _2768_/B1 _2767_/Y vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__o211a_1
X_4507_ _4683_/CLK _4507_/D vssd1 vssd1 vccd1 vccd1 _4507_/Q sky130_fd_sc_hd__dfxtp_1
X_2699_ _4497_/Q _4553_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__mux2_1
X_4438_ _4629_/CLK _4438_/D vssd1 vssd1 vccd1 vccd1 _4438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4369_ _4698_/CLK _4369_/D vssd1 vssd1 vccd1 vccd1 _4369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _2432_/X _3068_/B _3713_/A _3738_/X _3739_/X vssd1 vssd1 vccd1 vccd1 _3740_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3727_/S _3671_/B vssd1 vssd1 vccd1 vccd1 _3671_/Y sky130_fd_sc_hd__nor2_1
X_2622_ _3185_/A _2622_/B vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__or2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2553_ _2668_/A1 _2543_/Y _2547_/Y _2549_/Y _2551_/Y vssd1 vssd1 vccd1 vccd1 _3653_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2484_ _4477_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2484_/X sky130_fd_sc_hd__and3_1
X_4223_ _4662_/Q _3933_/B _4057_/X _4222_/X _4224_/A vssd1 vssd1 vccd1 vccd1 _4223_/X
+ sky130_fd_sc_hd__o311a_1
X_4154_ _4150_/X _4152_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _4154_/Y sky130_fd_sc_hd__o21ai_1
X_4085_ _4086_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4235_/A sky130_fd_sc_hd__nor2_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3105_ _3105_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _3105_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3036_ _3034_/X _3035_/X _3036_/S vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3938_/Y sky130_fd_sc_hd__nand2_2
X_3869_ _3936_/A _4671_/Q vssd1 vssd1 vccd1 vccd1 _3960_/B sky130_fd_sc_hd__and2b_4
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3723_ _3739_/B _3721_/X _3722_/X vssd1 vssd1 vccd1 vccd1 _3723_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3654_ _4486_/Q _3762_/B _3691_/C vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__or3_1
X_2605_ _2599_/X _2601_/X _2604_/X _2668_/A1 vssd1 vssd1 vccd1 vccd1 _2669_/C sky130_fd_sc_hd__o22a_4
X_3585_ _3993_/A _3585_/B vssd1 vssd1 vccd1 vccd1 _3585_/Y sky130_fd_sc_hd__nand2_4
X_2536_ _4446_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__and3_1
X_2467_ _3966_/B _2712_/B _2768_/B1 vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__o21a_1
X_4206_ _2225_/Y _3947_/X _4205_/Y _4203_/X vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2398_ _4646_/Q _2385_/Y _2396_/X vssd1 vssd1 vccd1 vccd1 _3318_/B sky130_fd_sc_hd__o21ai_4
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4059_/A _4136_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__o21a_1
X_4068_ input1/X _4270_/B _4272_/S vssd1 vssd1 vccd1 vccd1 _4068_/X sky130_fd_sc_hd__a21bo_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3019_ _3725_/B _3023_/B _3742_/A vssd1 vssd1 vccd1 vccd1 _3019_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout172 _4238_/A vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__buf_4
Xfanout150 _2758_/B vssd1 vssd1 vccd1 vccd1 _2812_/B sky130_fd_sc_hd__buf_4
Xfanout161 _3384_/Y vssd1 vssd1 vccd1 vccd1 _3739_/B sky130_fd_sc_hd__buf_8
Xfanout183 _2431_/Y vssd1 vssd1 vccd1 vccd1 _3731_/A1 sky130_fd_sc_hd__buf_6
Xfanout194 _2205_/X vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__buf_6
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3370_ _4424_/Q _3568_/A1 _3373_/S vssd1 vssd1 vccd1 vccd1 _4424_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2321_ _3384_/A _2424_/A vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__or2_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _3993_/A _4091_/A vssd1 vssd1 vccd1 vccd1 _4215_/A sky130_fd_sc_hd__nor2_4
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _4628_/Q vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3731_/A1 _2848_/C _3739_/B _3704_/X _3705_/Y vssd1 vssd1 vccd1 vccd1 _3706_/X
+ sky130_fd_sc_hd__a221o_4
X_4686_ _4697_/CLK _4686_/D vssd1 vssd1 vccd1 vccd1 _4686_/Q sky130_fd_sc_hd__dfxtp_2
X_3637_ _3754_/A1 _3635_/Y _3636_/X _4010_/A vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__o22a_1
X_3568_ _4576_/Q _3568_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4576_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2519_ _4484_/Q _4485_/Q vssd1 vssd1 vccd1 vccd1 _2519_/Y sky130_fd_sc_hd__xnor2_1
X_3499_ _4515_/Q _3571_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4515_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _4524_/Q _2934_/S _2869_/X _2937_/A1 vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_10_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4551_/CLK sky130_fd_sc_hd__clkbuf_16
X_4540_ _4576_/CLK _4540_/D vssd1 vssd1 vccd1 vccd1 _4540_/Q sky130_fd_sc_hd__dfxtp_1
X_4471_ _4667_/CLK _4471_/D vssd1 vssd1 vccd1 vccd1 _4471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3422_ _4446_/Q _3539_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4446_/D sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _4409_/Q _4316_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4409_/D sky130_fd_sc_hd__mux2_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2304_ _4439_/Q _3581_/C vssd1 vssd1 vccd1 vccd1 _2307_/C sky130_fd_sc_hd__nand2_1
X_3284_ _3210_/A _3283_/Y _3258_/Y _3209_/X vssd1 vssd1 vccd1 vccd1 _3290_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2235_ _2349_/B _2233_/Y _2234_/X _3989_/A vssd1 vssd1 vccd1 vccd1 _4438_/D sky130_fd_sc_hd__a22o_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2999_ _3288_/A _2994_/Y _2998_/Y _2860_/C vssd1 vssd1 vccd1 vccd1 _2999_/X sky130_fd_sc_hd__a211o_1
X_4669_ _4671_/CLK _4669_/D vssd1 vssd1 vccd1 vccd1 _4669_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ _3972_/A _4119_/B _4083_/A vssd1 vssd1 vccd1 vccd1 _4112_/A sky130_fd_sc_hd__a21o_1
X_2922_ _4357_/Q _2934_/S _2921_/X _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2922_/X sky130_fd_sc_hd__a211o_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2853_ _2820_/X _2821_/Y _2852_/X vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__o21a_2
X_2784_ _3689_/B _2783_/Y _2841_/S vssd1 vssd1 vccd1 vccd1 _2784_/X sky130_fd_sc_hd__mux2_1
X_4523_ _4579_/CLK _4523_/D vssd1 vssd1 vccd1 vccd1 _4523_/Q sky130_fd_sc_hd__dfxtp_1
X_4454_ _4481_/CLK _4454_/D vssd1 vssd1 vccd1 vccd1 _4454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3405_ _3405_/A _3405_/B _3417_/S vssd1 vssd1 vccd1 vccd1 _3405_/X sky130_fd_sc_hd__or3b_1
X_4385_ _4698_/CLK _4385_/D vssd1 vssd1 vccd1 vccd1 _4385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3336_ _4394_/Q _4337_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4394_/D sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3267_ _4387_/Q _4395_/Q _4411_/Q _4403_/Q _3264_/S _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3267_/X sky130_fd_sc_hd__mux4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2218_ _3826_/A _3989_/A vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__nor2_8
X_3198_ _3255_/S _3198_/B vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__or2_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4080_/S _2708_/B _4169_/Y _3407_/B vssd1 vssd1 vccd1 vccd1 _4170_/Y sky130_fd_sc_hd__o211ai_4
X_3121_ _3174_/A _3124_/B _3175_/A _3116_/X vssd1 vssd1 vccd1 vccd1 _3121_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3052_ _4583_/Q _4359_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3052_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3954_ _3956_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _3954_/Y sky130_fd_sc_hd__nor2_1
X_3885_ _4104_/B vssd1 vssd1 vccd1 vccd1 _3885_/Y sky130_fd_sc_hd__inv_2
X_2905_ _3013_/B _3174_/A _2906_/B vssd1 vssd1 vccd1 vccd1 _2907_/B sky130_fd_sc_hd__and3_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2836_ _2961_/A _3013_/A _2832_/X vssd1 vssd1 vccd1 vccd1 _2844_/B sky130_fd_sc_hd__o21ai_1
X_2767_ _2472_/Y _2766_/Y _2618_/B vssd1 vssd1 vccd1 vccd1 _2767_/Y sky130_fd_sc_hd__o21ai_1
X_2698_ _2937_/C1 _2691_/X _2693_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__a31o_2
X_4506_ _4570_/CLK _4506_/D vssd1 vssd1 vccd1 vccd1 _4506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4437_ _4613_/CLK _4437_/D vssd1 vssd1 vccd1 vccd1 _4437_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4697_/CLK _4368_/D vssd1 vssd1 vccd1 vccd1 _4368_/Q sky130_fd_sc_hd__dfxtp_1
X_4299_ _4661_/Q _4278_/Y _4298_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__a22o_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _4310_/B _3563_/C _3446_/C vssd1 vssd1 vccd1 vccd1 _3327_/S sky130_fd_sc_hd__and3_4
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ _3716_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__nand2_1
X_2621_ _2363_/B _2620_/X _2768_/B1 vssd1 vssd1 vccd1 vccd1 _2621_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2552_ _2668_/A1 _2543_/Y _2547_/Y _2549_/Y _2551_/Y vssd1 vssd1 vccd1 vccd1 _3652_/B
+ sky130_fd_sc_hd__a32oi_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4222_ _4104_/A _4216_/X _4217_/Y _4221_/X vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__a31o_1
X_2483_ _4493_/Q _4549_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__mux2_1
X_4153_ _4080_/S _2617_/D _4138_/Y _3407_/B vssd1 vssd1 vccd1 vccd1 _4153_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4084_ _4084_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4095_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3104_ _3935_/A _3259_/B _3160_/B1 vssd1 vssd1 vccd1 vccd1 _3104_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3035_ _4367_/Q _4696_/Q _4687_/Q _4415_/Q _3264_/S _3265_/A vssd1 vssd1 vccd1 vccd1
+ _3035_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3937_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _4127_/B sky130_fd_sc_hd__and2_1
X_3868_ _4188_/B _3907_/B vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__or2_4
X_3799_ _4606_/Q _4598_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__mux2_1
X_2819_ _2766_/A _2817_/D _2818_/X vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3722_ _3731_/A1 _2995_/A _3013_/C _3640_/A _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3722_/X
+ sky130_fd_sc_hd__a221o_1
X_3653_ _3727_/S _3653_/B vssd1 vssd1 vccd1 vccd1 _3653_/Y sky130_fd_sc_hd__nor2_1
X_2604_ _2602_/X _2603_/X _2889_/A vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_2
X_3584_ _4056_/B _3931_/A vssd1 vssd1 vccd1 vccd1 _3584_/Y sky130_fd_sc_hd__nor2_2
X_2535_ _4462_/Q _4470_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2466_ _2938_/A1 _2460_/Y _2465_/Y _2455_/Y _2448_/Y vssd1 vssd1 vccd1 vccd1 _2466_/X
+ sky130_fd_sc_hd__o32a_4
X_4205_ _4205_/A _4205_/B _4205_/C vssd1 vssd1 vccd1 vccd1 _4205_/Y sky130_fd_sc_hd__nand3_1
X_4136_ _3936_/A _4671_/Q _4057_/X _4128_/X _4135_/X vssd1 vssd1 vccd1 vccd1 _4136_/X
+ sky130_fd_sc_hd__o32a_1
X_2397_ _4646_/Q _2385_/Y _2396_/X vssd1 vssd1 vccd1 vccd1 _3299_/B sky130_fd_sc_hd__o21a_2
XFILLER_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4010_/A _4060_/X _4061_/Y _4240_/A _4066_/X vssd1 vssd1 vccd1 vccd1 _4067_/X
+ sky130_fd_sc_hd__o311a_1
X_3018_ _3938_/B _3017_/X _3232_/S vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout140 _2927_/C vssd1 vssd1 vccd1 vccd1 _2798_/C sky130_fd_sc_hd__clkbuf_2
Xfanout173 _2242_/X vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__buf_6
Xfanout151 _2863_/B vssd1 vssd1 vccd1 vccd1 _2758_/B sky130_fd_sc_hd__buf_4
Xfanout162 _3384_/Y vssd1 vssd1 vccd1 vccd1 _3749_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout195 _4300_/S vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__buf_6
Xfanout184 _2380_/A vssd1 vssd1 vccd1 vccd1 _2473_/C sky130_fd_sc_hd__buf_6
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2320_ _3384_/A _2424_/A vssd1 vssd1 vccd1 vccd1 _2384_/D sky130_fd_sc_hd__nor2_4
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2248_/Y _2250_/X _2366_/B vssd1 vssd1 vccd1 vccd1 _2263_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2182_ _4606_/Q vssd1 vssd1 vccd1 vccd1 _2182_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3705_ _3699_/B _3739_/B _3749_/C1 vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__o21bai_1
X_4685_ _4694_/CLK _4685_/D vssd1 vssd1 vccd1 vccd1 _4685_/Q sky130_fd_sc_hd__dfxtp_2
X_3636_ _3275_/S _3635_/Y _3727_/S vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__mux2_1
X_3567_ _4575_/Q _3567_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4575_/D sky130_fd_sc_hd__mux2_1
X_2518_ _2768_/B1 _2496_/X _2517_/X _2746_/A1 vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__a211o_1
X_3498_ _4514_/Q _3570_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4514_/D sky130_fd_sc_hd__mux2_1
X_2449_ _2798_/B _2798_/C _4428_/Q vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4119_ _4119_/A _4119_/B vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4481_/CLK _4470_/D vssd1 vssd1 vccd1 vccd1 _4470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3421_ _4445_/Q _3565_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4445_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3352_ _4408_/Q _4335_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4408_/D sky130_fd_sc_hd__mux2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _4620_/Q _3387_/B vssd1 vssd1 vccd1 vccd1 _3633_/B sky130_fd_sc_hd__nor2_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3283_/A _3286_/B vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__nand2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2234_ _4042_/A _2274_/A vssd1 vssd1 vccd1 vccd1 _2234_/X sky130_fd_sc_hd__and2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2998_ _2996_/X _2997_/X _3288_/A vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__a21oi_1
X_4668_ _4672_/CLK _4668_/D vssd1 vssd1 vccd1 vccd1 _4668_/Q sky130_fd_sc_hd__dfxtp_4
X_3619_ _3799_/S _3619_/B vssd1 vssd1 vccd1 vccd1 _3619_/X sky130_fd_sc_hd__or2_1
X_4599_ _4691_/CLK _4599_/D vssd1 vssd1 vccd1 vccd1 _4599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _4082_/A _4082_/B vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__and2_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2921_ _4581_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2921_/X sky130_fd_sc_hd__and3_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2852_ _2652_/A _2819_/Y _2851_/X _2655_/Y _2847_/Y vssd1 vssd1 vccd1 vccd1 _2852_/X
+ sky130_fd_sc_hd__o221a_1
X_2783_ _2783_/A _3689_/B vssd1 vssd1 vccd1 vccd1 _2783_/Y sky130_fd_sc_hd__xnor2_1
X_4522_ _4581_/CLK _4522_/D vssd1 vssd1 vccd1 vccd1 _4522_/Q sky130_fd_sc_hd__dfxtp_1
X_4453_ _4464_/CLK _4453_/D vssd1 vssd1 vccd1 vccd1 _4453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3404_ _2373_/B _4063_/A _4010_/A vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__mux2_1
X_4384_ _4683_/CLK _4384_/D vssd1 vssd1 vccd1 vccd1 _4384_/Q sky130_fd_sc_hd__dfxtp_1
X_3335_ _4393_/Q _4316_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4393_/D sky130_fd_sc_hd__mux2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3266_ _3266_/A1 _3263_/Y _3265_/Y _3261_/A vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__a211o_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _4062_/A _2217_/B vssd1 vssd1 vccd1 vccd1 _2217_/Y sky130_fd_sc_hd__nand2_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _4570_/Q _4530_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3198_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3040_/B _3742_/B _3173_/A vssd1 vssd1 vccd1 vccd1 _3124_/B sky130_fd_sc_hd__o21ai_1
X_3051_ _4679_/Q _4375_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _4266_/A _3953_/B vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__or2_1
X_3884_ _3881_/A _3883_/X _3899_/C vssd1 vssd1 vccd1 vccd1 _4104_/B sky130_fd_sc_hd__a21o_1
X_2904_ _2904_/A _2904_/B vssd1 vssd1 vccd1 vccd1 _2906_/B sky130_fd_sc_hd__nand2_1
X_2835_ _2961_/A _3013_/A vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__nor2_1
X_2766_ _2766_/A _2848_/B vssd1 vssd1 vccd1 vccd1 _2766_/Y sky130_fd_sc_hd__xnor2_1
X_2697_ _2805_/C1 _2694_/X _2696_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__o211a_2
X_4505_ _4584_/CLK _4505_/D vssd1 vssd1 vccd1 vccd1 _4505_/Q sky130_fd_sc_hd__dfxtp_1
X_4436_ _4702_/CLK _4436_/D vssd1 vssd1 vccd1 vccd1 _4436_/Q sky130_fd_sc_hd__dfxtp_1
X_4367_ _4696_/CLK _4367_/D vssd1 vssd1 vccd1 vccd1 _4367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3318_/A _3318_/B vssd1 vssd1 vccd1 vccd1 _3446_/C sky130_fd_sc_hd__nor2_4
X_4298_ _4645_/Q _2367_/Y _3629_/Y _4653_/Q vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__a22o_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3249_ _2443_/X _3244_/X _3246_/X _3248_/X _3249_/C1 vssd1 vssd1 vccd1 vccd1 _3249_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2620_ _2595_/Y _2622_/B _3288_/A vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__mux2_1
X_2551_ _2889_/A _2550_/X _2898_/A vssd1 vssd1 vccd1 vccd1 _2551_/Y sky130_fd_sc_hd__a21oi_4
X_2482_ _2937_/C1 _2479_/X _2481_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__a31o_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4221_ _4221_/A _4221_/B _4221_/C _4219_/X vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__or4b_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4152_ _3975_/Y _4151_/X _4228_/B vssd1 vssd1 vccd1 vccd1 _4152_/X sky130_fd_sc_hd__o21a_1
X_4083_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__or2_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3103_ _2655_/B _3102_/Y _3259_/B vssd1 vssd1 vccd1 vccd1 _3103_/X sky130_fd_sc_hd__o21a_1
X_3034_ _4383_/Q _4391_/Q _4407_/Q _4399_/Q _3216_/S _3266_/A1 vssd1 vssd1 vccd1 vccd1
+ _3034_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _3936_/A _4671_/Q vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__nand2_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3867_ _4188_/B _3907_/B vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__nor2_8
X_3798_ _3619_/B _3796_/X _3797_/X _2274_/A vssd1 vssd1 vccd1 vccd1 _4613_/D sky130_fd_sc_hd__o211a_1
X_2818_ _2766_/A _2848_/B _2848_/C vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__o21a_1
X_2749_ _4538_/Q _2927_/B _2927_/C vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__and3_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4419_ _4700_/CLK _4419_/D vssd1 vssd1 vccd1 vccd1 _4419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3721_ _3666_/B1 _3720_/X _2995_/A _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__a2bb2o_1
X_3652_ _3716_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3652_/Y sky130_fd_sc_hd__nand2_1
X_3583_ _3927_/A _4248_/A _2368_/B vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__o21ai_4
X_2603_ _4471_/Q _4463_/Q _4455_/Q _4447_/Q _2775_/S0 _2829_/S1 vssd1 vssd1 vccd1
+ vccd1 _2603_/X sky130_fd_sc_hd__mux4_1
X_2534_ _2814_/A1 _2531_/X _2533_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__o211a_1
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2465_ _2463_/X _2464_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2465_/Y sky130_fd_sc_hd__a21oi_1
X_4204_ _4204_/A _4204_/B _4204_/C vssd1 vssd1 vccd1 vccd1 _4204_/Y sky130_fd_sc_hd__nand3_1
X_2396_ _4666_/Q _2847_/A1 _2768_/B1 _4057_/B _2382_/X vssd1 vssd1 vccd1 vccd1 _2396_/X
+ sky130_fd_sc_hd__a221o_4
X_4135_ _4135_/A _4135_/B _4135_/C _4134_/X vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__or4b_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4066_ _4643_/Q _3931_/Y _4064_/Y _4065_/X vssd1 vssd1 vccd1 vccd1 _4066_/X sky130_fd_sc_hd__a211o_1
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3017_ _3231_/S _3023_/B _3176_/A _3016_/Y vssd1 vssd1 vccd1 vccd1 _3017_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _3972_/A _4082_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout130 _2369_/Y vssd1 vssd1 vccd1 vccd1 _3239_/A sky130_fd_sc_hd__buf_6
Xfanout152 _2863_/B vssd1 vssd1 vccd1 vccd1 _2990_/B sky130_fd_sc_hd__buf_4
Xfanout141 _2863_/C vssd1 vssd1 vccd1 vccd1 _2927_/C sky130_fd_sc_hd__buf_4
Xfanout174 _3773_/S vssd1 vssd1 vccd1 vccd1 _3720_/S sky130_fd_sc_hd__buf_6
Xfanout163 _2725_/X vssd1 vssd1 vccd1 vccd1 _3680_/B sky130_fd_sc_hd__buf_6
Xfanout196 _2204_/Y vssd1 vssd1 vccd1 vccd1 _4300_/S sky130_fd_sc_hd__buf_6
Xfanout185 _4256_/A1 vssd1 vssd1 vccd1 vccd1 _4080_/S sky130_fd_sc_hd__buf_6
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _3931_/A _2244_/X _2245_/X _4086_/A _2180_/Y vssd1 vssd1 vccd1 vccd1 _2250_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2181_ _4630_/Q vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3704_ _3666_/B1 _3703_/X _2848_/C _3747_/B2 vssd1 vssd1 vccd1 vccd1 _3704_/X sky130_fd_sc_hd__a2bb2o_1
X_4684_ _4684_/CLK _4684_/D vssd1 vssd1 vccd1 vccd1 _4684_/Q sky130_fd_sc_hd__dfxtp_4
X_3635_ _3927_/A _4061_/B _2511_/A vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__o21ai_1
X_3566_ _4574_/Q _3566_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4574_/D sky130_fd_sc_hd__mux2_1
X_2517_ _2385_/A _2385_/B _2517_/S vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__mux2_1
X_3497_ _4513_/Q _3569_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4513_/D sky130_fd_sc_hd__mux2_1
X_2448_ _2446_/X _2447_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2448_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2379_ _4238_/A _2277_/X _2378_/X _4050_/C _2306_/A vssd1 vssd1 vccd1 vccd1 _2380_/B
+ sky130_fd_sc_hd__o32a_4
X_4118_ _3921_/A _3921_/B _4260_/B vssd1 vssd1 vccd1 vccd1 _4118_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4049_ _3383_/B _4303_/B2 _3990_/B _2333_/B vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420_ _4444_/Q _3537_/A1 _3427_/S vssd1 vssd1 vccd1 vccd1 _4444_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3351_ _4407_/Q _4334_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4407_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2302_ _2302_/A _3991_/B vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__or2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A _3282_/B _3282_/C vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__nand3_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2233_ _4631_/Q _4011_/A _2233_/C vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__nor3_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ _3287_/A _2995_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__a21o_1
X_4667_ _4667_/CLK _4667_/D vssd1 vssd1 vccd1 vccd1 _4667_/Q sky130_fd_sc_hd__dfxtp_4
X_3618_ _3618_/A _3619_/B vssd1 vssd1 vccd1 vccd1 _3827_/S sky130_fd_sc_hd__nor2_8
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4598_ _4700_/CLK _4598_/D vssd1 vssd1 vccd1 vccd1 _4598_/Q sky130_fd_sc_hd__dfxtp_1
X_3549_ _4559_/Q _4314_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4559_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _4662_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2920_ _4356_/Q _4320_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4356_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _2886_/A _2851_/B vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__and2b_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2782_ _2348_/B _2780_/Y _2781_/X _3276_/B vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__o211a_1
X_4521_ _4545_/CLK _4521_/D vssd1 vssd1 vccd1 vccd1 _4521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4452_ _4555_/CLK _4452_/D vssd1 vssd1 vccd1 vccd1 _4452_/Q sky130_fd_sc_hd__dfxtp_1
X_3403_ _4003_/B _2190_/Y _4003_/A _3397_/Y _3834_/B vssd1 vssd1 vccd1 vccd1 _3417_/S
+ sky130_fd_sc_hd__o311a_4
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4383_ _4679_/CLK _4383_/D vssd1 vssd1 vccd1 vccd1 _4383_/Q sky130_fd_sc_hd__dfxtp_1
X_3334_ _4392_/Q _3577_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4392_/D sky130_fd_sc_hd__mux2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3265_ _3265_/A _3265_/B vssd1 vssd1 vccd1 vccd1 _3265_/Y sky130_fd_sc_hd__nor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _3623_/B _4619_/Q _3623_/C _3622_/B vssd1 vssd1 vccd1 vccd1 _2217_/B sky130_fd_sc_hd__a211o_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3252_/S _3196_/B vssd1 vssd1 vccd1 vccd1 _3196_/X sky130_fd_sc_hd__or2_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3282_/A _3048_/X _3049_/Y _3160_/B1 vssd1 vssd1 vccd1 vccd1 _3050_/X sky130_fd_sc_hd__a31o_1
XFILLER_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3952_ _3952_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3883_ _4072_/A _4074_/A vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__or2_2
X_2903_ _3760_/A _2330_/Y _2323_/Y vssd1 vssd1 vccd1 vccd1 _3174_/A sky130_fd_sc_hd__a21o_2
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2834_ _2834_/A _3680_/B _3689_/B _3699_/B vssd1 vssd1 vccd1 vccd1 _3013_/A sky130_fd_sc_hd__nand4_4
X_4504_ _4582_/CLK _4504_/D vssd1 vssd1 vccd1 vccd1 _4504_/Q sky130_fd_sc_hd__dfxtp_1
X_2765_ _2938_/A1 _2760_/X _2764_/X _2751_/X _2756_/X vssd1 vssd1 vccd1 vccd1 _2848_/B
+ sky130_fd_sc_hd__o32ai_4
X_2696_ _4545_/Q _2694_/S _2695_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__a211o_1
X_4435_ _4573_/CLK _4435_/D vssd1 vssd1 vccd1 vccd1 _4435_/Q sky130_fd_sc_hd__dfxtp_1
X_4366_ _4695_/CLK _4366_/D vssd1 vssd1 vccd1 vccd1 _4366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _4379_/Q _4338_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4379_/D sky130_fd_sc_hd__mux2_1
X_4297_ _4296_/X _4672_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4672_/D sky130_fd_sc_hd__mux2_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3255_/S _3247_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3179_ _3278_/A _3177_/Y _3178_/X _3280_/B1 vssd1 vssd1 vccd1 vccd1 _3182_/B sky130_fd_sc_hd__o211a_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2550_ _4470_/Q _4462_/Q _4454_/Q _4446_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2550_/X sky130_fd_sc_hd__mux4_2
XFILLER_5_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2481_ _4573_/Q _2694_/S _2480_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__a211o_1
X_4220_ _4229_/A _4245_/C _4212_/Y _4238_/B vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__a31o_1
X_4151_ _3962_/Y _3963_/X _3973_/A _3974_/Y vssd1 vssd1 vccd1 vccd1 _4151_/X sky130_fd_sc_hd__o211a_1
X_4082_ _4082_/A _4082_/B vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3102_ _3102_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _3102_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3033_ _3261_/A _3032_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3935_ _3935_/A _4672_/Q vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__nand2_2
X_3866_ _4672_/Q _3935_/A vssd1 vssd1 vccd1 vccd1 _3907_/B sky130_fd_sc_hd__and2b_4
X_3797_ _4613_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__or2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2817_ _2817_/A _2885_/B _2848_/A _2817_/D vssd1 vssd1 vccd1 vccd1 _3209_/A sky130_fd_sc_hd__or4_4
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2748_ _4426_/Q _4434_/Q _2800_/S vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__mux2_1
X_2679_ _2677_/X _2678_/X _2614_/S vssd1 vssd1 vccd1 vccd1 _2679_/Y sky130_fd_sc_hd__o21ai_1
X_4418_ _4696_/CLK _4418_/D vssd1 vssd1 vccd1 vccd1 _4418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4349_ _4544_/CLK _4349_/D vssd1 vssd1 vccd1 vccd1 _4349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3720_ _3718_/X _3719_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_40_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4570_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _4592_/Q _4329_/S _3649_/X _3650_/X vssd1 vssd1 vccd1 vccd1 _4592_/D sky130_fd_sc_hd__a22o_1
X_3582_ _2268_/B _2327_/C _3581_/X _2284_/X vssd1 vssd1 vccd1 vccd1 _3628_/A sky130_fd_sc_hd__a2bb2o_1
X_2602_ _4551_/Q _4495_/Q _4487_/Q _4479_/Q _2598_/S _2776_/S1 vssd1 vssd1 vccd1 vccd1
+ _2602_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2533_ _4486_/Q _2761_/S _2532_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__a211o_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _4452_/Q _2809_/S _2461_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__a211o_1
X_4203_ _4264_/B _4201_/X _4202_/Y _4191_/B _4123_/A vssd1 vssd1 vccd1 vccd1 _4203_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ _4647_/Q _2385_/Y _2393_/X vssd1 vssd1 vccd1 vccd1 _2859_/A sky130_fd_sc_hd__o21ai_4
X_4134_ _3872_/Y _4132_/Y _4133_/X vssd1 vssd1 vccd1 vccd1 _4134_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4065_ _3917_/A _3930_/Y _4063_/Y _4229_/A _4123_/A vssd1 vssd1 vccd1 vccd1 _4065_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3016_ _2964_/B _3119_/B _3231_/S vssd1 vssd1 vccd1 vccd1 _3016_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3918_ _2178_/Y _4074_/B _4072_/A vssd1 vssd1 vccd1 vccd1 _4088_/B sky130_fd_sc_hd__o21bai_2
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4689_/CLK sky130_fd_sc_hd__clkbuf_16
X_3849_ _3849_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _4637_/D sky130_fd_sc_hd__nor2_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout131 _2369_/Y vssd1 vssd1 vccd1 vccd1 _2746_/A1 sky130_fd_sc_hd__buf_4
Xfanout120 _3144_/S vssd1 vssd1 vccd1 vccd1 _2805_/C1 sky130_fd_sc_hd__buf_6
XFILLER_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout142 _2758_/C vssd1 vssd1 vccd1 vccd1 _2812_/C sky130_fd_sc_hd__buf_4
Xfanout164 _2513_/B vssd1 vssd1 vccd1 vccd1 _3643_/B sky130_fd_sc_hd__clkbuf_8
Xfanout153 _2863_/B vssd1 vssd1 vccd1 vccd1 _3192_/B sky130_fd_sc_hd__buf_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout186 _2307_/D vssd1 vssd1 vccd1 vccd1 _4256_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout175 _3773_/S vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__buf_8
Xfanout197 _2199_/Y vssd1 vssd1 vccd1 vccd1 _2412_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _4637_/Q vssd1 vssd1 vccd1 vccd1 _2180_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4481_/CLK sky130_fd_sc_hd__clkbuf_16
X_4683_ _4683_/CLK _4683_/D vssd1 vssd1 vccd1 vccd1 _4683_/Q sky130_fd_sc_hd__dfxtp_1
X_3703_ _4491_/Q _3762_/B _3691_/C _3702_/X vssd1 vssd1 vccd1 vccd1 _3703_/X sky130_fd_sc_hd__o31a_1
X_3634_ _3832_/B _3634_/B vssd1 vssd1 vccd1 vccd1 _3634_/Y sky130_fd_sc_hd__nand2_8
X_3565_ _4573_/Q _3565_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4573_/D sky130_fd_sc_hd__mux2_1
X_2516_ _3280_/B1 _2511_/Y _2515_/X _3282_/A vssd1 vssd1 vccd1 vccd1 _2516_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3496_ _4512_/Q _3568_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4512_/D sky130_fd_sc_hd__mux2_1
X_2447_ _4508_/Q _2694_/S _2442_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2447_/X sky130_fd_sc_hd__a211o_1
X_2378_ _4086_/A _3634_/B _3931_/A vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4117_ _4117_/A _4117_/B _4115_/X vssd1 vssd1 vccd1 vccd1 _4117_/X sky130_fd_sc_hd__or3b_1
X_4048_ _3847_/B _3399_/B _3804_/B _4047_/X vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__o211a_1
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3350_ _4406_/Q _4313_/A1 _3355_/S vssd1 vssd1 vccd1 vccd1 _4406_/D sky130_fd_sc_hd__mux2_1
X_2301_ _2473_/B _4046_/B _2360_/A vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__a21o_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _2511_/A _3274_/Y _3280_/Y vssd1 vssd1 vccd1 vccd1 _3282_/C sky130_fd_sc_hd__o21ai_1
X_2232_ _4632_/Q input12/X _4633_/Q vssd1 vssd1 vccd1 vccd1 _2233_/C sky130_fd_sc_hd__a21o_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4573_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2996_ _2996_/A _3068_/A _2886_/A vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__or3b_2
X_4666_ _4667_/CLK _4666_/D vssd1 vssd1 vccd1 vccd1 _4666_/Q sky130_fd_sc_hd__dfxtp_2
X_3617_ _3618_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__or2_1
X_4597_ _4629_/CLK _4597_/D vssd1 vssd1 vccd1 vccd1 _4597_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _4558_/Q _4333_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4558_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3479_ _4497_/Q _3542_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4497_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2850_ _2790_/A _2848_/B _2848_/C vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__a21o_1
X_2781_ _3933_/B _2837_/A vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__or2_1
X_4520_ _4537_/CLK _4520_/D vssd1 vssd1 vccd1 vccd1 _4520_/Q sky130_fd_sc_hd__dfxtp_1
X_4451_ _4555_/CLK _4451_/D vssd1 vssd1 vccd1 vccd1 _4451_/Q sky130_fd_sc_hd__dfxtp_1
X_3402_ _3846_/A _2277_/X _3401_/Y vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__o21ai_4
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4382_ _4582_/CLK _4382_/D vssd1 vssd1 vccd1 vccd1 _4382_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _4391_/Q _4314_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4391_/D sky130_fd_sc_hd__mux2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264_ _4379_/Q _4683_/Q _3264_/S vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__mux2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _3623_/B _4619_/Q _3623_/C _2360_/B vssd1 vssd1 vccd1 vccd1 _2432_/B sky130_fd_sc_hd__or4_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _4506_/Q _4562_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2979_ _4558_/Q _3089_/S _2978_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__a211o_1
X_4649_ _4667_/CLK _4649_/D vssd1 vssd1 vccd1 vccd1 _4649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ _3951_/A _4244_/B vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2902_ _3760_/A _2612_/S _2323_/Y vssd1 vssd1 vccd1 vccd1 _3231_/S sky130_fd_sc_hd__a21oi_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ _3972_/A _4082_/A vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__xor2_4
X_2833_ _2834_/A _3680_/B _3689_/B _3699_/B vssd1 vssd1 vccd1 vccd1 _2904_/B sky130_fd_sc_hd__and4_1
X_2764_ _2814_/A1 _2761_/X _2763_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__o211a_1
X_4503_ _4570_/CLK _4503_/D vssd1 vssd1 vccd1 vccd1 _4503_/Q sky130_fd_sc_hd__dfxtp_1
X_2695_ _4537_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__and3_1
X_4434_ _4580_/CLK _4434_/D vssd1 vssd1 vccd1 vccd1 _4434_/Q sky130_fd_sc_hd__dfxtp_1
X_4365_ _4694_/CLK _4365_/D vssd1 vssd1 vccd1 vccd1 _4365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _4378_/Q _4317_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4378_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ input8/X _4295_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__mux2_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _4571_/Q _4531_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3178_ _4673_/Q _3232_/S vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__or2_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _4517_/Q _2798_/B _2798_/C vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__and3_1
XFILLER_5_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4150_ _3922_/X _4149_/Y _4147_/X _4145_/X vssd1 vssd1 vccd1 vccd1 _4150_/X sky130_fd_sc_hd__o211a_1
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3101_ _3249_/C1 _3088_/X _3092_/X _3100_/X vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__o31ai_4
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4081_ _4081_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _4081_/Y sky130_fd_sc_hd__nand2_1
X_3032_ _4527_/Q _4567_/Q _4559_/Q _4503_/Q _3216_/S _3266_/A1 vssd1 vssd1 vccd1 vccd1
+ _3032_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3934_ _3934_/A _4673_/Q vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__nand2_2
X_3865_ _3935_/A _4672_/Q vssd1 vssd1 vccd1 vccd1 _4188_/B sky130_fd_sc_hd__and2b_4
X_2816_ _2848_/B _2848_/C vssd1 vssd1 vccd1 vccd1 _2817_/D sky130_fd_sc_hd__or2_1
X_3796_ _4605_/Q _4597_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3796_/X sky130_fd_sc_hd__mux2_1
X_2747_ _4353_/Q _3569_/A1 _2857_/S vssd1 vssd1 vccd1 vccd1 _4353_/D sky130_fd_sc_hd__mux2_1
X_2678_ _2904_/A _2678_/B vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__and2_1
X_4417_ _4689_/CLK _4417_/D vssd1 vssd1 vccd1 vccd1 _4417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _4576_/CLK _4348_/D vssd1 vssd1 vccd1 vccd1 _4348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4279_ _4303_/B2 _4277_/X _4278_/Y _3941_/A vssd1 vssd1 vccd1 vccd1 _4279_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3650_ _3731_/A1 _2617_/B _3640_/A _3648_/X vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__o2bb2a_2
X_3581_ _3623_/A _3581_/B _3581_/C _3581_/D vssd1 vssd1 vccd1 vccd1 _3581_/X sky130_fd_sc_hd__and4_1
X_2601_ _2953_/A _2600_/X _2412_/A vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__a21o_1
X_2532_ _4478_/Q _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__and3_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4202_ _3908_/B _4202_/B vssd1 vssd1 vccd1 vccd1 _4202_/Y sky130_fd_sc_hd__nand2b_1
X_2463_ _4468_/Q _2809_/S _2462_/X _2814_/A1 vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__a211o_1
X_2394_ _4647_/Q _2385_/Y _2393_/X vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__o21a_2
X_4133_ _4127_/A _4132_/A _4132_/B _3927_/B vssd1 vssd1 vccd1 vccd1 _4133_/X sky130_fd_sc_hd__a31o_1
XFILLER_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4064_ _2368_/A _4056_/B _4063_/Y vssd1 vssd1 vccd1 vccd1 _4064_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3015_ _3041_/A _3273_/A vssd1 vssd1 vccd1 vccd1 _3176_/A sky130_fd_sc_hd__or2_2
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3917_ _3917_/A _4082_/A vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__nand2_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3848_ _2368_/A _2180_/Y _3848_/S vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__mux2_1
X_3779_ _4607_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__or2_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout121 _2644_/S vssd1 vssd1 vccd1 vccd1 _2814_/A1 sky130_fd_sc_hd__buf_6
Xfanout110 _3251_/S vssd1 vssd1 vccd1 vccd1 _3201_/S sky130_fd_sc_hd__buf_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout165 _2472_/Y vssd1 vssd1 vccd1 vccd1 _2655_/B sky130_fd_sc_hd__buf_6
Xfanout154 _2439_/X vssd1 vssd1 vccd1 vccd1 _2863_/B sky130_fd_sc_hd__buf_4
Xfanout143 _2863_/C vssd1 vssd1 vccd1 vccd1 _2758_/C sky130_fd_sc_hd__buf_4
Xfanout132 _2332_/X vssd1 vssd1 vccd1 vccd1 _3183_/A sky130_fd_sc_hd__buf_4
XFILLER_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout187 _2302_/X vssd1 vssd1 vccd1 vccd1 _2307_/D sky130_fd_sc_hd__buf_4
Xfanout176 _3773_/S vssd1 vssd1 vccd1 vccd1 _3832_/B sky130_fd_sc_hd__buf_8
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout198 _3036_/S vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4682_ _4682_/CLK _4682_/D vssd1 vssd1 vccd1 vccd1 _4682_/Q sky130_fd_sc_hd__dfxtp_1
X_3702_ _3754_/A1 _3700_/Y _3701_/X _3720_/S vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__o22a_1
X_3633_ _3633_/A _3633_/B vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__or2_2
X_3564_ _4572_/Q _3564_/A1 _3571_/S vssd1 vssd1 vccd1 vccd1 _4572_/D sky130_fd_sc_hd__mux2_1
X_2515_ _4071_/A2 _2422_/A _3020_/S _2514_/X vssd1 vssd1 vccd1 vccd1 _2515_/X sky130_fd_sc_hd__a211o_1
X_3495_ _4511_/Q _3567_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4511_/D sky130_fd_sc_hd__mux2_1
X_2446_ _4572_/Q _2694_/S _2445_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__a211o_1
X_4116_ _4116_/A _4119_/A _4116_/C vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__and3_1
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2377_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4047_ _4011_/A _2290_/Y _4046_/Y _3608_/A vssd1 vssd1 vccd1 vccd1 _4047_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2300_ _2300_/A _2300_/B _2300_/C vssd1 vssd1 vccd1 vccd1 _3987_/B sky130_fd_sc_hd__or3_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _2511_/A _3272_/Y _3280_/B1 vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__a21oi_1
X_2231_ _4437_/Q _2286_/C _3581_/D _2206_/X vssd1 vssd1 vccd1 vccd1 _4439_/D sky130_fd_sc_hd__a31o_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2995_ _2995_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _3068_/A sky130_fd_sc_hd__nand2_2
X_4665_ _4665_/CLK _4665_/D vssd1 vssd1 vccd1 vccd1 _4665_/Q sky130_fd_sc_hd__dfxtp_4
X_3616_ _3802_/A _4588_/Q vssd1 vssd1 vccd1 vccd1 _3619_/B sky130_fd_sc_hd__nand2_8
X_4596_ _4626_/CLK _4596_/D vssd1 vssd1 vccd1 vccd1 _4596_/Q sky130_fd_sc_hd__dfxtp_1
X_3547_ _4557_/Q _4312_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4557_/D sky130_fd_sc_hd__mux2_1
X_3478_ _4496_/Q _3541_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4496_/D sky130_fd_sc_hd__mux2_1
X_2429_ _3384_/A _2243_/A _2307_/D _2428_/X vssd1 vssd1 vccd1 vccd1 _3612_/D sky130_fd_sc_hd__o31a_1
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2780_ _2780_/A _3690_/B vssd1 vssd1 vccd1 vccd1 _2780_/Y sky130_fd_sc_hd__xnor2_1
X_4450_ _4553_/CLK _4450_/D vssd1 vssd1 vccd1 vccd1 _4450_/Q sky130_fd_sc_hd__dfxtp_1
X_3401_ _4003_/B _3987_/A vssd1 vssd1 vccd1 vccd1 _3401_/Y sky130_fd_sc_hd__nor2_4
X_4381_ _4678_/CLK _4381_/D vssd1 vssd1 vccd1 vccd1 _4381_/Q sky130_fd_sc_hd__dfxtp_1
X_3332_ _4390_/Q _4313_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4390_/D sky130_fd_sc_hd__mux2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3263_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__inv_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2473_/A _2302_/A vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__nor2_4
X_3194_ _3255_/S _3191_/X _3193_/X _3194_/C1 vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__o211a_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2978_ _4502_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__and3_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4648_ _4667_/CLK _4648_/D vssd1 vssd1 vccd1 vccd1 _4648_/Q sky130_fd_sc_hd__dfxtp_1
X_4579_ _4579_/CLK _4579_/D vssd1 vssd1 vccd1 vccd1 _4579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3950_ _3259_/A _3857_/B _4262_/B vssd1 vssd1 vccd1 vccd1 _3950_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2901_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2913_/B sky130_fd_sc_hd__xnor2_2
X_3881_ _3881_/A _4119_/A vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__and2_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2832_ _3275_/S _2834_/A _3680_/B _3689_/B _3699_/B vssd1 vssd1 vccd1 vccd1 _2832_/X
+ sky130_fd_sc_hd__a41o_1
X_2763_ _4458_/Q _2761_/S _2762_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__a211o_1
X_4502_ _4695_/CLK _4502_/D vssd1 vssd1 vccd1 vccd1 _4502_/Q sky130_fd_sc_hd__dfxtp_1
X_2694_ _4425_/Q _4433_/Q _2694_/S vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4433_ _4537_/CLK _4433_/D vssd1 vssd1 vccd1 vccd1 _4433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4364_ _4697_/CLK _4364_/D vssd1 vssd1 vccd1 vccd1 _4364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4295_ _4660_/Q _4278_/Y _4294_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__a22o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _4377_/Q _4316_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4377_/D sky130_fd_sc_hd__mux2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3252_/S _3246_/B vssd1 vssd1 vccd1 vccd1 _3246_/X sky130_fd_sc_hd__or2_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _3231_/S _3183_/B _3174_/X _3175_/Y vssd1 vssd1 vccd1 vccd1 _3177_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3100_ _3194_/C1 _3095_/X _3099_/X _3257_/A1 vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__a211o_1
XFILLER_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _2617_/B _4079_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3031_ _3028_/X _3029_/X _3030_/X _3266_/A1 _3036_/S vssd1 vssd1 vccd1 vccd1 _3031_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _4662_/Q _3933_/B vssd1 vssd1 vccd1 vccd1 _4261_/B sky130_fd_sc_hd__nand2_2
X_3864_ _3956_/A _3905_/A vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__nand2_2
X_2815_ _2938_/A1 _2810_/X _2814_/X _2801_/X _2806_/X vssd1 vssd1 vccd1 vccd1 _2848_/C
+ sky130_fd_sc_hd__o32ai_4
X_3795_ _3619_/B _3793_/X _3794_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4612_/D sky130_fd_sc_hd__o211a_1
X_2746_ _2746_/A1 _2744_/Y _2794_/B _2743_/X vssd1 vssd1 vccd1 vccd1 _2746_/Y sky130_fd_sc_hd__a31oi_4
X_2677_ _3276_/B _2681_/B _2676_/X _3041_/A vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__o211a_1
X_4416_ _4697_/CLK _4416_/D vssd1 vssd1 vccd1 vccd1 _4416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4347_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4667_/D sky130_fd_sc_hd__and2_1
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4278_ _2368_/B _4278_/B vssd1 vssd1 vccd1 vccd1 _4278_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_100_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3229_ _3229_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3230_/B sky130_fd_sc_hd__xor2_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3580_ _4587_/Q _3580_/A1 _3580_/S vssd1 vssd1 vccd1 vccd1 _4587_/D sky130_fd_sc_hd__mux2_1
X_2600_ _4575_/Q _4519_/Q _4511_/Q _4351_/Q _2892_/S _2893_/A vssd1 vssd1 vccd1 vccd1
+ _2600_/X sky130_fd_sc_hd__mux4_1
X_2531_ _4494_/Q _4550_/Q _2761_/S vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__mux2_1
X_4201_ _3894_/A _4202_/B _3908_/A vssd1 vssd1 vccd1 vccd1 _4201_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2462_ _4460_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__and3_1
X_2393_ _4667_/Q _2847_/A1 _3160_/B1 _3716_/A _2382_/X vssd1 vssd1 vccd1 vccd1 _2393_/X
+ sky130_fd_sc_hd__a221o_2
X_4132_ _4132_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4132_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4063_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _4063_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3014_ _2961_/A _3273_/A _3012_/Y vssd1 vssd1 vccd1 vccd1 _3023_/B sky130_fd_sc_hd__o21a_1
XFILLER_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3916_ _3916_/A _3916_/B vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__nor2_1
X_3847_ _4238_/A _3847_/B _3846_/X vssd1 vssd1 vccd1 vccd1 _3848_/S sky130_fd_sc_hd__or3b_1
X_3778_ _4599_/Q _4591_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__mux2_1
X_2729_ _2961_/A _2783_/A _2728_/X vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout122 _3144_/S vssd1 vssd1 vccd1 vccd1 _2644_/S sky130_fd_sc_hd__buf_4
Xfanout100 _3251_/S vssd1 vssd1 vccd1 vccd1 _2800_/S sky130_fd_sc_hd__buf_4
Xfanout111 _2441_/Y vssd1 vssd1 vccd1 vccd1 _3251_/S sky130_fd_sc_hd__buf_6
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout133 _2330_/Y vssd1 vssd1 vccd1 vccd1 _2612_/S sky130_fd_sc_hd__buf_6
Xfanout144 _2863_/C vssd1 vssd1 vccd1 vccd1 _2990_/C sky130_fd_sc_hd__buf_4
Xfanout155 _2414_/Y vssd1 vssd1 vccd1 vccd1 _3275_/S sky130_fd_sc_hd__buf_6
Xfanout188 _2225_/Y vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__buf_4
Xfanout177 _2241_/Y vssd1 vssd1 vccd1 vccd1 _3773_/S sky130_fd_sc_hd__buf_6
Xfanout166 _4017_/S vssd1 vssd1 vccd1 vccd1 _3691_/C sky130_fd_sc_hd__clkbuf_8
Xfanout199 _3269_/S vssd1 vssd1 vccd1 vccd1 _3036_/S sky130_fd_sc_hd__buf_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4681_ _4681_/CLK _4681_/D vssd1 vssd1 vccd1 vccd1 _4681_/Q sky130_fd_sc_hd__dfxtp_1
X_3701_ _3699_/B _3700_/Y _3727_/S vssd1 vssd1 vccd1 vccd1 _3701_/X sky130_fd_sc_hd__mux2_1
X_3632_ _4010_/A _2331_/A _4013_/S _3633_/B vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__a31o_2
X_3563_ _3563_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3571_/S sky130_fd_sc_hd__and3_4
XFILLER_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2514_ _2904_/A _2512_/X _2513_/Y _2345_/Y vssd1 vssd1 vccd1 vccd1 _2514_/X sky130_fd_sc_hd__o211a_1
X_3494_ _4510_/Q _3566_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4510_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2445_ _4516_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__and3_1
X_4115_ _4119_/A _4116_/C _4116_/A vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__a21o_1
X_2376_ _4050_/C _2375_/X _2306_/A _2473_/C vssd1 vssd1 vccd1 vccd1 _2652_/A sky130_fd_sc_hd__a211o_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4046_ _4046_/A _4046_/B vssd1 vssd1 vccd1 vccd1 _4046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2373_/C _2230_/B vssd1 vssd1 vccd1 vccd1 _2351_/B sky130_fd_sc_hd__or2_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2994_ _2994_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _2994_/Y sky130_fd_sc_hd__xnor2_1
X_4664_ _4672_/CLK _4664_/D vssd1 vssd1 vccd1 vccd1 _4664_/Q sky130_fd_sc_hd__dfxtp_2
X_3615_ _4590_/Q _3617_/B vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__nor2_4
X_4595_ _4629_/CLK _4595_/D vssd1 vssd1 vccd1 vccd1 _4595_/Q sky130_fd_sc_hd__dfxtp_1
X_3546_ _4556_/Q _4320_/A1 _3553_/S vssd1 vssd1 vccd1 vccd1 _4556_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3477_ _4495_/Q _3540_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4495_/D sky130_fd_sc_hd__mux2_1
X_2428_ _3384_/A _3989_/A _4224_/A _2217_/B vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__or4b_2
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2359_ _2290_/Y _2473_/C _2440_/B vssd1 vssd1 vccd1 vccd1 _2860_/D sky130_fd_sc_hd__o21ai_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4029_ _4037_/A _4029_/B vssd1 vssd1 vccd1 vccd1 _4651_/D sky130_fd_sc_hd__and2_1
XFILLER_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3400_ _2293_/A _3991_/B _3399_/X _3771_/S vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__o211ai_4
X_4380_ _4584_/CLK _4380_/D vssd1 vssd1 vccd1 vccd1 _4380_/Q sky130_fd_sc_hd__dfxtp_1
X_3331_ _4389_/Q _4312_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4389_/D sky130_fd_sc_hd__mux2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3262_ _4363_/Q _4587_/Q _3264_/S vssd1 vssd1 vccd1 vccd1 _3263_/A sky130_fd_sc_hd__mux2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _3623_/C _2302_/A vssd1 vssd1 vccd1 vccd1 _2290_/B sky130_fd_sc_hd__nor2_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193_ _4362_/Q _3247_/S _3192_/X _3252_/S vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__a211o_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2977_ _4526_/Q _3089_/S _2976_/X _3086_/A vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__a211o_1
X_4647_ _4665_/CLK _4647_/D vssd1 vssd1 vccd1 vccd1 _4647_/Q sky130_fd_sc_hd__dfxtp_4
X_4578_ _4581_/CLK _4578_/D vssd1 vssd1 vccd1 vccd1 _4578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3529_ _4541_/Q _3565_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4541_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2900_ _3013_/B vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__clkinv_2
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _4082_/A _3972_/A vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__nand2b_4
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2831_ _2825_/X _2827_/X _2830_/X _2898_/A vssd1 vssd1 vccd1 vccd1 _3699_/B sky130_fd_sc_hd__o22a_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2762_ _4450_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__and3_1
X_4501_ _4581_/CLK _4501_/D vssd1 vssd1 vccd1 vccd1 _4501_/Q sky130_fd_sc_hd__dfxtp_1
X_2693_ _4513_/Q _2694_/S _2692_/X _2635_/A vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__a211o_1
X_4432_ _4544_/CLK _4432_/D vssd1 vssd1 vccd1 vccd1 _4432_/Q sky130_fd_sc_hd__dfxtp_1
X_4363_ _4698_/CLK _4363_/D vssd1 vssd1 vccd1 vccd1 _4363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4294_ _4644_/Q _2367_/Y _3629_/Y _4652_/Q vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__a22o_1
X_3314_ _4376_/Q _3577_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4376_/D sky130_fd_sc_hd__mux2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _4507_/Q _4563_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3246_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3176_ _3176_/A _3273_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3223_/A sky130_fd_sc_hd__or3_1
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_52_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4545_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3030_ _4375_/Q _4679_/Q _3216_/S vssd1 vssd1 vccd1 vccd1 _3030_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3932_ _3966_/B _4267_/A2 _4267_/B1 _3855_/B vssd1 vssd1 vccd1 vccd1 _3993_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_43_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4681_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3863_ _3956_/A _3905_/A vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__and2_2
X_2814_ _2814_/A1 _2811_/X _2813_/X _2814_/C1 vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__o211a_1
X_3794_ _4612_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__or2_1
X_2745_ _4488_/Q _4489_/Q _2745_/C vssd1 vssd1 vccd1 vccd1 _2794_/B sky130_fd_sc_hd__or3_4
X_2676_ _2837_/A _2674_/X _2675_/Y _2612_/S vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__a211o_1
X_4415_ _4698_/CLK _4415_/D vssd1 vssd1 vccd1 vccd1 _4415_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4347_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _4666_/D sky130_fd_sc_hd__and2_1
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4277_ _4664_/Q _2367_/Y _3629_/Y _4648_/Q vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__a22o_1
X_3228_ _3185_/A _3211_/B _2382_/X vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3159_ _3288_/A _3158_/X _3154_/Y _2860_/C vssd1 vssd1 vccd1 vccd1 _3159_/X sky130_fd_sc_hd__a211o_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4696_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clkbuf_opt_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4702_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_as1802_283 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_283/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2530_ _2937_/C1 _2523_/X _2525_/X _2984_/B1 vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__a31o_2
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2461_ _4444_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2461_/X sky130_fd_sc_hd__and3_1
X_4200_ _4200_/A _4200_/B vssd1 vssd1 vccd1 vccd1 _4200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2392_ _2858_/A _3328_/B vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__nor2_8
X_4131_ _3935_/A _4267_/A2 _4267_/B1 _4658_/Q _4221_/A vssd1 vssd1 vccd1 vccd1 _4135_/C
+ sky130_fd_sc_hd__a221o_1
X_4062_ _4062_/A _4062_/B vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__and2_4
X_3013_ _3013_/A _3013_/B _3013_/C _3119_/B vssd1 vssd1 vccd1 vccd1 _3273_/A sky130_fd_sc_hd__or4_4
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4667_/CLK sky130_fd_sc_hd__clkbuf_16
X_3915_ _4082_/A _4116_/A vssd1 vssd1 vccd1 vccd1 _3916_/B sky130_fd_sc_hd__and2_1
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3846_ _3846_/A _3846_/B _3930_/A vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__and3_1
X_3777_ _4606_/Q _3741_/S _3776_/X vssd1 vssd1 vccd1 vccd1 _4606_/D sky130_fd_sc_hd__a21o_1
X_2728_ _2414_/Y _2834_/A _3680_/B vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__a21o_1
X_2659_ _2661_/S _4544_/Q vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__and2b_1
Xfanout112 _2936_/C1 vssd1 vssd1 vccd1 vccd1 _2635_/A sky130_fd_sc_hd__buf_6
Xfanout101 _2811_/S vssd1 vssd1 vccd1 vccd1 _2809_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4329_ _4328_/X _4692_/Q _4329_/S vssd1 vssd1 vccd1 vccd1 _4692_/D sky130_fd_sc_hd__mux2_1
Xfanout134 _2323_/Y vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__clkbuf_8
Xfanout123 _3144_/S vssd1 vssd1 vccd1 vccd1 _3255_/S sky130_fd_sc_hd__buf_6
Xfanout145 _2863_/C vssd1 vssd1 vccd1 vccd1 _3192_/C sky130_fd_sc_hd__buf_2
Xfanout156 _2413_/X vssd1 vssd1 vccd1 vccd1 _2961_/A sky130_fd_sc_hd__buf_6
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout178 _3931_/Y vssd1 vssd1 vccd1 vccd1 _4267_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout167 _4017_/S vssd1 vssd1 vccd1 vccd1 _4013_/S sky130_fd_sc_hd__buf_6
Xfanout189 _3771_/S vssd1 vssd1 vccd1 vccd1 _3727_/S sky130_fd_sc_hd__buf_6
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _3716_/A _2848_/C _3699_/Y vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _4683_/CLK _4680_/D vssd1 vssd1 vccd1 vccd1 _4680_/Q sky130_fd_sc_hd__dfxtp_1
X_3631_ _3987_/A _2367_/Y _3633_/B vssd1 vssd1 vccd1 vccd1 _3631_/X sky130_fd_sc_hd__o21ba_4
X_3562_ _4571_/Q _4338_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4571_/D sky130_fd_sc_hd__mux2_1
X_2513_ _2904_/A _2513_/B vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__nand2_1
X_3493_ _4509_/Q _3565_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4509_/D sky130_fd_sc_hd__mux2_1
X_2444_ _4646_/Q _4057_/B _2454_/S vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__mux2_2
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4548_/CLK sky130_fd_sc_hd__clkbuf_16
X_2375_ _3931_/A _4086_/A _2277_/X _3987_/A vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__a211o_1
X_4114_ _4229_/A _4114_/B _4114_/C vssd1 vssd1 vccd1 vccd1 _4123_/C sky130_fd_sc_hd__and3_1
XFILLER_83_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4300_/S _4044_/X _4043_/X _3605_/X vssd1 vssd1 vccd1 vccd1 _4045_/X sky130_fd_sc_hd__o211a_1
XFILLER_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3829_ _3383_/B _4632_/Q input12/X _4062_/A _4631_/Q vssd1 vssd1 vccd1 vccd1 _3829_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2993_ _3257_/A1 _2988_/X _2992_/X _2983_/X _2984_/X vssd1 vssd1 vccd1 vccd1 _3072_/B
+ sky130_fd_sc_hd__o32ai_4
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4663_ _4674_/CLK _4663_/D vssd1 vssd1 vccd1 vccd1 _4663_/Q sky130_fd_sc_hd__dfxtp_1
X_3614_ _3618_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3614_/Y sky130_fd_sc_hd__nand2_1
X_4594_ _4613_/CLK _4594_/D vssd1 vssd1 vccd1 vccd1 _4594_/Q sky130_fd_sc_hd__dfxtp_1
X_3545_ _3563_/A _4319_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _3553_/S sky130_fd_sc_hd__and3_4
X_3476_ _4494_/Q _3539_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4494_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2427_ _2418_/Y _3280_/B1 _2426_/X _2847_/A1 vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2358_ _2360_/B _2473_/C _2357_/Y vssd1 vssd1 vccd1 vccd1 _2440_/B sky130_fd_sc_hd__or3b_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ _4437_/Q _4439_/Q _2265_/Y _3384_/B _4062_/A vssd1 vssd1 vccd1 vccd1 _2289_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4028_ _4667_/Q _4651_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4029_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3330_ _4388_/Q _4331_/A1 _3337_/S vssd1 vssd1 vccd1 vccd1 _4388_/D sky130_fd_sc_hd__mux2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3261_/A _3261_/B vssd1 vssd1 vccd1 vccd1 _3261_/Y sky130_fd_sc_hd__nand2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2212_ _3623_/B _4619_/Q vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__or2_4
X_3192_ _4586_/Q _3192_/B _3192_/C vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__and3_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2976_ _4566_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__and3_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4646_ _4665_/CLK _4646_/D vssd1 vssd1 vccd1 vccd1 _4646_/Q sky130_fd_sc_hd__dfxtp_4
X_4577_ _4579_/CLK _4577_/D vssd1 vssd1 vccd1 vccd1 _4577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3528_ _4540_/Q _3564_/A1 _3535_/S vssd1 vssd1 vccd1 vccd1 _4540_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3459_ _4479_/Q _3540_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4479_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2830_ _2828_/X _2829_/X _4442_/Q vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__mux2_1
X_2761_ _4466_/Q _4474_/Q _2761_/S vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__mux2_1
X_2692_ _4353_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__and3_1
X_4500_ _4580_/CLK _4500_/D vssd1 vssd1 vccd1 vccd1 _4500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4431_ _4543_/CLK _4431_/D vssd1 vssd1 vccd1 vccd1 _4431_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _4675_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4362_ _4683_/CLK _4362_/D vssd1 vssd1 vccd1 vccd1 _4362_/Q sky130_fd_sc_hd__dfxtp_1
X_4293_ _4292_/X _4671_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4671_/D sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _4375_/Q _4314_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4375_/D sky130_fd_sc_hd__mux2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3242_/X _3243_/X _3255_/S vssd1 vssd1 vccd1 vccd1 _3244_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3175_ _3175_/A _3273_/C vssd1 vssd1 vccd1 vccd1 _3175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2959_ _3231_/S _2959_/B _3716_/B vssd1 vssd1 vccd1 vccd1 _2964_/C sky130_fd_sc_hd__or3_1
X_4629_ _4629_/CLK _4629_/D vssd1 vssd1 vccd1 vccd1 _4629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _3931_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _3931_/Y sky130_fd_sc_hd__nor2_2
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3862_ _4673_/Q _3934_/A vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__nand2b_4
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2813_ _4491_/Q _2809_/S _2812_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__a211o_1
X_3793_ _4604_/Q _4596_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__mux2_1
X_2744_ _4488_/Q _2745_/C _4489_/Q vssd1 vssd1 vccd1 vccd1 _2744_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2675_ _4672_/Q _2837_/A vssd1 vssd1 vccd1 vccd1 _2675_/Y sky130_fd_sc_hd__nor2_1
X_4414_ _4695_/CLK _4414_/D vssd1 vssd1 vccd1 vccd1 _4414_/Q sky130_fd_sc_hd__dfxtp_1
X_4345_ _4665_/Q _3417_/S _3409_/Y vssd1 vssd1 vccd1 vccd1 _4665_/D sky130_fd_sc_hd__o21a_1
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4276_ _3608_/A _3633_/A _3832_/X _4275_/X vssd1 vssd1 vccd1 vccd1 _4309_/S sky130_fd_sc_hd__o31ai_4
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3227_ _3290_/A _3227_/B vssd1 vssd1 vccd1 vccd1 _3227_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3158_ _3155_/X _3210_/A vssd1 vssd1 vccd1 vccd1 _3158_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _4680_/Q _4376_/Q _3089_/S vssd1 vssd1 vccd1 vccd1 _3089_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_as1802_284 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_284/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2460_ _2458_/X _2459_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2460_/Y sky130_fd_sc_hd__a21oi_1
X_4130_ _3585_/Y _4177_/B _4127_/A _2371_/C vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__a2bb2o_1
X_2391_ _4644_/Q _2385_/Y _2388_/X vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__o21ai_4
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4061_ _4080_/S _4061_/B vssd1 vssd1 vccd1 vccd1 _4061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3012_ _3119_/A _3119_/B vssd1 vssd1 vccd1 vccd1 _3012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3914_ _4082_/A _4116_/A vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3845_ _3619_/X _3844_/Y _3849_/A vssd1 vssd1 vccd1 vccd1 _4636_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ _2432_/X _3286_/B _3713_/A _3774_/X _3775_/Y vssd1 vssd1 vccd1 vccd1 _3776_/X
+ sky130_fd_sc_hd__o221a_1
X_2727_ _2961_/A _2783_/A vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__nor2_1
X_2658_ _2889_/A _2658_/B vssd1 vssd1 vccd1 vccd1 _2658_/Y sky130_fd_sc_hd__nand2_2
XFILLER_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2589_ _4455_/Q _2761_/S _2588_/X _2641_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__a211o_1
Xfanout113 _2931_/C1 vssd1 vssd1 vccd1 vccd1 _2936_/C1 sky130_fd_sc_hd__buf_6
Xfanout102 _2761_/S vssd1 vssd1 vccd1 vccd1 _2699_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4328_ _3384_/A _4303_/B2 _3587_/A _3390_/B vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__a2bb2o_1
Xfanout146 _2440_/Y vssd1 vssd1 vccd1 vccd1 _2863_/C sky130_fd_sc_hd__buf_4
Xfanout135 _3634_/Y vssd1 vssd1 vccd1 vccd1 _3754_/A1 sky130_fd_sc_hd__buf_6
Xfanout124 _3144_/S vssd1 vssd1 vccd1 vccd1 _3086_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _4264_/A _3903_/X _3904_/Y _3925_/Y vssd1 vssd1 vccd1 vccd1 _4260_/C sky130_fd_sc_hd__a211o_1
Xfanout179 _3877_/Y vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__clkbuf_4
Xfanout157 _3930_/Y vssd1 vssd1 vccd1 vccd1 _4267_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout168 _2368_/X vssd1 vssd1 vccd1 vccd1 _4017_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _3630_/A _3630_/B _3630_/C _3851_/C vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__or4b_4
X_3561_ _4570_/Q _4317_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4570_/D sky130_fd_sc_hd__mux2_1
X_2512_ _2509_/X _2511_/Y _2612_/S vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3492_ _4508_/Q _3564_/A1 _3499_/S vssd1 vssd1 vccd1 vccd1 _4508_/D sky130_fd_sc_hd__mux2_1
X_2443_ _2177_/Y _3993_/A _2454_/S vssd1 vssd1 vccd1 vccd1 _2443_/X sky130_fd_sc_hd__mux2_8
X_2374_ _3993_/B _2384_/C vssd1 vssd1 vccd1 vccd1 _4050_/C sky130_fd_sc_hd__nand2_4
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4113_ _4116_/A _4113_/B vssd1 vssd1 vccd1 vccd1 _4114_/C sky130_fd_sc_hd__or2_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4044_ _4589_/Q _4588_/Q _4590_/Q vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3828_ _3828_/A _3828_/B vssd1 vssd1 vccd1 vccd1 _4630_/D sky130_fd_sc_hd__nand2_1
X_3759_ _4604_/Q _3741_/S _3758_/Y vssd1 vssd1 vccd1 vccd1 _4604_/D sky130_fd_sc_hd__a21o_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ _3086_/A _2989_/X _2991_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__o211a_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4662_ _4662_/CLK _4662_/D vssd1 vssd1 vccd1 vccd1 _4662_/Q sky130_fd_sc_hd__dfxtp_4
X_3613_ _3589_/X _3600_/Y _3613_/C _3613_/D vssd1 vssd1 vccd1 vccd1 _4588_/D sky130_fd_sc_hd__and4bb_1
X_4593_ _4626_/CLK _4593_/D vssd1 vssd1 vccd1 vccd1 _4593_/Q sky130_fd_sc_hd__dfxtp_1
X_3544_ _4555_/Q _3544_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4555_/D sky130_fd_sc_hd__mux2_1
X_3475_ _4493_/Q _3538_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4493_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2426_ _4668_/Q _2422_/A _2422_/Y _3020_/S vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2357_ _2473_/B _4046_/B _3623_/C vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2288_ _4042_/A _4437_/Q vssd1 vssd1 vccd1 vccd1 _2288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4037_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4650_/D sky130_fd_sc_hd__and2_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _4531_/Q _4571_/Q _4563_/Q _4507_/Q _3216_/S _3266_/A1 vssd1 vssd1 vccd1 vccd1
+ _3261_/B sky130_fd_sc_hd__mux4_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2211_ _3623_/B _4619_/Q vssd1 vssd1 vccd1 vccd1 _4046_/B sky130_fd_sc_hd__nand2b_4
X_3191_ _4682_/Q _4378_/Q _3204_/S vssd1 vssd1 vccd1 vccd1 _3191_/X sky130_fd_sc_hd__mux2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _4686_/Q _3080_/C vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__xnor2_1
X_4645_ _4673_/CLK _4645_/D vssd1 vssd1 vccd1 vccd1 _4645_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4576_ _4576_/CLK _4576_/D vssd1 vssd1 vccd1 vccd1 _4576_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _3563_/B _4319_/A _4310_/A vssd1 vssd1 vccd1 vccd1 _3535_/S sky130_fd_sc_hd__and3_4
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3458_ _4478_/Q _3566_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4478_/D sky130_fd_sc_hd__mux2_1
X_3389_ _4050_/A _3623_/C _4046_/B _4062_/A vssd1 vssd1 vccd1 vccd1 _3396_/A sky130_fd_sc_hd__o31a_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2409_ _4468_/Q _4460_/Q _4452_/Q _4444_/Q _2546_/S _2829_/S1 vssd1 vssd1 vccd1 vccd1
+ _2409_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2760_ _2644_/S _2757_/X _2759_/X _2933_/C1 vssd1 vssd1 vccd1 vccd1 _2760_/X sky130_fd_sc_hd__o211a_1
X_2691_ _4577_/Q _2694_/S _2690_/X _2805_/C1 vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__a211o_1
X_4430_ _4574_/CLK _4430_/D vssd1 vssd1 vccd1 vccd1 _4430_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 _2725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4361_ _4681_/CLK _4361_/D vssd1 vssd1 vccd1 vccd1 _4361_/Q sky130_fd_sc_hd__dfxtp_1
X_4292_ input7/X _4291_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__mux2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _4374_/Q _4313_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4374_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _4587_/Q _4363_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3243_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3174_ _3174_/A _3175_/A _3273_/C vssd1 vssd1 vccd1 vccd1 _3174_/X sky130_fd_sc_hd__and3_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2958_ _2959_/B _3716_/B vssd1 vssd1 vccd1 vccd1 _2964_/B sky130_fd_sc_hd__nand2_1
X_4628_ _4630_/CLK _4628_/D vssd1 vssd1 vccd1 vccd1 _4628_/Q sky130_fd_sc_hd__dfxtp_1
X_2889_ _2889_/A _2889_/B vssd1 vssd1 vccd1 vccd1 _2889_/Y sky130_fd_sc_hd__nand2_1
X_4559_ _4570_/CLK _4559_/D vssd1 vssd1 vccd1 vccd1 _4559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3930_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _3930_/Y sky130_fd_sc_hd__nor2_2
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _3934_/A _4673_/Q vssd1 vssd1 vccd1 vccd1 _3956_/A sky130_fd_sc_hd__nand2b_4
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3792_ _3619_/B _3790_/X _3791_/X _3828_/A vssd1 vssd1 vccd1 vccd1 _4611_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2812_ _4483_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2812_/X sky130_fd_sc_hd__and3_1
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2743_ _2364_/Y _2711_/X _2712_/Y _2742_/X vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__o31a_2
X_2674_ _3275_/S _2834_/A _2673_/Y vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__a21o_1
X_4413_ _4694_/CLK _4413_/D vssd1 vssd1 vccd1 vccd1 _4413_/Q sky130_fd_sc_hd__dfxtp_1
X_4344_ _4664_/Q _3417_/S _3405_/X _4037_/A vssd1 vssd1 vccd1 vccd1 _4664_/D sky130_fd_sc_hd__o211a_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _4050_/A _2293_/B _3987_/A _3587_/A _4274_/X vssd1 vssd1 vccd1 vccd1 _4275_/X
+ sky130_fd_sc_hd__o41a_2
X_3226_ _3860_/A _2860_/C _3211_/Y _3225_/Y _2364_/Y vssd1 vssd1 vccd1 vccd1 _3226_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3157_ _3209_/A _3209_/B _3209_/C vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__or3_2
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3088_ _3139_/A _3087_/X _3086_/X _3065_/S vssd1 vssd1 vccd1 vccd1 _3088_/X sky130_fd_sc_hd__o211a_2
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapped_as1802_285 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_285/HI io_out[10] sky130_fd_sc_hd__conb_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _4644_/Q _2385_/Y _2388_/X vssd1 vssd1 vccd1 vccd1 _3298_/B sky130_fd_sc_hd__o21a_4
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4060_ _4224_/A _2996_/A _4059_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__o211a_1
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _3725_/B vssd1 vssd1 vccd1 vccd1 _3119_/B sky130_fd_sc_hd__clkinv_2
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3913_ _4127_/A _4132_/A vssd1 vssd1 vccd1 vccd1 _3913_/Y sky130_fd_sc_hd__nand2_1
X_3844_ _4590_/Q _3614_/Y _4636_/Q vssd1 vssd1 vccd1 vccd1 _3844_/Y sky130_fd_sc_hd__o21ai_1
X_3775_ _3276_/C _3713_/A _3775_/B1 vssd1 vssd1 vccd1 vccd1 _3775_/Y sky130_fd_sc_hd__a21oi_1
X_2726_ _2834_/A _3680_/B vssd1 vssd1 vccd1 vccd1 _2783_/A sky130_fd_sc_hd__nand2_2
X_2657_ _4576_/Q _4520_/Q _4512_/Q _4352_/Q _2661_/S _2825_/B2 vssd1 vssd1 vccd1 vccd1
+ _2658_/B sky130_fd_sc_hd__mux4_2
X_2588_ _4447_/Q _2812_/B _2812_/C vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__and3_1
Xfanout103 _2811_/S vssd1 vssd1 vccd1 vccd1 _2761_/S sky130_fd_sc_hd__buf_6
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout114 _2759_/C1 vssd1 vssd1 vccd1 vccd1 _2641_/S sky130_fd_sc_hd__buf_6
Xfanout125 _2437_/X vssd1 vssd1 vccd1 vccd1 _3144_/S sky130_fd_sc_hd__buf_8
Xfanout136 _3633_/X vssd1 vssd1 vccd1 vccd1 _3666_/B1 sky130_fd_sc_hd__buf_4
Xfanout147 _2927_/B vssd1 vssd1 vccd1 vccd1 _2804_/B sky130_fd_sc_hd__buf_4
X_4327_ _4691_/Q _4338_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4691_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4258_ _4257_/X _4258_/B vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__and2b_1
XFILLER_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout158 _4278_/B vssd1 vssd1 vccd1 vccd1 _4303_/B2 sky130_fd_sc_hd__buf_6
Xfanout169 _2242_/X vssd1 vssd1 vccd1 vccd1 _3762_/B sky130_fd_sc_hd__buf_6
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ _3209_/A _3209_/B _3209_/C _4224_/B vssd1 vssd1 vccd1 vccd1 _3209_/X sky130_fd_sc_hd__or4_1
X_4189_ _4662_/Q _4267_/A2 _4267_/B1 _4660_/Q vssd1 vssd1 vccd1 vccd1 _4191_/B sky130_fd_sc_hd__a22o_1
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3560_ _4569_/Q _4316_/A1 _3562_/S vssd1 vssd1 vccd1 vccd1 _4569_/D sky130_fd_sc_hd__mux2_1
X_2511_ _2511_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__xnor2_1
X_3491_ _3563_/A _3563_/B _4319_/A vssd1 vssd1 vccd1 vccd1 _3499_/S sky130_fd_sc_hd__and3_4
X_2442_ _4348_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2442_/X sky130_fd_sc_hd__and3_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2373_ _3846_/A _2373_/B _2373_/C _3930_/A vssd1 vssd1 vccd1 vccd1 _2373_/Y sky130_fd_sc_hd__nor4_2
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4112_ _4112_/A _4112_/B vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__or2_1
X_4043_ _3618_/A _3604_/A _2274_/A _3802_/A vssd1 vssd1 vccd1 vccd1 _4043_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3827_ _2181_/Y _2182_/Y _3827_/S vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__mux2_1
X_3758_ _3739_/B _3756_/X _3757_/X vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__a21oi_1
X_2709_ _2709_/A _2848_/A vssd1 vssd1 vccd1 vccd1 _2710_/B sky130_fd_sc_hd__nand2_1
X_3689_ _3689_/A _3689_/B vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _4406_/Q _3089_/S _2990_/X _3139_/A vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4661_ _4673_/CLK _4661_/D vssd1 vssd1 vccd1 vccd1 _4661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3612_ _3608_/Y _3610_/Y _3612_/C _3612_/D vssd1 vssd1 vccd1 vccd1 _3613_/D sky130_fd_sc_hd__and4bb_1
X_4592_ _4626_/CLK _4592_/D vssd1 vssd1 vccd1 vccd1 _4592_/Q sky130_fd_sc_hd__dfxtp_1
X_3543_ _4554_/Q _3543_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4554_/D sky130_fd_sc_hd__mux2_1
X_3474_ _4492_/Q _3537_/A1 _3481_/S vssd1 vssd1 vccd1 vccd1 _4492_/D sky130_fd_sc_hd__mux2_1
X_2425_ _2425_/A _2473_/C vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__nor2_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2356_ _3826_/A _2356_/B vssd1 vssd1 vccd1 vccd1 _3259_/B sky130_fd_sc_hd__or2_4
X_2287_ _2234_/X _2269_/X _2275_/X _2286_/X vssd1 vssd1 vccd1 vccd1 _4437_/D sky130_fd_sc_hd__a211o_1
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _4666_/Q _4650_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4027_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _4619_/Q _3623_/B vssd1 vssd1 vccd1 vccd1 _2473_/B sky130_fd_sc_hd__nand2b_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3190_ _4361_/Q _4316_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4361_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2974_ _4357_/Q _4312_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4357_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4644_ _4665_/CLK _4644_/D vssd1 vssd1 vccd1 vccd1 _4644_/Q sky130_fd_sc_hd__dfxtp_4
X_4575_ _4694_/CLK _4575_/D vssd1 vssd1 vccd1 vccd1 _4575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3526_ _4539_/Q _3571_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4539_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3457_ _4477_/Q _3538_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4477_/D sky130_fd_sc_hd__mux2_1
X_3388_ _4046_/B _4011_/A _4046_/A vssd1 vssd1 vccd1 vccd1 _3624_/C sky130_fd_sc_hd__and3b_1
X_2408_ _2953_/A _2404_/Y _2406_/Y _2407_/Y vssd1 vssd1 vccd1 vccd1 _2414_/A sky130_fd_sc_hd__a31o_4
X_2339_ _3383_/B _2339_/B vssd1 vssd1 vccd1 vccd1 _2341_/B sky130_fd_sc_hd__or2_4
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4009_ _4665_/Q _4673_/Q _4013_/S vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2690_ _4521_/Q _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__and3_1
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _3286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _4582_/CLK _4360_/D vssd1 vssd1 vccd1 vccd1 _4360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3311_ _4373_/Q _4312_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4373_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4291_ _4659_/Q _4278_/Y _4290_/X _4303_/B2 vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__a22o_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _4683_/Q _4379_/Q _3247_/S vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3173_/A _3273_/C vssd1 vssd1 vccd1 vccd1 _3183_/B sky130_fd_sc_hd__xnor2_2
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4580_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2957_ _3716_/B vssd1 vssd1 vccd1 vccd1 _3013_/C sky130_fd_sc_hd__inv_2
X_2888_ _4524_/Q _4564_/Q _4556_/Q _4500_/Q _2950_/S _2893_/A vssd1 vssd1 vccd1 vccd1
+ _2889_/B sky130_fd_sc_hd__mux4_1
X_4627_ _4700_/CLK _4627_/D vssd1 vssd1 vccd1 vccd1 _4627_/Q sky130_fd_sc_hd__dfxtp_1
X_4558_ _4695_/CLK _4558_/D vssd1 vssd1 vccd1 vccd1 _4558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3509_ _3563_/A _4310_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3517_/S sky130_fd_sc_hd__and3_4
X_4489_ _4490_/CLK _4489_/D vssd1 vssd1 vccd1 vccd1 _4489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _4679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk _4662_/CLK vssd1 vssd1 vccd1 vccd1 _4629_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _3860_/A _3933_/B vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__nor2_4
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3791_ _4611_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__or2_1
X_2811_ _4499_/Q _4555_/Q _2811_/S vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__mux2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2742_ _2652_/A _2710_/Y _2715_/Y _2655_/Y _2741_/Y vssd1 vssd1 vccd1 vccd1 _2742_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2673_ _3275_/S _2670_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _2673_/Y sky130_fd_sc_hd__a21oi_1
X_4412_ _4694_/CLK _4412_/D vssd1 vssd1 vccd1 vccd1 _4412_/Q sky130_fd_sc_hd__dfxtp_1
X_4343_ _3837_/B _4341_/B _4342_/S _4702_/Q vssd1 vssd1 vccd1 vccd1 _4702_/D sky130_fd_sc_hd__a22o_1
X_4274_ _2243_/A _3396_/B _4045_/X _4047_/X _4273_/X vssd1 vssd1 vccd1 vccd1 _4274_/X
+ sky130_fd_sc_hd__o2111a_1
X_3225_ _2655_/B _3227_/B _2860_/C vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3156_ _4157_/B _4184_/B vssd1 vssd1 vccd1 vccd1 _3209_/C sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_19_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _4672_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3087_ _4504_/Q _4560_/Q _3140_/S vssd1 vssd1 vccd1 vccd1 _3087_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _3989_/A _3989_/B _3989_/C _2425_/A vssd1 vssd1 vccd1 vccd1 _3990_/D sky130_fd_sc_hd__or4b_1
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_as1802_286 vssd1 vssd1 vccd1 vccd1 wrapped_as1802_286/HI io_out[11] sky130_fd_sc_hd__conb_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3010_ _3004_/X _3006_/X _3009_/X _3270_/A vssd1 vssd1 vccd1 vccd1 _3725_/B sky130_fd_sc_hd__o22a_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3912_ _4127_/A _4132_/A vssd1 vssd1 vccd1 vccd1 _3912_/X sky130_fd_sc_hd__or2_1
X_3843_ _4042_/C _3843_/B vssd1 vssd1 vccd1 vccd1 _4635_/D sky130_fd_sc_hd__nand2_1
X_3774_ _3286_/B _3631_/X _3989_/B _3773_/X vssd1 vssd1 vccd1 vccd1 _3774_/X sky130_fd_sc_hd__o22a_1
X_2725_ _2719_/X _2721_/X _2724_/X _2898_/A vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_leaf_8_clk clkbuf_leaf_8_clk/A vssd1 vssd1 vccd1 vccd1 _4684_/CLK sky130_fd_sc_hd__clkbuf_16
X_2656_ _2653_/Y _2654_/X _2655_/Y vssd1 vssd1 vccd1 vccd1 _2656_/Y sky130_fd_sc_hd__a21oi_1
X_2587_ _4463_/Q _4471_/Q _2761_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
Xfanout104 _3251_/S vssd1 vssd1 vccd1 vccd1 _2811_/S sky130_fd_sc_hd__buf_6
Xfanout137 _3633_/X vssd1 vssd1 vccd1 vccd1 _3989_/B sky130_fd_sc_hd__clkbuf_4
Xfanout126 _2424_/X vssd1 vssd1 vccd1 vccd1 _3280_/B1 sky130_fd_sc_hd__buf_6
Xfanout115 _2931_/C1 vssd1 vssd1 vccd1 vccd1 _2759_/C1 sky130_fd_sc_hd__clkbuf_8
X_4326_ _4690_/Q _4337_/A1 _4327_/S vssd1 vssd1 vccd1 vccd1 _4690_/D sky130_fd_sc_hd__mux2_1
X_4257_ _3953_/X _3955_/X _4228_/A _4084_/A vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__a31o_1
Xfanout159 _3385_/Y vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__buf_6
Xfanout148 _2927_/B vssd1 vssd1 vccd1 vccd1 _2798_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4188_ _4205_/A _4188_/B _4188_/C vssd1 vssd1 vccd1 vccd1 _4188_/X sky130_fd_sc_hd__or3_1
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3208_ _3283_/A vssd1 vssd1 vccd1 vccd1 _4224_/B sky130_fd_sc_hd__inv_2
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3139_ _3139_/A _3139_/B vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__or2_1
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2510_ _2511_/A _2513_/B vssd1 vssd1 vccd1 vccd1 _2555_/S sky130_fd_sc_hd__nand2_1
X_3490_ _4507_/Q _4338_/A1 _3490_/S vssd1 vssd1 vccd1 vccd1 _4507_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2441_ _2804_/B _2804_/C vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__nand2_1
X_2372_ _3927_/A _4248_/A _2372_/C vssd1 vssd1 vccd1 vccd1 _3290_/A sky130_fd_sc_hd__or3_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4111_ _4080_/S _2617_/C _4110_/X _3407_/B vssd1 vssd1 vccd1 vccd1 _4111_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4042_ _4042_/A _4692_/Q _4042_/C vssd1 vssd1 vccd1 vccd1 _4042_/X sky130_fd_sc_hd__or3_2
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3826_ _3826_/A _3826_/B vssd1 vssd1 vccd1 vccd1 _4629_/D sky130_fd_sc_hd__or2_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _2431_/Y _4184_/B _3273_/C _3713_/A _3775_/B1 vssd1 vssd1 vccd1 vccd1 _3757_/X
+ sky130_fd_sc_hd__a221o_1
X_2708_ _2817_/A _2708_/B _2848_/A vssd1 vssd1 vccd1 vccd1 _2766_/A sky130_fd_sc_hd__or3_4
X_3688_ _4596_/Q _3741_/S _3687_/X vssd1 vssd1 vccd1 vccd1 _4596_/D sky130_fd_sc_hd__a21bo_1
X_2639_ _4480_/Q _4488_/Q _2699_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4309_ _4308_/X _4675_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4675_/D sky130_fd_sc_hd__mux2_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _4398_/Q _2990_/B _2990_/C vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__and3_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4660_ _4672_/CLK _4660_/D vssd1 vssd1 vccd1 vccd1 _4660_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3611_ _2339_/B _3391_/B _3399_/B _3847_/B vssd1 vssd1 vccd1 vccd1 _3612_/C sky130_fd_sc_hd__a31o_1
X_4591_ _4626_/CLK _4591_/D vssd1 vssd1 vccd1 vccd1 _4591_/Q sky130_fd_sc_hd__dfxtp_1
X_3542_ _4553_/Q _3542_/A1 _3544_/S vssd1 vssd1 vccd1 vccd1 _4553_/D sky130_fd_sc_hd__mux2_1
X_3473_ _3536_/A _4330_/B _4330_/C vssd1 vssd1 vccd1 vccd1 _3481_/S sky130_fd_sc_hd__and3_4
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2424_ _2424_/A _2424_/B vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__or2_2
X_2355_ _3826_/A _2356_/B vssd1 vssd1 vccd1 vccd1 _2860_/C sky130_fd_sc_hd__nor2_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2286_ _2284_/X _3581_/D _2286_/C _4042_/A vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__and4b_1
X_4025_ _4037_/A _4025_/B vssd1 vssd1 vccd1 vccd1 _4649_/D sky130_fd_sc_hd__and2_1
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3809_ _4619_/Q input8/X _3812_/S vssd1 vssd1 vccd1 vccd1 _4619_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _3080_/C _2972_/Y _2970_/X vssd1 vssd1 vccd1 vccd1 _2973_/Y sky130_fd_sc_hd__a21oi_1
X_4643_ _4643_/CLK _4643_/D vssd1 vssd1 vccd1 vccd1 _4643_/Q sky130_fd_sc_hd__dfxtp_4
X_4574_ _4574_/CLK _4574_/D vssd1 vssd1 vccd1 vccd1 _4574_/Q sky130_fd_sc_hd__dfxtp_1
X_3525_ _4538_/Q _3570_/A1 _3526_/S vssd1 vssd1 vccd1 vccd1 _4538_/D sky130_fd_sc_hd__mux2_1
X_3456_ _4476_/Q _3564_/A1 _3463_/S vssd1 vssd1 vccd1 vccd1 _4476_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3387_ _4046_/B _3387_/B vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__or2_4
X_2407_ _2953_/A _2402_/X _2898_/A vssd1 vssd1 vccd1 vccd1 _2407_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2338_ _3581_/B _3385_/B vssd1 vssd1 vccd1 vccd1 _2339_/B sky130_fd_sc_hd__or2_1
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2269_ _2295_/B _2243_/Y _2268_/X vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _4644_/Q _4019_/S _4007_/X _4347_/A vssd1 vssd1 vccd1 vccd1 _4644_/D sky130_fd_sc_hd__o211a_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _3749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _4372_/Q _4320_/A1 _3317_/S vssd1 vssd1 vccd1 vccd1 _4372_/D sky130_fd_sc_hd__mux2_1
X_4290_ _4667_/Q _2367_/Y _3629_/Y _4651_/Q vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__a22o_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3241_ _4362_/Q _4317_/A1 _3297_/S vssd1 vssd1 vccd1 vccd1 _4362_/D sky130_fd_sc_hd__mux2_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3172_ _3173_/A _3273_/C vssd1 vssd1 vccd1 vccd1 _3229_/A sky130_fd_sc_hd__or2_4
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2412_/A _2947_/X _2951_/X _2953_/X _2955_/X vssd1 vssd1 vccd1 vccd1 _3716_/B
+ sky130_fd_sc_hd__o32a_4
X_2887_ _3287_/A _2886_/Y _2655_/Y vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__o21ba_1
X_4626_ _4626_/CLK _4626_/D vssd1 vssd1 vccd1 vccd1 _4626_/Q sky130_fd_sc_hd__dfxtp_1
X_4557_ _4581_/CLK _4557_/D vssd1 vssd1 vccd1 vccd1 _4557_/Q sky130_fd_sc_hd__dfxtp_1
X_4488_ _4551_/CLK _4488_/D vssd1 vssd1 vccd1 vccd1 _4488_/Q sky130_fd_sc_hd__dfxtp_4
X_3508_ _4523_/Q _3571_/A1 _3508_/S vssd1 vssd1 vccd1 vccd1 _4523_/D sky130_fd_sc_hd__mux2_1
X_3439_ _4461_/Q _3538_/A1 _3445_/S vssd1 vssd1 vccd1 vccd1 _4461_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput30 _4701_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_4
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _4603_/Q _4595_/Q _3799_/S vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2810_ _2814_/A1 _2809_/X _2808_/X _2645_/S vssd1 vssd1 vccd1 vccd1 _2810_/X sky130_fd_sc_hd__o211a_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _3282_/A _2740_/X _3239_/A vssd1 vssd1 vccd1 vccd1 _2741_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2672_ _3671_/B _2678_/B _2841_/S vssd1 vssd1 vccd1 vccd1 _2681_/B sky130_fd_sc_hd__mux2_1
X_4411_ _4698_/CLK _4411_/D vssd1 vssd1 vccd1 vccd1 _4411_/Q sky130_fd_sc_hd__dfxtp_1
X_4342_ _3601_/B _4701_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4701_/D sky130_fd_sc_hd__mux2_1
X_4273_ _4062_/B _3847_/B _4042_/X _2189_/Y _3804_/B vssd1 vssd1 vccd1 vccd1 _4273_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3224_ _3770_/S _3761_/B vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__nor2_1
.ends

