magic
tech sky130B
magscale 1 2
timestamp 1674824008
<< viali >>
rect 3433 27557 3467 27591
rect 8585 27557 8619 27591
rect 9321 27557 9355 27591
rect 11897 27557 11931 27591
rect 20821 27557 20855 27591
rect 23305 27557 23339 27591
rect 25789 27557 25823 27591
rect 3985 27421 4019 27455
rect 6561 27421 6595 27455
rect 7205 27421 7239 27455
rect 9137 27421 9171 27455
rect 10425 27421 10459 27455
rect 11713 27421 11747 27455
rect 12633 27421 12667 27455
rect 12817 27421 12851 27455
rect 14289 27421 14323 27455
rect 14933 27421 14967 27455
rect 17049 27421 17083 27455
rect 17509 27421 17543 27455
rect 19625 27421 19659 27455
rect 20085 27421 20119 27455
rect 21465 27421 21499 27455
rect 23949 27421 23983 27455
rect 26433 27421 26467 27455
rect 27721 27421 27755 27455
rect 28365 27421 28399 27455
rect 13277 27353 13311 27387
rect 4169 27285 4203 27319
rect 6745 27285 6779 27319
rect 9873 27285 9907 27319
rect 10885 27285 10919 27319
rect 12817 27285 12851 27319
rect 14473 27285 14507 27319
rect 16865 27285 16899 27319
rect 19441 27285 19475 27319
rect 21281 27285 21315 27319
rect 23765 27285 23799 27319
rect 26249 27285 26283 27319
rect 28181 27285 28215 27319
rect 8861 27081 8895 27115
rect 9505 27013 9539 27047
rect 12265 27013 12299 27047
rect 13921 27013 13955 27047
rect 9321 26945 9355 26979
rect 9597 26945 9631 26979
rect 10793 26945 10827 26979
rect 10977 26945 11011 26979
rect 12081 26945 12115 26979
rect 12357 26945 12391 26979
rect 13001 26945 13035 26979
rect 13829 26945 13863 26979
rect 14105 26945 14139 26979
rect 13093 26877 13127 26911
rect 12081 26809 12115 26843
rect 9321 26741 9355 26775
rect 10057 26741 10091 26775
rect 10977 26741 11011 26775
rect 13277 26741 13311 26775
rect 14105 26741 14139 26775
rect 15853 26741 15887 26775
rect 17049 26741 17083 26775
rect 10609 26537 10643 26571
rect 11161 26537 11195 26571
rect 12357 26537 12391 26571
rect 11529 26401 11563 26435
rect 13001 26401 13035 26435
rect 13369 26401 13403 26435
rect 15117 26401 15151 26435
rect 16589 26401 16623 26435
rect 16773 26401 16807 26435
rect 17785 26401 17819 26435
rect 17969 26401 18003 26435
rect 8401 26333 8435 26367
rect 8585 26333 8619 26367
rect 9413 26333 9447 26367
rect 9597 26333 9631 26367
rect 10425 26333 10459 26367
rect 10609 26333 10643 26367
rect 11069 26333 11103 26367
rect 12081 26333 12115 26367
rect 12357 26333 12391 26367
rect 12909 26333 12943 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 14289 26333 14323 26367
rect 14473 26333 14507 26367
rect 15301 26333 15335 26367
rect 16497 26333 16531 26367
rect 17693 26333 17727 26367
rect 19625 26333 19659 26367
rect 25421 26333 25455 26367
rect 4077 26265 4111 26299
rect 8493 26265 8527 26299
rect 12173 26265 12207 26299
rect 15209 26265 15243 26299
rect 19533 26265 19567 26299
rect 25329 26265 25363 26299
rect 2145 26197 2179 26231
rect 2605 26197 2639 26231
rect 3341 26197 3375 26231
rect 5365 26197 5399 26231
rect 7941 26197 7975 26231
rect 9781 26197 9815 26231
rect 10241 26197 10275 26231
rect 14381 26197 14415 26231
rect 15669 26197 15703 26231
rect 16129 26197 16163 26231
rect 17325 26197 17359 26231
rect 18613 26197 18647 26231
rect 4905 25993 4939 26027
rect 10609 25993 10643 26027
rect 10885 25993 10919 26027
rect 10977 25993 11011 26027
rect 12541 25993 12575 26027
rect 17785 25993 17819 26027
rect 10149 25925 10183 25959
rect 13093 25925 13127 25959
rect 14657 25925 14691 25959
rect 17877 25925 17911 25959
rect 8217 25857 8251 25891
rect 8401 25857 8435 25891
rect 8953 25857 8987 25891
rect 9045 25857 9079 25891
rect 9965 25857 9999 25891
rect 10793 25857 10827 25891
rect 11713 25857 11747 25891
rect 11897 25857 11931 25891
rect 12817 25857 12851 25891
rect 13185 25857 13219 25891
rect 14013 25857 14047 25891
rect 14841 25857 14875 25891
rect 16221 25857 16255 25891
rect 2513 25789 2547 25823
rect 7113 25789 7147 25823
rect 9229 25789 9263 25823
rect 9689 25789 9723 25823
rect 12725 25789 12759 25823
rect 13921 25789 13955 25823
rect 18061 25789 18095 25823
rect 1961 25721 1995 25755
rect 8401 25721 8435 25755
rect 11161 25721 11195 25755
rect 13645 25721 13679 25755
rect 15577 25721 15611 25755
rect 3433 25653 3467 25687
rect 3893 25653 3927 25687
rect 5549 25653 5583 25687
rect 7665 25653 7699 25687
rect 9781 25653 9815 25687
rect 12081 25653 12115 25687
rect 15025 25653 15059 25687
rect 16037 25653 16071 25687
rect 16957 25653 16991 25687
rect 17417 25653 17451 25687
rect 18705 25653 18739 25687
rect 8401 25449 8435 25483
rect 8585 25449 8619 25483
rect 11805 25449 11839 25483
rect 13369 25449 13403 25483
rect 5825 25313 5859 25347
rect 7205 25313 7239 25347
rect 9965 25313 9999 25347
rect 10701 25313 10735 25347
rect 12633 25313 12667 25347
rect 12909 25313 12943 25347
rect 14381 25313 14415 25347
rect 3065 25245 3099 25279
rect 7757 25245 7791 25279
rect 9321 25245 9355 25279
rect 9505 25245 9539 25279
rect 10588 25245 10622 25279
rect 10793 25245 10827 25279
rect 11713 25245 11747 25279
rect 11897 25245 11931 25279
rect 12541 25245 12575 25279
rect 13553 25245 13587 25279
rect 13645 25245 13679 25279
rect 14473 25245 14507 25279
rect 16221 25245 16255 25279
rect 17141 25245 17175 25279
rect 17601 25245 17635 25279
rect 2513 25177 2547 25211
rect 8217 25177 8251 25211
rect 8433 25177 8467 25211
rect 9137 25177 9171 25211
rect 10701 25177 10735 25211
rect 10977 25177 11011 25211
rect 1961 25109 1995 25143
rect 3985 25109 4019 25143
rect 4629 25109 4663 25143
rect 5089 25109 5123 25143
rect 6561 25109 6595 25143
rect 14841 25109 14875 25143
rect 15669 25109 15703 25143
rect 16405 25109 16439 25143
rect 16957 25109 16991 25143
rect 17785 25109 17819 25143
rect 3525 24905 3559 24939
rect 8401 24905 8435 24939
rect 12541 24905 12575 24939
rect 22477 24905 22511 24939
rect 9137 24837 9171 24871
rect 7288 24769 7322 24803
rect 8953 24769 8987 24803
rect 9229 24769 9263 24803
rect 9357 24769 9391 24803
rect 9873 24769 9907 24803
rect 10057 24769 10091 24803
rect 10149 24769 10183 24803
rect 10609 24769 10643 24803
rect 10793 24769 10827 24803
rect 11713 24769 11747 24803
rect 11897 24769 11931 24803
rect 12357 24769 12391 24803
rect 12541 24769 12575 24803
rect 13277 24769 13311 24803
rect 13461 24769 13495 24803
rect 13645 24769 13679 24803
rect 15200 24769 15234 24803
rect 17785 24769 17819 24803
rect 17969 24769 18003 24803
rect 18705 24769 18739 24803
rect 18889 24769 18923 24803
rect 19349 24769 19383 24803
rect 19441 24769 19475 24803
rect 19625 24769 19659 24803
rect 21281 24769 21315 24803
rect 21465 24769 21499 24803
rect 22480 24769 22514 24803
rect 23305 24769 23339 24803
rect 1961 24701 1995 24735
rect 7021 24701 7055 24735
rect 14933 24701 14967 24735
rect 22017 24701 22051 24735
rect 23213 24701 23247 24735
rect 4169 24633 4203 24667
rect 9873 24633 9907 24667
rect 16313 24633 16347 24667
rect 17877 24633 17911 24667
rect 19625 24633 19659 24667
rect 2513 24565 2547 24599
rect 2973 24565 3007 24599
rect 4629 24565 4663 24599
rect 5549 24565 5583 24599
rect 8953 24565 8987 24599
rect 10701 24565 10735 24599
rect 11805 24565 11839 24599
rect 14381 24565 14415 24599
rect 16865 24565 16899 24599
rect 18797 24565 18831 24599
rect 21465 24565 21499 24599
rect 22109 24565 22143 24599
rect 22661 24565 22695 24599
rect 23673 24565 23707 24599
rect 5733 24361 5767 24395
rect 16589 24361 16623 24395
rect 17601 24361 17635 24395
rect 19717 24361 19751 24395
rect 20453 24361 20487 24395
rect 23121 24361 23155 24395
rect 23581 24361 23615 24395
rect 3433 24293 3467 24327
rect 19901 24293 19935 24327
rect 22017 24293 22051 24327
rect 9321 24225 9355 24259
rect 9505 24225 9539 24259
rect 11989 24225 12023 24259
rect 13093 24225 13127 24259
rect 22753 24225 22787 24259
rect 22845 24225 22879 24259
rect 24685 24225 24719 24259
rect 2973 24157 3007 24191
rect 3249 24157 3283 24191
rect 4905 24157 4939 24191
rect 5181 24157 5215 24191
rect 6193 24157 6227 24191
rect 6469 24157 6503 24191
rect 7113 24157 7147 24191
rect 9413 24157 9447 24191
rect 9597 24157 9631 24191
rect 10149 24157 10183 24191
rect 10977 24157 11011 24191
rect 11161 24157 11195 24191
rect 11897 24157 11931 24191
rect 12173 24157 12207 24191
rect 12265 24157 12299 24191
rect 13553 24157 13587 24191
rect 13737 24157 13771 24191
rect 15209 24157 15243 24191
rect 17325 24157 17359 24191
rect 18613 24157 18647 24191
rect 18889 24157 18923 24191
rect 20361 24157 20395 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 21833 24157 21867 24191
rect 22477 24157 22511 24191
rect 22661 24157 22695 24191
rect 22937 24157 22971 24191
rect 23581 24157 23615 24191
rect 23673 24157 23707 24191
rect 24777 24157 24811 24191
rect 3065 24089 3099 24123
rect 6285 24089 6319 24123
rect 7380 24089 7414 24123
rect 10333 24089 10367 24123
rect 15476 24089 15510 24123
rect 19533 24089 19567 24123
rect 19733 24089 19767 24123
rect 1777 24021 1811 24055
rect 2237 24021 2271 24055
rect 4169 24021 4203 24055
rect 4721 24021 4755 24055
rect 5089 24021 5123 24055
rect 6653 24021 6687 24055
rect 8493 24021 8527 24055
rect 9137 24021 9171 24055
rect 10517 24021 10551 24055
rect 10977 24021 11011 24055
rect 12449 24021 12483 24055
rect 13645 24021 13679 24055
rect 14289 24021 14323 24055
rect 17785 24021 17819 24055
rect 18429 24021 18463 24055
rect 18797 24021 18831 24055
rect 23949 24021 23983 24055
rect 25145 24021 25179 24055
rect 5641 23817 5675 23851
rect 9045 23817 9079 23851
rect 10793 23817 10827 23851
rect 15761 23817 15795 23851
rect 16129 23817 16163 23851
rect 17049 23817 17083 23851
rect 17417 23817 17451 23851
rect 18521 23817 18555 23851
rect 20177 23817 20211 23851
rect 21189 23817 21223 23851
rect 1685 23749 1719 23783
rect 1869 23749 1903 23783
rect 9413 23749 9447 23783
rect 14749 23749 14783 23783
rect 18613 23749 18647 23783
rect 21465 23749 21499 23783
rect 2145 23681 2179 23715
rect 4353 23681 4387 23715
rect 5549 23681 5583 23715
rect 5825 23681 5859 23715
rect 6837 23681 6871 23715
rect 9229 23681 9263 23715
rect 9505 23681 9539 23715
rect 10149 23681 10183 23715
rect 10701 23681 10735 23715
rect 10977 23681 11011 23715
rect 12081 23681 12115 23715
rect 12357 23681 12391 23715
rect 12541 23681 12575 23715
rect 13001 23681 13035 23715
rect 15945 23681 15979 23715
rect 16221 23681 16255 23715
rect 17233 23681 17267 23715
rect 17509 23681 17543 23715
rect 19441 23681 19475 23715
rect 20085 23681 20119 23715
rect 20269 23681 20303 23715
rect 21097 23681 21131 23715
rect 21373 23681 21407 23715
rect 22201 23681 22235 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 22845 23681 22879 23715
rect 23397 23681 23431 23715
rect 23581 23681 23615 23715
rect 23673 23681 23707 23715
rect 24317 23681 24351 23715
rect 24501 23681 24535 23715
rect 25053 23681 25087 23715
rect 25237 23681 25271 23715
rect 18337 23613 18371 23647
rect 23489 23613 23523 23647
rect 4997 23545 5031 23579
rect 8125 23545 8159 23579
rect 18981 23545 19015 23579
rect 22845 23545 22879 23579
rect 24317 23545 24351 23579
rect 1869 23477 1903 23511
rect 3065 23477 3099 23511
rect 6009 23477 6043 23511
rect 10057 23477 10091 23511
rect 11161 23477 11195 23511
rect 11897 23477 11931 23511
rect 15209 23477 15243 23511
rect 19533 23477 19567 23511
rect 21281 23477 21315 23511
rect 23857 23477 23891 23511
rect 25145 23477 25179 23511
rect 7481 23273 7515 23307
rect 9137 23273 9171 23307
rect 16405 23273 16439 23307
rect 17325 23273 17359 23307
rect 18061 23273 18095 23307
rect 19441 23273 19475 23307
rect 22937 23273 22971 23307
rect 12449 23205 12483 23239
rect 22109 23205 22143 23239
rect 23397 23205 23431 23239
rect 7021 23137 7055 23171
rect 12173 23137 12207 23171
rect 13277 23137 13311 23171
rect 18429 23137 18463 23171
rect 18521 23137 18555 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 2513 23069 2547 23103
rect 3157 23069 3191 23103
rect 3433 23069 3467 23103
rect 4353 23069 4387 23103
rect 4629 23069 4663 23103
rect 5273 23069 5307 23103
rect 7665 23069 7699 23103
rect 8309 23069 8343 23103
rect 8585 23069 8619 23103
rect 9321 23069 9355 23103
rect 9597 23069 9631 23103
rect 10517 23069 10551 23103
rect 10793 23069 10827 23103
rect 11253 23069 11287 23103
rect 11437 23069 11471 23103
rect 12081 23069 12115 23103
rect 13369 23069 13403 23103
rect 14473 23069 14507 23103
rect 18245 23069 18279 23103
rect 18337 23069 18371 23103
rect 19625 23069 19659 23103
rect 19717 23069 19751 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 20913 23069 20947 23103
rect 21097 23069 21131 23103
rect 21281 23069 21315 23103
rect 21925 23069 21959 23103
rect 22017 23069 22051 23103
rect 22201 23069 22235 23103
rect 22385 23069 22419 23103
rect 22845 23069 22879 23103
rect 23213 23069 23247 23103
rect 23857 23069 23891 23103
rect 24041 23069 24075 23103
rect 26249 23069 26283 23103
rect 14289 23001 14323 23035
rect 15117 23001 15151 23035
rect 25329 23001 25363 23035
rect 2053 22933 2087 22967
rect 2421 22933 2455 22967
rect 2973 22933 3007 22967
rect 3341 22933 3375 22967
rect 4445 22933 4479 22967
rect 4813 22933 4847 22967
rect 8125 22933 8159 22967
rect 8493 22933 8527 22967
rect 9505 22933 9539 22967
rect 10333 22933 10367 22967
rect 10701 22933 10735 22967
rect 11437 22933 11471 22967
rect 13737 22933 13771 22967
rect 14657 22933 14691 22967
rect 21741 22933 21775 22967
rect 23949 22933 23983 22967
rect 25421 22933 25455 22967
rect 25789 22933 25823 22967
rect 26341 22933 26375 22967
rect 7941 22729 7975 22763
rect 8493 22729 8527 22763
rect 9137 22729 9171 22763
rect 9505 22729 9539 22763
rect 13369 22729 13403 22763
rect 14105 22729 14139 22763
rect 20177 22729 20211 22763
rect 22017 22729 22051 22763
rect 22937 22729 22971 22763
rect 4322 22661 4356 22695
rect 6806 22661 6840 22695
rect 8953 22661 8987 22695
rect 9965 22661 9999 22695
rect 10977 22661 11011 22695
rect 18337 22661 18371 22695
rect 18429 22661 18463 22695
rect 18567 22661 18601 22695
rect 21097 22661 21131 22695
rect 2421 22593 2455 22627
rect 2605 22593 2639 22627
rect 2697 22593 2731 22627
rect 3341 22593 3375 22627
rect 3525 22593 3559 22627
rect 3617 22593 3651 22627
rect 4077 22593 4111 22627
rect 9229 22593 9263 22627
rect 9321 22593 9355 22627
rect 10149 22593 10183 22627
rect 10241 22593 10275 22627
rect 10701 22593 10735 22627
rect 10885 22593 10919 22627
rect 11089 22593 11123 22627
rect 11713 22593 11747 22627
rect 11805 22593 11839 22627
rect 11989 22593 12023 22627
rect 13093 22593 13127 22627
rect 13277 22593 13311 22627
rect 13553 22593 13587 22627
rect 14013 22593 14047 22627
rect 14289 22593 14323 22627
rect 15200 22593 15234 22627
rect 17325 22593 17359 22627
rect 18245 22593 18279 22627
rect 19165 22593 19199 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 19901 22593 19935 22627
rect 22201 22593 22235 22627
rect 22845 22593 22879 22627
rect 23029 22593 23063 22627
rect 23581 22593 23615 22627
rect 23857 22593 23891 22627
rect 25237 22593 25271 22627
rect 26157 22593 26191 22627
rect 6561 22525 6595 22559
rect 10977 22525 11011 22559
rect 14933 22525 14967 22559
rect 17509 22525 17543 22559
rect 17601 22525 17635 22559
rect 18705 22525 18739 22559
rect 20177 22525 20211 22559
rect 20637 22525 20671 22559
rect 22385 22525 22419 22559
rect 23673 22525 23707 22559
rect 25421 22525 25455 22559
rect 25513 22525 25547 22559
rect 26065 22525 26099 22559
rect 1777 22457 1811 22491
rect 10241 22457 10275 22491
rect 20729 22457 20763 22491
rect 2237 22389 2271 22423
rect 3157 22389 3191 22423
rect 5457 22389 5491 22423
rect 5917 22389 5951 22423
rect 12173 22389 12207 22423
rect 14473 22389 14507 22423
rect 16313 22389 16347 22423
rect 17141 22389 17175 22423
rect 18061 22389 18095 22423
rect 24041 22389 24075 22423
rect 25053 22389 25087 22423
rect 26433 22389 26467 22423
rect 6009 22185 6043 22219
rect 12725 22185 12759 22219
rect 13737 22185 13771 22219
rect 18245 22185 18279 22219
rect 19441 22185 19475 22219
rect 20729 22185 20763 22219
rect 21281 22185 21315 22219
rect 22017 22185 22051 22219
rect 23765 22185 23799 22219
rect 16405 22117 16439 22151
rect 19717 22117 19751 22151
rect 12725 22049 12759 22083
rect 23765 22049 23799 22083
rect 26525 22049 26559 22083
rect 2053 21981 2087 22015
rect 4077 21981 4111 22015
rect 4344 21981 4378 22015
rect 6469 21981 6503 22015
rect 6736 21981 6770 22015
rect 9137 21981 9171 22015
rect 9321 21981 9355 22015
rect 9505 21981 9539 22015
rect 12633 21981 12667 22015
rect 13553 21981 13587 22015
rect 14289 21981 14323 22015
rect 14381 21981 14415 22015
rect 15025 21981 15059 22015
rect 15292 21981 15326 22015
rect 16865 21981 16899 22015
rect 18705 21981 18739 22015
rect 19625 21981 19659 22015
rect 19809 21981 19843 22015
rect 19901 21981 19935 22015
rect 20085 21981 20119 22015
rect 20545 21981 20579 22015
rect 20729 21981 20763 22015
rect 21189 21981 21223 22015
rect 21373 21981 21407 22015
rect 21833 21981 21867 22015
rect 22017 21981 22051 22015
rect 23673 21981 23707 22015
rect 24593 21981 24627 22015
rect 24686 21981 24720 22015
rect 25058 21981 25092 22015
rect 25697 21981 25731 22015
rect 25881 21981 25915 22015
rect 26709 21981 26743 22015
rect 2320 21913 2354 21947
rect 9413 21913 9447 21947
rect 12173 21913 12207 21947
rect 14565 21913 14599 21947
rect 17132 21913 17166 21947
rect 24869 21913 24903 21947
rect 24961 21913 24995 21947
rect 3433 21845 3467 21879
rect 5457 21845 5491 21879
rect 7849 21845 7883 21879
rect 8585 21845 8619 21879
rect 9689 21845 9723 21879
rect 10885 21845 10919 21879
rect 13001 21845 13035 21879
rect 14466 21845 14500 21879
rect 22477 21845 22511 21879
rect 24041 21845 24075 21879
rect 25237 21845 25271 21879
rect 25789 21845 25823 21879
rect 26617 21845 26651 21879
rect 27077 21845 27111 21879
rect 2237 21641 2271 21675
rect 9321 21641 9355 21675
rect 11161 21641 11195 21675
rect 13093 21641 13127 21675
rect 14105 21641 14139 21675
rect 15577 21641 15611 21675
rect 15945 21641 15979 21675
rect 19073 21641 19107 21675
rect 19257 21641 19291 21675
rect 24409 21641 24443 21675
rect 26433 21641 26467 21675
rect 3157 21573 3191 21607
rect 10048 21573 10082 21607
rect 11980 21573 12014 21607
rect 13737 21573 13771 21607
rect 17132 21573 17166 21607
rect 19717 21573 19751 21607
rect 20177 21573 20211 21607
rect 20729 21573 20763 21607
rect 23397 21573 23431 21607
rect 2053 21505 2087 21539
rect 2329 21505 2363 21539
rect 2973 21505 3007 21539
rect 3249 21505 3283 21539
rect 5825 21505 5859 21539
rect 7205 21505 7239 21539
rect 7389 21505 7423 21539
rect 7481 21505 7515 21539
rect 8197 21505 8231 21539
rect 9781 21505 9815 21539
rect 13921 21505 13955 21539
rect 14841 21505 14875 21539
rect 15025 21505 15059 21539
rect 15761 21505 15795 21539
rect 16037 21505 16071 21539
rect 18705 21505 18739 21539
rect 19901 21505 19935 21539
rect 19993 21505 20027 21539
rect 20637 21505 20671 21539
rect 22845 21505 22879 21539
rect 22937 21505 22971 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 24317 21505 24351 21539
rect 25421 21505 25455 21539
rect 26249 21505 26283 21539
rect 26525 21505 26559 21539
rect 27169 21505 27203 21539
rect 27353 21505 27387 21539
rect 7941 21437 7975 21471
rect 11713 21437 11747 21471
rect 15117 21437 15151 21471
rect 16865 21437 16899 21471
rect 19809 21437 19843 21471
rect 24685 21437 24719 21471
rect 24777 21437 24811 21471
rect 25329 21437 25363 21471
rect 18245 21369 18279 21403
rect 24593 21369 24627 21403
rect 26249 21369 26283 21403
rect 1869 21301 1903 21335
rect 2789 21301 2823 21335
rect 4353 21301 4387 21335
rect 7021 21301 7055 21335
rect 19073 21301 19107 21335
rect 21281 21301 21315 21335
rect 22017 21301 22051 21335
rect 25697 21301 25731 21335
rect 27261 21301 27295 21335
rect 6561 21097 6595 21131
rect 7481 21097 7515 21131
rect 13277 21097 13311 21131
rect 13461 21097 13495 21131
rect 16957 21097 16991 21131
rect 23673 21097 23707 21131
rect 24961 21097 24995 21131
rect 26985 21097 27019 21131
rect 25421 21029 25455 21063
rect 8585 20961 8619 20995
rect 14933 20961 14967 20995
rect 21741 20961 21775 20995
rect 23397 20961 23431 20995
rect 24593 20961 24627 20995
rect 5273 20893 5307 20927
rect 7665 20893 7699 20927
rect 8125 20893 8159 20927
rect 8401 20893 8435 20927
rect 10425 20893 10459 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 14841 20893 14875 20927
rect 18337 20893 18371 20927
rect 20361 20893 20395 20927
rect 23029 20893 23063 20927
rect 23213 20893 23247 20927
rect 23305 20893 23339 20927
rect 23489 20893 23523 20927
rect 24777 20893 24811 20927
rect 25605 20893 25639 20927
rect 25697 20893 25731 20927
rect 26341 20893 26375 20927
rect 26525 20893 26559 20927
rect 27261 20893 27295 20927
rect 27445 20893 27479 20927
rect 27905 20893 27939 20927
rect 28089 20893 28123 20927
rect 1593 20825 1627 20859
rect 4721 20825 4755 20859
rect 9229 20825 9263 20859
rect 13093 20825 13127 20859
rect 13277 20825 13311 20859
rect 15669 20825 15703 20859
rect 19533 20825 19567 20859
rect 22569 20825 22603 20859
rect 25421 20825 25455 20859
rect 26433 20825 26467 20859
rect 2881 20757 2915 20791
rect 4629 20757 4663 20791
rect 8217 20757 8251 20791
rect 9321 20757 9355 20791
rect 11713 20757 11747 20791
rect 14289 20757 14323 20791
rect 18521 20757 18555 20791
rect 19809 20757 19843 20791
rect 20545 20757 20579 20791
rect 27169 20757 27203 20791
rect 27997 20757 28031 20791
rect 3249 20553 3283 20587
rect 8677 20553 8711 20587
rect 12265 20553 12299 20587
rect 22477 20553 22511 20587
rect 27537 20553 27571 20587
rect 2513 20485 2547 20519
rect 2697 20485 2731 20519
rect 3433 20485 3467 20519
rect 3617 20485 3651 20519
rect 8309 20485 8343 20519
rect 8401 20485 8435 20519
rect 10250 20485 10284 20519
rect 14657 20485 14691 20519
rect 15669 20485 15703 20519
rect 16865 20485 16899 20519
rect 25237 20485 25271 20519
rect 27629 20485 27663 20519
rect 1777 20417 1811 20451
rect 2237 20417 2271 20451
rect 4344 20417 4378 20451
rect 7297 20417 7331 20451
rect 7481 20417 7515 20451
rect 7573 20417 7607 20451
rect 8033 20417 8067 20451
rect 8181 20417 8215 20451
rect 8539 20417 8573 20451
rect 10517 20417 10551 20451
rect 10977 20417 11011 20451
rect 11161 20417 11195 20451
rect 11897 20417 11931 20451
rect 12081 20417 12115 20451
rect 12816 20417 12850 20451
rect 13000 20417 13034 20451
rect 14289 20417 14323 20451
rect 15577 20417 15611 20451
rect 15853 20417 15887 20451
rect 19073 20417 19107 20451
rect 19349 20417 19383 20451
rect 19441 20417 19475 20451
rect 19901 20417 19935 20451
rect 20085 20417 20119 20451
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 21189 20417 21223 20451
rect 22017 20417 22051 20451
rect 22937 20417 22971 20451
rect 25145 20417 25179 20451
rect 25329 20417 25363 20451
rect 26249 20417 26283 20451
rect 26433 20417 26467 20451
rect 4077 20349 4111 20383
rect 11805 20349 11839 20383
rect 11989 20349 12023 20383
rect 12908 20349 12942 20383
rect 13093 20349 13127 20383
rect 14197 20349 14231 20383
rect 14565 20349 14599 20383
rect 20637 20349 20671 20383
rect 23857 20349 23891 20383
rect 24685 20349 24719 20383
rect 27445 20349 27479 20383
rect 11161 20281 11195 20315
rect 22293 20281 22327 20315
rect 1593 20213 1627 20247
rect 2513 20213 2547 20247
rect 3433 20213 3467 20247
rect 5457 20213 5491 20247
rect 6009 20213 6043 20247
rect 6561 20213 6595 20247
rect 7113 20213 7147 20247
rect 9137 20213 9171 20247
rect 13277 20213 13311 20247
rect 14013 20213 14047 20247
rect 16037 20213 16071 20247
rect 18153 20213 18187 20247
rect 19901 20213 19935 20247
rect 21281 20213 21315 20247
rect 23029 20213 23063 20247
rect 26341 20213 26375 20247
rect 27997 20213 28031 20247
rect 4537 20009 4571 20043
rect 5733 20009 5767 20043
rect 11713 20009 11747 20043
rect 12081 20009 12115 20043
rect 13369 20009 13403 20043
rect 15485 20009 15519 20043
rect 17877 20009 17911 20043
rect 22201 20009 22235 20043
rect 24041 20009 24075 20043
rect 25329 20009 25363 20043
rect 27905 20009 27939 20043
rect 3433 19941 3467 19975
rect 17325 19941 17359 19975
rect 22017 19941 22051 19975
rect 2053 19873 2087 19907
rect 7573 19873 7607 19907
rect 9505 19873 9539 19907
rect 9689 19873 9723 19907
rect 12541 19873 12575 19907
rect 14933 19873 14967 19907
rect 21741 19873 21775 19907
rect 25973 19873 26007 19907
rect 2320 19805 2354 19839
rect 7021 19805 7055 19839
rect 7849 19805 7883 19839
rect 8033 19805 8067 19839
rect 9413 19805 9447 19839
rect 9597 19805 9631 19839
rect 10885 19805 10919 19839
rect 11713 19805 11747 19839
rect 11805 19805 11839 19839
rect 12633 19805 12667 19839
rect 12909 19805 12943 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14473 19805 14507 19839
rect 14565 19805 14599 19839
rect 14841 19805 14875 19839
rect 15945 19805 15979 19839
rect 16201 19805 16235 19839
rect 18061 19805 18095 19839
rect 18337 19805 18371 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 22753 19805 22787 19839
rect 23029 19805 23063 19839
rect 23489 19805 23523 19839
rect 23581 19805 23615 19839
rect 23765 19805 23799 19839
rect 23857 19805 23891 19839
rect 24593 19805 24627 19839
rect 24777 19805 24811 19839
rect 25237 19805 25271 19839
rect 25421 19805 25455 19839
rect 25881 19805 25915 19839
rect 27077 19805 27111 19839
rect 27445 19805 27479 19839
rect 28181 19805 28215 19839
rect 4353 19737 4387 19771
rect 7731 19737 7765 19771
rect 7940 19737 7974 19771
rect 11253 19737 11287 19771
rect 14289 19737 14323 19771
rect 20453 19737 20487 19771
rect 22937 19737 22971 19771
rect 26893 19737 26927 19771
rect 27905 19737 27939 19771
rect 4537 19669 4571 19703
rect 4721 19669 4755 19703
rect 8217 19669 8251 19703
rect 9873 19669 9907 19703
rect 13737 19669 13771 19703
rect 14749 19669 14783 19703
rect 18245 19669 18279 19703
rect 18797 19669 18831 19703
rect 19441 19669 19475 19703
rect 19809 19669 19843 19703
rect 20545 19669 20579 19703
rect 22851 19669 22885 19703
rect 24685 19669 24719 19703
rect 27169 19669 27203 19703
rect 27261 19669 27295 19703
rect 28089 19669 28123 19703
rect 3433 19465 3467 19499
rect 4261 19465 4295 19499
rect 8033 19465 8067 19499
rect 12725 19465 12759 19499
rect 13461 19465 13495 19499
rect 18429 19465 18463 19499
rect 19165 19465 19199 19499
rect 19717 19465 19751 19499
rect 27537 19465 27571 19499
rect 2320 19397 2354 19431
rect 5365 19397 5399 19431
rect 5457 19397 5491 19431
rect 6920 19397 6954 19431
rect 9505 19397 9539 19431
rect 10333 19397 10367 19431
rect 17316 19397 17350 19431
rect 25145 19397 25179 19431
rect 25329 19397 25363 19431
rect 27169 19397 27203 19431
rect 27369 19397 27403 19431
rect 2053 19329 2087 19363
rect 4169 19329 4203 19363
rect 4445 19329 4479 19363
rect 5273 19329 5307 19363
rect 5641 19329 5675 19363
rect 6653 19329 6687 19363
rect 8677 19329 8711 19363
rect 9137 19329 9171 19363
rect 9230 19329 9264 19363
rect 9413 19329 9447 19363
rect 9643 19329 9677 19363
rect 11713 19329 11747 19363
rect 12357 19329 12391 19363
rect 13829 19329 13863 19363
rect 14473 19329 14507 19363
rect 17049 19329 17083 19363
rect 18981 19329 19015 19363
rect 19257 19329 19291 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 21189 19329 21223 19363
rect 22201 19329 22235 19363
rect 22385 19329 22419 19363
rect 23581 19329 23615 19363
rect 24961 19329 24995 19363
rect 25881 19329 25915 19363
rect 25973 19329 26007 19363
rect 26065 19329 26099 19363
rect 12449 19261 12483 19295
rect 13645 19261 13679 19295
rect 13737 19261 13771 19295
rect 13914 19261 13948 19295
rect 23489 19261 23523 19295
rect 24409 19261 24443 19295
rect 22385 19193 22419 19227
rect 4629 19125 4663 19159
rect 5089 19125 5123 19159
rect 8493 19125 8527 19159
rect 9781 19125 9815 19159
rect 10425 19125 10459 19159
rect 11897 19125 11931 19159
rect 12449 19125 12483 19159
rect 15761 19125 15795 19159
rect 18981 19125 19015 19159
rect 20453 19125 20487 19159
rect 21005 19125 21039 19159
rect 26249 19125 26283 19159
rect 27353 19125 27387 19159
rect 6101 18921 6135 18955
rect 13645 18921 13679 18955
rect 15577 18921 15611 18955
rect 18061 18921 18095 18955
rect 21649 18921 21683 18955
rect 23949 18921 23983 18955
rect 26709 18921 26743 18955
rect 16589 18853 16623 18887
rect 23489 18853 23523 18887
rect 20729 18785 20763 18819
rect 22845 18785 22879 18819
rect 24961 18785 24995 18819
rect 26249 18785 26283 18819
rect 27537 18785 27571 18819
rect 1685 18717 1719 18751
rect 4261 18717 4295 18751
rect 4721 18717 4755 18751
rect 4988 18717 5022 18751
rect 8309 18717 8343 18751
rect 9597 18717 9631 18751
rect 11713 18717 11747 18751
rect 13737 18717 13771 18751
rect 16681 18717 16715 18751
rect 17325 18717 17359 18751
rect 17601 18717 17635 18751
rect 18245 18717 18279 18751
rect 18429 18717 18463 18751
rect 18521 18717 18555 18751
rect 19625 18717 19659 18751
rect 19717 18717 19751 18751
rect 19901 18717 19935 18751
rect 19993 18717 20027 18751
rect 20821 18717 20855 18751
rect 22385 18717 22419 18751
rect 23305 18717 23339 18751
rect 23489 18717 23523 18751
rect 25145 18717 25179 18751
rect 25329 18717 25363 18751
rect 25881 18717 25915 18751
rect 25973 18717 26007 18751
rect 26341 18717 26375 18751
rect 26801 18717 26835 18751
rect 27629 18717 27663 18751
rect 9864 18649 9898 18683
rect 11980 18649 12014 18683
rect 14289 18649 14323 18683
rect 17509 18649 17543 18683
rect 2973 18581 3007 18615
rect 4077 18581 4111 18615
rect 7021 18581 7055 18615
rect 10977 18581 11011 18615
rect 13093 18581 13127 18615
rect 17141 18581 17175 18615
rect 19441 18581 19475 18615
rect 21189 18581 21223 18615
rect 22477 18581 22511 18615
rect 22569 18581 22603 18615
rect 27261 18581 27295 18615
rect 3065 18377 3099 18411
rect 5457 18377 5491 18411
rect 8125 18377 8159 18411
rect 8677 18377 8711 18411
rect 10885 18377 10919 18411
rect 11897 18377 11931 18411
rect 19809 18377 19843 18411
rect 20821 18377 20855 18411
rect 22201 18377 22235 18411
rect 23581 18377 23615 18411
rect 4353 18309 4387 18343
rect 7012 18309 7046 18343
rect 9045 18309 9079 18343
rect 9750 18309 9784 18343
rect 12265 18309 12299 18343
rect 14749 18309 14783 18343
rect 15761 18309 15795 18343
rect 16129 18309 16163 18343
rect 17110 18309 17144 18343
rect 1685 18241 1719 18275
rect 1777 18241 1811 18275
rect 1961 18241 1995 18275
rect 4813 18241 4847 18275
rect 4906 18241 4940 18275
rect 5089 18241 5123 18275
rect 5181 18241 5215 18275
rect 5319 18241 5353 18275
rect 8585 18241 8619 18275
rect 8861 18241 8895 18275
rect 12081 18241 12115 18275
rect 12357 18241 12391 18275
rect 13001 18241 13035 18275
rect 15669 18241 15703 18275
rect 15945 18241 15979 18275
rect 18889 18241 18923 18275
rect 18981 18241 19015 18275
rect 19165 18241 19199 18275
rect 19257 18241 19291 18275
rect 19901 18241 19935 18275
rect 20085 18241 20119 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 21465 18241 21499 18275
rect 22017 18241 22051 18275
rect 22293 18241 22327 18275
rect 22385 18241 22419 18275
rect 23213 18241 23247 18275
rect 23581 18241 23615 18275
rect 26157 18241 26191 18275
rect 27353 18241 27387 18275
rect 6745 18173 6779 18207
rect 9505 18173 9539 18207
rect 16865 18173 16899 18207
rect 18705 18173 18739 18207
rect 23765 18173 23799 18207
rect 25605 18173 25639 18207
rect 26249 18173 26283 18207
rect 27261 18173 27295 18207
rect 22569 18105 22603 18139
rect 24777 18105 24811 18139
rect 27721 18105 27755 18139
rect 2145 18037 2179 18071
rect 5917 18037 5951 18071
rect 18245 18037 18279 18071
rect 24317 18037 24351 18071
rect 3433 17833 3467 17867
rect 6745 17833 6779 17867
rect 13737 17833 13771 17867
rect 21557 17833 21591 17867
rect 25973 17833 26007 17867
rect 26065 17833 26099 17867
rect 27077 17833 27111 17867
rect 9781 17765 9815 17799
rect 16589 17765 16623 17799
rect 23489 17765 23523 17799
rect 9229 17697 9263 17731
rect 17509 17697 17543 17731
rect 19441 17697 19475 17731
rect 23765 17697 23799 17731
rect 24685 17697 24719 17731
rect 26157 17697 26191 17731
rect 2053 17629 2087 17663
rect 2320 17629 2354 17663
rect 3985 17629 4019 17663
rect 4261 17629 4295 17663
rect 4353 17629 4387 17663
rect 7665 17629 7699 17663
rect 7941 17629 7975 17663
rect 8401 17629 8435 17663
rect 8585 17629 8619 17663
rect 9137 17629 9171 17663
rect 9321 17629 9355 17663
rect 9965 17629 9999 17663
rect 10241 17629 10275 17663
rect 12449 17629 12483 17663
rect 13185 17629 13219 17663
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 14565 17629 14599 17663
rect 18245 17629 18279 17663
rect 18337 17629 18371 17663
rect 18613 17629 18647 17663
rect 19625 17629 19659 17663
rect 20637 17629 20671 17663
rect 21557 17629 21591 17663
rect 21961 17629 21995 17663
rect 22661 17629 22695 17663
rect 22937 17629 22971 17663
rect 23397 17629 23431 17663
rect 24593 17629 24627 17663
rect 24777 17629 24811 17663
rect 25881 17629 25915 17663
rect 26985 17629 27019 17663
rect 27169 17629 27203 17663
rect 4169 17561 4203 17595
rect 5273 17561 5307 17595
rect 7849 17561 7883 17595
rect 10149 17561 10183 17595
rect 13369 17561 13403 17595
rect 13461 17561 13495 17595
rect 15301 17561 15335 17595
rect 18797 17561 18831 17595
rect 18889 17561 18923 17595
rect 20269 17561 20303 17595
rect 20453 17561 20487 17595
rect 21741 17561 21775 17595
rect 21833 17561 21867 17595
rect 23489 17561 23523 17595
rect 4537 17493 4571 17527
rect 7481 17493 7515 17527
rect 8493 17493 8527 17527
rect 11161 17493 11195 17527
rect 14381 17493 14415 17527
rect 14749 17493 14783 17527
rect 19809 17493 19843 17527
rect 22477 17493 22511 17527
rect 22845 17493 22879 17527
rect 23581 17493 23615 17527
rect 1685 17289 1719 17323
rect 11069 17289 11103 17323
rect 12541 17289 12575 17323
rect 15301 17289 15335 17323
rect 19349 17289 19383 17323
rect 22217 17289 22251 17323
rect 23489 17289 23523 17323
rect 2412 17221 2446 17255
rect 10701 17221 10735 17255
rect 10885 17221 10919 17255
rect 12173 17221 12207 17255
rect 13001 17221 13035 17255
rect 15945 17221 15979 17255
rect 18705 17221 18739 17255
rect 21373 17221 21407 17255
rect 22017 17221 22051 17255
rect 22937 17221 22971 17255
rect 24501 17221 24535 17255
rect 21143 17187 21177 17221
rect 3985 17153 4019 17187
rect 4629 17153 4663 17187
rect 4896 17153 4930 17187
rect 6561 17153 6595 17187
rect 6654 17153 6688 17187
rect 6837 17153 6871 17187
rect 6929 17153 6963 17187
rect 7067 17153 7101 17187
rect 7849 17153 7883 17187
rect 10057 17153 10091 17187
rect 10241 17153 10275 17187
rect 11897 17153 11931 17187
rect 11990 17153 12024 17187
rect 12273 17153 12307 17187
rect 12403 17153 12437 17187
rect 15209 17153 15243 17187
rect 15393 17153 15427 17187
rect 15853 17153 15887 17187
rect 16129 17153 16163 17187
rect 17121 17153 17155 17187
rect 19073 17153 19107 17187
rect 20085 17153 20119 17187
rect 20361 17153 20395 17187
rect 22845 17153 22879 17187
rect 23029 17153 23063 17187
rect 23857 17153 23891 17187
rect 23949 17153 23983 17187
rect 24685 17153 24719 17187
rect 25329 17153 25363 17187
rect 25513 17153 25547 17187
rect 27261 17153 27295 17187
rect 27445 17153 27479 17187
rect 27905 17153 27939 17187
rect 2145 17085 2179 17119
rect 14749 17085 14783 17119
rect 16865 17085 16899 17119
rect 19165 17085 19199 17119
rect 20177 17085 20211 17119
rect 23673 17085 23707 17119
rect 23765 17085 23799 17119
rect 3525 17017 3559 17051
rect 6009 17017 6043 17051
rect 7205 17017 7239 17051
rect 9137 17017 9171 17051
rect 10057 17017 10091 17051
rect 20269 17017 20303 17051
rect 21005 17017 21039 17051
rect 24869 17017 24903 17051
rect 4169 16949 4203 16983
rect 10885 16949 10919 16983
rect 16313 16949 16347 16983
rect 18245 16949 18279 16983
rect 20545 16949 20579 16983
rect 21189 16949 21223 16983
rect 22201 16949 22235 16983
rect 22385 16949 22419 16983
rect 25697 16949 25731 16983
rect 27353 16949 27387 16983
rect 27997 16949 28031 16983
rect 5549 16745 5583 16779
rect 8401 16745 8435 16779
rect 11345 16745 11379 16779
rect 18521 16745 18555 16779
rect 21373 16745 21407 16779
rect 24593 16745 24627 16779
rect 27813 16745 27847 16779
rect 13737 16677 13771 16711
rect 27905 16677 27939 16711
rect 9321 16609 9355 16643
rect 12725 16609 12759 16643
rect 15301 16609 15335 16643
rect 17141 16609 17175 16643
rect 19625 16609 19659 16643
rect 19717 16609 19751 16643
rect 25421 16609 25455 16643
rect 25605 16609 25639 16643
rect 26065 16609 26099 16643
rect 27997 16609 28031 16643
rect 2053 16541 2087 16575
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4353 16541 4387 16575
rect 7849 16541 7883 16575
rect 7941 16541 7975 16575
rect 8125 16541 8159 16575
rect 8217 16541 8251 16575
rect 14381 16541 14415 16575
rect 14565 16541 14599 16575
rect 15568 16541 15602 16575
rect 17397 16541 17431 16575
rect 20085 16541 20119 16575
rect 20545 16541 20579 16575
rect 20729 16541 20763 16575
rect 21649 16541 21683 16575
rect 22109 16541 22143 16575
rect 22385 16541 22419 16575
rect 23305 16541 23339 16575
rect 23581 16541 23615 16575
rect 25329 16541 25363 16575
rect 25697 16541 25731 16575
rect 26157 16541 26191 16575
rect 26893 16541 26927 16575
rect 27261 16541 27295 16575
rect 27721 16541 27755 16575
rect 2320 16473 2354 16507
rect 4169 16473 4203 16507
rect 7021 16473 7055 16507
rect 9588 16473 9622 16507
rect 12480 16473 12514 16507
rect 13369 16473 13403 16507
rect 13553 16473 13587 16507
rect 21373 16473 21407 16507
rect 22201 16473 22235 16507
rect 26709 16473 26743 16507
rect 3433 16405 3467 16439
rect 4537 16405 4571 16439
rect 10701 16405 10735 16439
rect 14565 16405 14599 16439
rect 16681 16405 16715 16439
rect 19441 16405 19475 16439
rect 19901 16405 19935 16439
rect 19993 16405 20027 16439
rect 20637 16405 20671 16439
rect 21557 16405 21591 16439
rect 22286 16405 22320 16439
rect 23121 16405 23155 16439
rect 23489 16405 23523 16439
rect 26985 16405 27019 16439
rect 27077 16405 27111 16439
rect 2881 16201 2915 16235
rect 9137 16201 9171 16235
rect 10793 16201 10827 16235
rect 14289 16201 14323 16235
rect 16129 16201 16163 16235
rect 16957 16201 16991 16235
rect 18521 16201 18555 16235
rect 22661 16201 22695 16235
rect 27537 16201 27571 16235
rect 1593 16133 1627 16167
rect 6009 16133 6043 16167
rect 10425 16133 10459 16167
rect 13001 16133 13035 16167
rect 15761 16133 15795 16167
rect 21005 16133 21039 16167
rect 22753 16133 22787 16167
rect 26065 16133 26099 16167
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 6837 16065 6871 16099
rect 6929 16065 6963 16099
rect 7849 16065 7883 16099
rect 10149 16065 10183 16099
rect 10297 16065 10331 16099
rect 10517 16065 10551 16099
rect 10655 16065 10689 16099
rect 11713 16065 11747 16099
rect 12173 16065 12207 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 16957 16065 16991 16099
rect 17141 16065 17175 16099
rect 17969 16065 18003 16099
rect 18429 16065 18463 16099
rect 18705 16065 18739 16099
rect 19901 16065 19935 16099
rect 19993 16065 20027 16099
rect 21189 16065 21223 16099
rect 22477 16065 22511 16099
rect 23397 16065 23431 16099
rect 23489 16065 23523 16099
rect 24961 16065 24995 16099
rect 25145 16065 25179 16099
rect 25237 16065 25271 16099
rect 25881 16065 25915 16099
rect 26157 16065 26191 16099
rect 19809 15997 19843 16031
rect 20085 15997 20119 16031
rect 21465 15997 21499 16031
rect 23305 15997 23339 16031
rect 23581 15997 23615 16031
rect 24869 15997 24903 16031
rect 27629 15997 27663 16031
rect 27721 15997 27755 16031
rect 21373 15929 21407 15963
rect 23765 15929 23799 15963
rect 27169 15929 27203 15963
rect 4721 15861 4755 15895
rect 7113 15861 7147 15895
rect 11805 15861 11839 15895
rect 17785 15861 17819 15895
rect 18889 15861 18923 15895
rect 19625 15861 19659 15895
rect 22293 15861 22327 15895
rect 24225 15861 24259 15895
rect 24869 15861 24903 15895
rect 25697 15861 25731 15895
rect 2053 15657 2087 15691
rect 8493 15657 8527 15691
rect 10885 15657 10919 15691
rect 15025 15657 15059 15691
rect 15945 15657 15979 15691
rect 21373 15657 21407 15691
rect 26525 15657 26559 15691
rect 27537 15657 27571 15691
rect 28089 15657 28123 15691
rect 19717 15589 19751 15623
rect 22293 15589 22327 15623
rect 23305 15589 23339 15623
rect 5273 15521 5307 15555
rect 18245 15521 18279 15555
rect 19441 15521 19475 15555
rect 22109 15521 22143 15555
rect 22569 15521 22603 15555
rect 23489 15521 23523 15555
rect 27353 15521 27387 15555
rect 4353 15453 4387 15487
rect 4629 15453 4663 15487
rect 7021 15453 7055 15487
rect 7849 15453 7883 15487
rect 7997 15453 8031 15487
rect 8217 15453 8251 15487
rect 8314 15453 8348 15487
rect 9137 15453 9171 15487
rect 9230 15453 9264 15487
rect 9602 15453 9636 15487
rect 12173 15453 12207 15487
rect 13093 15453 13127 15487
rect 13461 15453 13495 15487
rect 15116 15453 15150 15487
rect 15209 15453 15243 15487
rect 17417 15453 17451 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 18429 15453 18463 15487
rect 20361 15453 20395 15487
rect 20545 15453 20579 15487
rect 21373 15453 21407 15487
rect 21649 15453 21683 15487
rect 23581 15453 23615 15487
rect 23673 15453 23707 15487
rect 23765 15453 23799 15487
rect 24961 15453 24995 15487
rect 25237 15453 25271 15487
rect 25697 15453 25731 15487
rect 25789 15453 25823 15487
rect 25973 15453 26007 15487
rect 26433 15453 26467 15487
rect 26617 15453 26651 15487
rect 27261 15453 27295 15487
rect 28089 15453 28123 15487
rect 28273 15453 28307 15487
rect 3341 15385 3375 15419
rect 4445 15385 4479 15419
rect 8125 15385 8159 15419
rect 9413 15385 9447 15419
rect 9505 15385 9539 15419
rect 13277 15385 13311 15419
rect 20453 15385 20487 15419
rect 21557 15385 21591 15419
rect 24777 15385 24811 15419
rect 25145 15385 25179 15419
rect 4813 15317 4847 15351
rect 9781 15317 9815 15351
rect 14289 15317 14323 15351
rect 18613 15317 18647 15351
rect 19901 15317 19935 15351
rect 25697 15317 25731 15351
rect 1685 15113 1719 15147
rect 6009 15113 6043 15147
rect 8309 15113 8343 15147
rect 10793 15113 10827 15147
rect 13093 15113 13127 15147
rect 15669 15113 15703 15147
rect 16221 15113 16255 15147
rect 20085 15113 20119 15147
rect 21373 15113 21407 15147
rect 22661 15113 22695 15147
rect 23949 15113 23983 15147
rect 25605 15113 25639 15147
rect 27353 15113 27387 15147
rect 4077 15045 4111 15079
rect 6837 15045 6871 15079
rect 10977 15045 11011 15079
rect 14749 15045 14783 15079
rect 19257 15045 19291 15079
rect 22845 15045 22879 15079
rect 25697 15045 25731 15079
rect 25881 15045 25915 15079
rect 1869 14977 1903 15011
rect 4629 14977 4663 15011
rect 4885 14977 4919 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 6929 14977 6963 15011
rect 9597 14977 9631 15011
rect 11980 14977 12014 15011
rect 14013 14977 14047 15011
rect 14565 14977 14599 15011
rect 15393 14977 15427 15011
rect 15577 14977 15611 15011
rect 17049 14977 17083 15011
rect 17325 14977 17359 15011
rect 18337 14977 18371 15011
rect 18429 14977 18463 15011
rect 18613 14977 18647 15011
rect 18797 14977 18831 15011
rect 19533 14977 19567 15011
rect 19993 14977 20027 15011
rect 20177 14977 20211 15011
rect 20821 14977 20855 15011
rect 21281 14977 21315 15011
rect 21465 14977 21499 15011
rect 22569 14977 22603 15011
rect 23305 14977 23339 15011
rect 23949 14977 23983 15011
rect 24133 14977 24167 15011
rect 25605 14977 25639 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 11713 14909 11747 14943
rect 13737 14909 13771 14943
rect 16865 14909 16899 14943
rect 19257 14909 19291 14943
rect 19441 14909 19475 14943
rect 23397 14909 23431 14943
rect 28365 14909 28399 14943
rect 7113 14841 7147 14875
rect 18521 14841 18555 14875
rect 22845 14841 22879 14875
rect 2789 14773 2823 14807
rect 10609 14773 10643 14807
rect 10793 14773 10827 14807
rect 13921 14773 13955 14807
rect 14841 14773 14875 14807
rect 18153 14773 18187 14807
rect 20729 14773 20763 14807
rect 22109 14773 22143 14807
rect 24593 14773 24627 14807
rect 3433 14569 3467 14603
rect 21189 14569 21223 14603
rect 23581 14569 23615 14603
rect 25237 14569 25271 14603
rect 5641 14501 5675 14535
rect 15393 14501 15427 14535
rect 21833 14501 21867 14535
rect 23121 14501 23155 14535
rect 2053 14433 2087 14467
rect 25789 14433 25823 14467
rect 2320 14365 2354 14399
rect 4261 14365 4295 14399
rect 6101 14365 6135 14399
rect 8585 14365 8619 14399
rect 9321 14365 9355 14399
rect 9505 14365 9539 14399
rect 9689 14365 9723 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 13277 14365 13311 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 15945 14365 15979 14399
rect 18245 14365 18279 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 19625 14365 19659 14399
rect 19901 14365 19935 14399
rect 20361 14365 20395 14399
rect 21097 14365 21131 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22845 14365 22879 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 4528 14297 4562 14331
rect 9413 14297 9447 14331
rect 10609 14297 10643 14331
rect 14657 14297 14691 14331
rect 16221 14297 16255 14331
rect 18521 14297 18555 14331
rect 19809 14297 19843 14331
rect 20453 14297 20487 14331
rect 20637 14297 20671 14331
rect 23121 14297 23155 14331
rect 7389 14229 7423 14263
rect 8401 14229 8435 14263
rect 9137 14229 9171 14263
rect 11897 14229 11931 14263
rect 12817 14229 12851 14263
rect 17693 14229 17727 14263
rect 18797 14229 18831 14263
rect 19901 14229 19935 14263
rect 20361 14229 20395 14263
rect 22937 14229 22971 14263
rect 24593 14229 24627 14263
rect 1869 14025 1903 14059
rect 7297 14025 7331 14059
rect 10057 14025 10091 14059
rect 10425 14025 10459 14059
rect 11069 14025 11103 14059
rect 13093 14025 13127 14059
rect 14657 14025 14691 14059
rect 16957 14025 16991 14059
rect 19993 14025 20027 14059
rect 9597 13957 9631 13991
rect 11980 13957 12014 13991
rect 13921 13957 13955 13991
rect 16238 13957 16272 13991
rect 17693 13957 17727 13991
rect 19625 13957 19659 13991
rect 25697 13957 25731 13991
rect 1777 13889 1811 13923
rect 1961 13889 1995 13923
rect 2677 13889 2711 13923
rect 4445 13889 4479 13923
rect 4701 13889 4735 13923
rect 6653 13889 6687 13923
rect 6746 13889 6780 13923
rect 6929 13889 6963 13923
rect 7029 13889 7063 13923
rect 7159 13889 7193 13923
rect 10241 13889 10275 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 11161 13889 11195 13923
rect 13737 13889 13771 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 15945 13889 15979 13923
rect 16042 13889 16076 13923
rect 16865 13889 16899 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 19533 13889 19567 13923
rect 19809 13889 19843 13923
rect 22477 13889 22511 13923
rect 23213 13889 23247 13923
rect 24225 13889 24259 13923
rect 25053 13889 25087 13923
rect 25237 13889 25271 13923
rect 2421 13821 2455 13855
rect 11713 13821 11747 13855
rect 19073 13821 19107 13855
rect 20545 13821 20579 13855
rect 23305 13821 23339 13855
rect 24317 13821 24351 13855
rect 3801 13753 3835 13787
rect 18061 13753 18095 13787
rect 20821 13753 20855 13787
rect 23581 13753 23615 13787
rect 24593 13753 24627 13787
rect 5825 13685 5859 13719
rect 8309 13685 8343 13719
rect 13553 13685 13587 13719
rect 21005 13685 21039 13719
rect 22385 13685 22419 13719
rect 25145 13685 25179 13719
rect 3433 13481 3467 13515
rect 7941 13481 7975 13515
rect 11713 13481 11747 13515
rect 12633 13481 12667 13515
rect 13645 13481 13679 13515
rect 14565 13481 14599 13515
rect 16208 13481 16242 13515
rect 19809 13481 19843 13515
rect 21005 13481 21039 13515
rect 24593 13481 24627 13515
rect 8493 13413 8527 13447
rect 18797 13413 18831 13447
rect 21741 13413 21775 13447
rect 19717 13345 19751 13379
rect 24961 13345 24995 13379
rect 2053 13277 2087 13311
rect 3985 13277 4019 13311
rect 4721 13277 4755 13311
rect 6561 13277 6595 13311
rect 6828 13277 6862 13311
rect 8401 13277 8435 13311
rect 9137 13277 9171 13311
rect 9230 13277 9264 13311
rect 9602 13277 9636 13311
rect 10425 13277 10459 13311
rect 12817 13277 12851 13311
rect 13093 13277 13127 13311
rect 13553 13277 13587 13311
rect 14381 13277 14415 13311
rect 14657 13277 14691 13311
rect 15945 13277 15979 13311
rect 18613 13277 18647 13311
rect 19441 13277 19475 13311
rect 20545 13277 20579 13311
rect 20821 13277 20855 13311
rect 21465 13277 21499 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22569 13277 22603 13311
rect 24777 13277 24811 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 25605 13277 25639 13311
rect 25973 13277 26007 13311
rect 2298 13209 2332 13243
rect 4988 13209 5022 13243
rect 9413 13209 9447 13243
rect 9505 13209 9539 13243
rect 15117 13209 15151 13243
rect 15301 13209 15335 13243
rect 17969 13209 18003 13243
rect 20637 13209 20671 13243
rect 22836 13209 22870 13243
rect 25789 13209 25823 13243
rect 26433 13209 26467 13243
rect 4169 13141 4203 13175
rect 6101 13141 6135 13175
rect 9781 13141 9815 13175
rect 13001 13141 13035 13175
rect 15485 13141 15519 13175
rect 19993 13141 20027 13175
rect 23949 13141 23983 13175
rect 1869 12937 1903 12971
rect 3065 12937 3099 12971
rect 8309 12937 8343 12971
rect 11161 12937 11195 12971
rect 12265 12937 12299 12971
rect 15393 12937 15427 12971
rect 19441 12937 19475 12971
rect 19993 12937 20027 12971
rect 23213 12937 23247 12971
rect 1685 12869 1719 12903
rect 4353 12869 4387 12903
rect 5825 12869 5859 12903
rect 6009 12869 6043 12903
rect 7113 12869 7147 12903
rect 9597 12869 9631 12903
rect 13001 12869 13035 12903
rect 16313 12869 16347 12903
rect 18061 12869 18095 12903
rect 2145 12801 2179 12835
rect 4813 12801 4847 12835
rect 6883 12801 6917 12835
rect 7021 12801 7055 12835
rect 7296 12801 7330 12835
rect 7389 12801 7423 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 12265 12801 12299 12835
rect 12541 12801 12575 12835
rect 15209 12801 15243 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 16957 12801 16991 12835
rect 17141 12801 17175 12835
rect 17693 12801 17727 12835
rect 17877 12801 17911 12835
rect 18521 12801 18555 12835
rect 19245 12801 19279 12835
rect 21106 12801 21140 12835
rect 22017 12801 22051 12835
rect 23397 12801 23431 12835
rect 23489 12801 23523 12835
rect 23581 12801 23615 12835
rect 23699 12801 23733 12835
rect 24501 12801 24535 12835
rect 25513 12801 25547 12835
rect 16865 12733 16899 12767
rect 21373 12733 21407 12767
rect 22293 12733 22327 12767
rect 23857 12733 23891 12767
rect 24409 12733 24443 12767
rect 24593 12733 24627 12767
rect 24685 12733 24719 12767
rect 25697 12733 25731 12767
rect 26157 12733 26191 12767
rect 5641 12665 5675 12699
rect 6745 12665 6779 12699
rect 22201 12665 22235 12699
rect 1869 12597 1903 12631
rect 4997 12597 5031 12631
rect 5825 12597 5859 12631
rect 10057 12597 10091 12631
rect 14473 12597 14507 12631
rect 18705 12597 18739 12631
rect 22109 12597 22143 12631
rect 24869 12597 24903 12631
rect 25329 12597 25363 12631
rect 2053 12393 2087 12427
rect 6745 12393 6779 12427
rect 11621 12393 11655 12427
rect 18705 12393 18739 12427
rect 20637 12393 20671 12427
rect 22385 12393 22419 12427
rect 23581 12393 23615 12427
rect 7205 12325 7239 12359
rect 12633 12325 12667 12359
rect 13645 12325 13679 12359
rect 21373 12325 21407 12359
rect 25697 12325 25731 12359
rect 15669 12257 15703 12291
rect 19441 12257 19475 12291
rect 20085 12257 20119 12291
rect 20361 12257 20395 12291
rect 3433 12189 3467 12223
rect 6193 12189 6227 12223
rect 6561 12189 6595 12223
rect 8585 12189 8619 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 13369 12189 13403 12223
rect 13645 12189 13679 12223
rect 14565 12189 14599 12223
rect 14749 12189 14783 12223
rect 15393 12189 15427 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 19993 12189 20027 12223
rect 20453 12189 20487 12223
rect 21097 12189 21131 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 23121 12189 23155 12223
rect 23397 12189 23431 12223
rect 24961 12189 24995 12223
rect 25053 12189 25087 12223
rect 25973 12189 26007 12223
rect 3188 12121 3222 12155
rect 3985 12121 4019 12155
rect 6377 12121 6411 12155
rect 6469 12121 6503 12155
rect 8318 12121 8352 12155
rect 10333 12121 10367 12155
rect 14381 12121 14415 12155
rect 18061 12121 18095 12155
rect 18889 12121 18923 12155
rect 24593 12121 24627 12155
rect 24685 12121 24719 12155
rect 25697 12121 25731 12155
rect 25881 12121 25915 12155
rect 5273 12053 5307 12087
rect 9597 12053 9631 12087
rect 17141 12053 17175 12087
rect 18521 12053 18555 12087
rect 18689 12053 18723 12087
rect 20269 12053 20303 12087
rect 21833 12053 21867 12087
rect 23213 12053 23247 12087
rect 25237 12053 25271 12087
rect 2145 11849 2179 11883
rect 3985 11849 4019 11883
rect 10701 11849 10735 11883
rect 11989 11849 12023 11883
rect 19165 11849 19199 11883
rect 21373 11849 21407 11883
rect 24777 11849 24811 11883
rect 26341 11849 26375 11883
rect 1777 11781 1811 11815
rect 6653 11781 6687 11815
rect 12173 11781 12207 11815
rect 13461 11781 13495 11815
rect 15853 11781 15887 11815
rect 16221 11781 16255 11815
rect 19809 11781 19843 11815
rect 23664 11781 23698 11815
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 2872 11713 2906 11747
rect 4896 11713 4930 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 8594 11713 8628 11747
rect 9321 11713 9355 11747
rect 9588 11713 9622 11747
rect 12633 11713 12667 11747
rect 19165 11713 19199 11747
rect 20729 11713 20763 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 22753 11713 22787 11747
rect 25513 11713 25547 11747
rect 25605 11713 25639 11747
rect 25789 11713 25823 11747
rect 2605 11645 2639 11679
rect 4629 11645 4663 11679
rect 7021 11645 7055 11679
rect 8861 11645 8895 11679
rect 13185 11645 13219 11679
rect 15209 11645 15243 11679
rect 16865 11645 16899 11679
rect 17141 11645 17175 11679
rect 18613 11645 18647 11679
rect 20269 11645 20303 11679
rect 23397 11645 23431 11679
rect 25697 11645 25731 11679
rect 20177 11577 20211 11611
rect 20821 11577 20855 11611
rect 25329 11577 25363 11611
rect 6009 11509 6043 11543
rect 7481 11509 7515 11543
rect 11805 11509 11839 11543
rect 11989 11509 12023 11543
rect 22109 11509 22143 11543
rect 22845 11509 22879 11543
rect 2053 11305 2087 11339
rect 5733 11305 5767 11339
rect 8585 11305 8619 11339
rect 14979 11305 15013 11339
rect 19901 11305 19935 11339
rect 21649 11305 21683 11339
rect 22845 11305 22879 11339
rect 23949 11305 23983 11339
rect 25145 11305 25179 11339
rect 10885 11237 10919 11271
rect 13461 11237 13495 11271
rect 17877 11237 17911 11271
rect 21005 11237 21039 11271
rect 25697 11237 25731 11271
rect 9505 11169 9539 11203
rect 11989 11169 12023 11203
rect 15669 11169 15703 11203
rect 18429 11169 18463 11203
rect 19993 11169 20027 11203
rect 24869 11169 24903 11203
rect 4353 11101 4387 11135
rect 8401 11101 8435 11135
rect 11713 11101 11747 11135
rect 15209 11101 15243 11135
rect 18245 11101 18279 11135
rect 18337 11101 18371 11135
rect 20177 11101 20211 11135
rect 21097 11101 21131 11135
rect 21557 11101 21591 11135
rect 21741 11101 21775 11135
rect 22201 11101 22235 11135
rect 22385 11101 22419 11135
rect 23673 11101 23707 11135
rect 23949 11101 23983 11135
rect 24777 11101 24811 11135
rect 25605 11101 25639 11135
rect 25789 11101 25823 11135
rect 26801 11101 26835 11135
rect 3341 11033 3375 11067
rect 4620 11033 4654 11067
rect 6193 11033 6227 11067
rect 9750 11033 9784 11067
rect 17417 11033 17451 11067
rect 19901 11033 19935 11067
rect 26249 11033 26283 11067
rect 7481 10965 7515 10999
rect 20361 10965 20395 10999
rect 22293 10965 22327 10999
rect 23765 10965 23799 10999
rect 2145 10761 2179 10795
rect 3065 10761 3099 10795
rect 4997 10761 5031 10795
rect 5549 10761 5583 10795
rect 5917 10761 5951 10795
rect 7021 10761 7055 10795
rect 7573 10761 7607 10795
rect 12817 10761 12851 10795
rect 19625 10761 19659 10795
rect 21005 10761 21039 10795
rect 21465 10761 21499 10795
rect 24317 10761 24351 10795
rect 1777 10693 1811 10727
rect 8708 10693 8742 10727
rect 11161 10693 11195 10727
rect 13277 10693 13311 10727
rect 16865 10693 16899 10727
rect 23489 10693 23523 10727
rect 25513 10693 25547 10727
rect 1685 10625 1719 10659
rect 1961 10625 1995 10659
rect 4353 10625 4387 10659
rect 4905 10625 4939 10659
rect 5089 10625 5123 10659
rect 5733 10625 5767 10659
rect 6009 10625 6043 10659
rect 6837 10625 6871 10659
rect 7113 10625 7147 10659
rect 8953 10625 8987 10659
rect 9413 10625 9447 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 12633 10625 12667 10659
rect 19073 10625 19107 10659
rect 19441 10625 19475 10659
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 21097 10625 21131 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 23397 10625 23431 10659
rect 24041 10625 24075 10659
rect 25053 10625 25087 10659
rect 16037 10557 16071 10591
rect 16313 10557 16347 10591
rect 20913 10557 20947 10591
rect 24317 10557 24351 10591
rect 24777 10557 24811 10591
rect 12173 10489 12207 10523
rect 22753 10489 22787 10523
rect 24133 10489 24167 10523
rect 26065 10489 26099 10523
rect 6653 10421 6687 10455
rect 14565 10421 14599 10455
rect 18153 10421 18187 10455
rect 19349 10421 19383 10455
rect 20085 10421 20119 10455
rect 22017 10421 22051 10455
rect 24869 10421 24903 10455
rect 24961 10421 24995 10455
rect 1869 10217 1903 10251
rect 4261 10217 4295 10251
rect 6561 10217 6595 10251
rect 7665 10217 7699 10251
rect 12449 10217 12483 10251
rect 16681 10217 16715 10251
rect 19717 10217 19751 10251
rect 21097 10217 21131 10251
rect 21833 10217 21867 10251
rect 24593 10217 24627 10251
rect 24777 10217 24811 10251
rect 26709 10217 26743 10251
rect 8125 10149 8159 10183
rect 9229 10149 9263 10183
rect 21649 10149 21683 10183
rect 23029 10149 23063 10183
rect 25421 10149 25455 10183
rect 27261 10149 27295 10183
rect 14381 10081 14415 10115
rect 16129 10081 16163 10115
rect 17233 10081 17267 10115
rect 18337 10081 18371 10115
rect 23581 10081 23615 10115
rect 3341 10013 3375 10047
rect 4445 10013 4479 10047
rect 4721 10013 4755 10047
rect 5273 10013 5307 10047
rect 7481 10009 7515 10043
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 13737 10013 13771 10047
rect 18061 10013 18095 10047
rect 19901 10013 19935 10047
rect 20085 10013 20119 10047
rect 20821 10013 20855 10047
rect 20913 10013 20947 10047
rect 21189 10013 21223 10047
rect 21833 10013 21867 10047
rect 21925 10013 21959 10047
rect 22753 10013 22787 10047
rect 23673 10013 23707 10047
rect 25697 10013 25731 10047
rect 4629 9945 4663 9979
rect 8493 9945 8527 9979
rect 9781 9945 9815 9979
rect 11529 9945 11563 9979
rect 14657 9945 14691 9979
rect 17141 9945 17175 9979
rect 20177 9945 20211 9979
rect 22109 9945 22143 9979
rect 23029 9945 23063 9979
rect 24761 9945 24795 9979
rect 24961 9945 24995 9979
rect 25421 9945 25455 9979
rect 17049 9877 17083 9911
rect 20637 9877 20671 9911
rect 22845 9877 22879 9911
rect 24041 9877 24075 9911
rect 25605 9877 25639 9911
rect 26249 9877 26283 9911
rect 7941 9673 7975 9707
rect 14657 9673 14691 9707
rect 18337 9673 18371 9707
rect 18705 9673 18739 9707
rect 26065 9673 26099 9707
rect 4629 9605 4663 9639
rect 4997 9605 5031 9639
rect 5825 9605 5859 9639
rect 6009 9605 6043 9639
rect 8769 9605 8803 9639
rect 17509 9605 17543 9639
rect 18797 9605 18831 9639
rect 21189 9605 21223 9639
rect 23489 9605 23523 9639
rect 2053 9537 2087 9571
rect 2320 9537 2354 9571
rect 3985 9537 4019 9571
rect 4813 9537 4847 9571
rect 5089 9537 5123 9571
rect 6828 9537 6862 9571
rect 8585 9537 8619 9571
rect 8861 9537 8895 9571
rect 11805 9537 11839 9571
rect 12081 9537 12115 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 13369 9537 13403 9571
rect 16129 9537 16163 9571
rect 17877 9537 17911 9571
rect 22201 9537 22235 9571
rect 23121 9537 23155 9571
rect 23213 9537 23247 9571
rect 23397 9537 23431 9571
rect 23581 9537 23615 9571
rect 24409 9537 24443 9571
rect 24593 9537 24627 9571
rect 24685 9537 24719 9571
rect 25421 9537 25455 9571
rect 6561 9469 6595 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 11161 9469 11195 9503
rect 15853 9469 15887 9503
rect 18889 9469 18923 9503
rect 19717 9469 19751 9503
rect 21465 9469 21499 9503
rect 22109 9469 22143 9503
rect 22293 9469 22327 9503
rect 22385 9469 22419 9503
rect 25237 9469 25271 9503
rect 25605 9469 25639 9503
rect 3433 9401 3467 9435
rect 4169 9401 4203 9435
rect 8401 9401 8435 9435
rect 12817 9401 12851 9435
rect 15945 9401 15979 9435
rect 22569 9401 22603 9435
rect 24501 9401 24535 9435
rect 5641 9333 5675 9367
rect 5825 9333 5859 9367
rect 11989 9333 12023 9367
rect 16313 9333 16347 9367
rect 17325 9333 17359 9367
rect 17509 9333 17543 9367
rect 23765 9333 23799 9367
rect 24225 9333 24259 9367
rect 2513 9129 2547 9163
rect 2973 9129 3007 9163
rect 4905 9129 4939 9163
rect 7481 9129 7515 9163
rect 12817 9129 12851 9163
rect 13553 9129 13587 9163
rect 21465 9129 21499 9163
rect 25697 9129 25731 9163
rect 1869 9061 1903 9095
rect 10149 9061 10183 9095
rect 21649 9061 21683 9095
rect 8217 8993 8251 9027
rect 8401 8993 8435 9027
rect 11069 8993 11103 9027
rect 14565 8993 14599 9027
rect 17049 8993 17083 9027
rect 17325 8993 17359 9027
rect 18061 8993 18095 9027
rect 22201 8993 22235 9027
rect 23857 8993 23891 9027
rect 24685 8993 24719 9027
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 5089 8925 5123 8959
rect 5365 8925 5399 8959
rect 6101 8925 6135 8959
rect 6368 8925 6402 8959
rect 8125 8925 8159 8959
rect 8309 8925 8343 8959
rect 9229 8925 9263 8959
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 14289 8925 14323 8959
rect 17785 8925 17819 8959
rect 20177 8925 20211 8959
rect 20361 8925 20395 8959
rect 20821 8925 20855 8959
rect 22109 8925 22143 8959
rect 23397 8925 23431 8959
rect 23489 8925 23523 8959
rect 24777 8925 24811 8959
rect 25605 8925 25639 8959
rect 25789 8925 25823 8959
rect 4353 8857 4387 8891
rect 5273 8857 5307 8891
rect 11345 8857 11379 8891
rect 13737 8857 13771 8891
rect 21281 8857 21315 8891
rect 21481 8857 21515 8891
rect 23765 8857 23799 8891
rect 3341 8789 3375 8823
rect 7941 8789 7975 8823
rect 9321 8789 9355 8823
rect 13369 8789 13403 8823
rect 13537 8789 13571 8823
rect 16037 8789 16071 8823
rect 19533 8789 19567 8823
rect 23213 8789 23247 8823
rect 25145 8789 25179 8823
rect 4077 8585 4111 8619
rect 4261 8585 4295 8619
rect 5549 8585 5583 8619
rect 5917 8585 5951 8619
rect 6653 8585 6687 8619
rect 7757 8585 7791 8619
rect 16129 8585 16163 8619
rect 17325 8585 17359 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 20729 8585 20763 8619
rect 22201 8585 22235 8619
rect 24133 8585 24167 8619
rect 25697 8585 25731 8619
rect 1961 8517 1995 8551
rect 3065 8517 3099 8551
rect 3433 8517 3467 8551
rect 4445 8517 4479 8551
rect 12341 8517 12375 8551
rect 12541 8517 12575 8551
rect 14749 8517 14783 8551
rect 15209 8517 15243 8551
rect 18613 8517 18647 8551
rect 20053 8517 20087 8551
rect 20269 8517 20303 8551
rect 23020 8517 23054 8551
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 5733 8449 5767 8483
rect 6009 8449 6043 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 7849 8449 7883 8483
rect 8769 8449 8803 8483
rect 9413 8449 9447 8483
rect 15393 8449 15427 8483
rect 15577 8449 15611 8483
rect 16313 8449 16347 8483
rect 18245 8449 18279 8483
rect 18429 8449 18463 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 20913 8449 20947 8483
rect 21097 8449 21131 8483
rect 22017 8449 22051 8483
rect 22753 8449 22787 8483
rect 25053 8449 25087 8483
rect 7573 8381 7607 8415
rect 11161 8381 11195 8415
rect 15669 8381 15703 8415
rect 17233 8381 17267 8415
rect 19073 8381 19107 8415
rect 24685 8381 24719 8415
rect 25145 8381 25179 8415
rect 2513 8313 2547 8347
rect 4997 8313 5031 8347
rect 8217 8313 8251 8347
rect 12173 8313 12207 8347
rect 13461 8313 13495 8347
rect 4261 8245 4295 8279
rect 7021 8245 7055 8279
rect 8953 8245 8987 8279
rect 9676 8245 9710 8279
rect 12357 8245 12391 8279
rect 19901 8245 19935 8279
rect 20085 8245 20119 8279
rect 2881 8041 2915 8075
rect 3985 8041 4019 8075
rect 6561 8041 6595 8075
rect 9321 8041 9355 8075
rect 10149 8041 10183 8075
rect 10793 8041 10827 8075
rect 18889 8041 18923 8075
rect 22937 8041 22971 8075
rect 24593 8041 24627 8075
rect 2053 7973 2087 8007
rect 9137 7973 9171 8007
rect 12725 7973 12759 8007
rect 20361 7973 20395 8007
rect 23489 7973 23523 8007
rect 24041 7973 24075 8007
rect 3433 7905 3467 7939
rect 7757 7905 7791 7939
rect 8217 7905 8251 7939
rect 12311 7905 12345 7939
rect 13369 7905 13403 7939
rect 14933 7905 14967 7939
rect 21097 7905 21131 7939
rect 4169 7837 4203 7871
rect 4445 7837 4479 7871
rect 5273 7837 5307 7871
rect 7849 7837 7883 7871
rect 9689 7837 9723 7871
rect 10701 7837 10735 7871
rect 10977 7837 11011 7871
rect 12173 7837 12207 7871
rect 12449 7837 12483 7871
rect 13185 7837 13219 7871
rect 14749 7837 14783 7871
rect 17417 7837 17451 7871
rect 18061 7837 18095 7871
rect 18153 7837 18187 7871
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 21925 7837 21959 7871
rect 22109 7837 22143 7871
rect 22753 7837 22787 7871
rect 22937 7837 22971 7871
rect 4353 7769 4387 7803
rect 8125 7769 8159 7803
rect 9321 7769 9355 7803
rect 17877 7769 17911 7803
rect 19441 7769 19475 7803
rect 22293 7769 22327 7803
rect 7573 7701 7607 7735
rect 7941 7701 7975 7735
rect 11529 7701 11563 7735
rect 16129 7701 16163 7735
rect 2053 7497 2087 7531
rect 3709 7497 3743 7531
rect 4261 7497 4295 7531
rect 5457 7497 5491 7531
rect 7757 7497 7791 7531
rect 8493 7497 8527 7531
rect 11161 7497 11195 7531
rect 16313 7497 16347 7531
rect 23489 7497 23523 7531
rect 5917 7429 5951 7463
rect 7389 7429 7423 7463
rect 3157 7361 3191 7395
rect 5273 7361 5307 7395
rect 6653 7361 6687 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 8309 7361 8343 7395
rect 9137 7361 9171 7395
rect 9321 7361 9355 7395
rect 10048 7361 10082 7395
rect 11713 7361 11747 7395
rect 13369 7361 13403 7395
rect 13553 7361 13587 7395
rect 19257 7361 19291 7395
rect 22201 7361 22235 7395
rect 22753 7361 22787 7395
rect 9781 7293 9815 7327
rect 12357 7293 12391 7327
rect 12495 7293 12529 7327
rect 12633 7293 12667 7327
rect 14013 7293 14047 7327
rect 14289 7293 14323 7327
rect 16865 7293 16899 7327
rect 17141 7293 17175 7327
rect 19717 7293 19751 7327
rect 21189 7293 21223 7327
rect 21465 7293 21499 7327
rect 22017 7293 22051 7327
rect 4813 7225 4847 7259
rect 9229 7225 9263 7259
rect 12909 7225 12943 7259
rect 15761 7225 15795 7259
rect 19073 7225 19107 7259
rect 22845 7225 22879 7259
rect 6837 7157 6871 7191
rect 18613 7157 18647 7191
rect 7389 6953 7423 6987
rect 7573 6953 7607 6987
rect 8401 6953 8435 6987
rect 11069 6953 11103 6987
rect 12909 6953 12943 6987
rect 16589 6885 16623 6919
rect 22385 6885 22419 6919
rect 1961 6817 1995 6851
rect 3433 6817 3467 6851
rect 4353 6817 4387 6851
rect 4997 6817 5031 6851
rect 9137 6817 9171 6851
rect 11529 6817 11563 6851
rect 13553 6817 13587 6851
rect 14289 6817 14323 6851
rect 17141 6817 17175 6851
rect 6101 6749 6135 6783
rect 6929 6749 6963 6783
rect 9689 6749 9723 6783
rect 13461 6749 13495 6783
rect 13645 6749 13679 6783
rect 16497 6749 16531 6783
rect 16681 6749 16715 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 20453 6749 20487 6783
rect 22569 6749 22603 6783
rect 5549 6681 5583 6715
rect 6837 6681 6871 6715
rect 7757 6681 7791 6715
rect 8217 6681 8251 6715
rect 9956 6681 9990 6715
rect 11774 6681 11808 6715
rect 14565 6681 14599 6715
rect 17417 6681 17451 6715
rect 2513 6613 2547 6647
rect 6193 6613 6227 6647
rect 7557 6613 7591 6647
rect 8417 6613 8451 6647
rect 8585 6613 8619 6647
rect 16037 6613 16071 6647
rect 18889 6613 18923 6647
rect 19625 6613 19659 6647
rect 21879 6613 21913 6647
rect 3341 6409 3375 6443
rect 5457 6409 5491 6443
rect 7021 6409 7055 6443
rect 9229 6409 9263 6443
rect 11161 6409 11195 6443
rect 16313 6409 16347 6443
rect 19257 6409 19291 6443
rect 21281 6409 21315 6443
rect 4353 6341 4387 6375
rect 10048 6341 10082 6375
rect 11713 6341 11747 6375
rect 13001 6341 13035 6375
rect 17877 6341 17911 6375
rect 20821 6341 20855 6375
rect 2329 6273 2363 6307
rect 3801 6273 3835 6307
rect 6929 6273 6963 6307
rect 8585 6273 8619 6307
rect 9781 6273 9815 6307
rect 11897 6273 11931 6307
rect 12081 6273 12115 6307
rect 15945 6273 15979 6307
rect 17049 6273 17083 6307
rect 18337 6273 18371 6307
rect 18521 6273 18555 6307
rect 19349 6273 19383 6307
rect 20545 6273 20579 6307
rect 20729 6273 20763 6307
rect 8401 6205 8435 6239
rect 14749 6205 14783 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 16957 6205 16991 6239
rect 17509 6205 17543 6239
rect 19073 6205 19107 6239
rect 7849 6137 7883 6171
rect 8769 6137 8803 6171
rect 1777 6069 1811 6103
rect 5917 6069 5951 6103
rect 17417 6069 17451 6103
rect 18429 6069 18463 6103
rect 19717 6069 19751 6103
rect 7849 5865 7883 5899
rect 14381 5865 14415 5899
rect 14933 5865 14967 5899
rect 17877 5865 17911 5899
rect 19441 5865 19475 5899
rect 20729 5865 20763 5899
rect 2789 5797 2823 5831
rect 4537 5797 4571 5831
rect 5089 5797 5123 5831
rect 5733 5797 5767 5831
rect 8585 5797 8619 5831
rect 10885 5797 10919 5831
rect 21373 5797 21407 5831
rect 2329 5729 2363 5763
rect 3433 5729 3467 5763
rect 4077 5729 4111 5763
rect 6285 5729 6319 5763
rect 12541 5729 12575 5763
rect 12817 5729 12851 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 19993 5729 20027 5763
rect 7297 5661 7331 5695
rect 8401 5661 8435 5695
rect 9505 5661 9539 5695
rect 12265 5661 12299 5695
rect 12424 5661 12458 5695
rect 13277 5661 13311 5695
rect 13461 5661 13495 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 18245 5661 18279 5695
rect 19809 5661 19843 5695
rect 20729 5661 20763 5695
rect 21557 5661 21591 5695
rect 6837 5593 6871 5627
rect 9772 5593 9806 5627
rect 15669 5593 15703 5627
rect 11621 5525 11655 5559
rect 16957 5525 16991 5559
rect 19901 5525 19935 5559
rect 22109 5525 22143 5559
rect 2605 5321 2639 5355
rect 3525 5321 3559 5355
rect 4077 5321 4111 5355
rect 4537 5321 4571 5355
rect 5181 5321 5215 5355
rect 5917 5321 5951 5355
rect 8217 5321 8251 5355
rect 10701 5321 10735 5355
rect 15577 5321 15611 5355
rect 17141 5321 17175 5355
rect 19441 5321 19475 5355
rect 14464 5253 14498 5287
rect 17233 5253 17267 5287
rect 18306 5253 18340 5287
rect 22201 5253 22235 5287
rect 7021 5185 7055 5219
rect 8861 5185 8895 5219
rect 9321 5185 9355 5219
rect 9588 5185 9622 5219
rect 13553 5185 13587 5219
rect 16037 5185 16071 5219
rect 19901 5185 19935 5219
rect 21097 5185 21131 5219
rect 22017 5185 22051 5219
rect 22385 5185 22419 5219
rect 23489 5185 23523 5219
rect 12357 5117 12391 5151
rect 12495 5117 12529 5151
rect 12633 5117 12667 5151
rect 12909 5117 12943 5151
rect 13369 5117 13403 5151
rect 14197 5117 14231 5151
rect 16957 5117 16991 5151
rect 18061 5117 18095 5151
rect 20177 5117 20211 5151
rect 7665 5049 7699 5083
rect 21005 5049 21039 5083
rect 8677 4981 8711 5015
rect 11713 4981 11747 5015
rect 16221 4981 16255 5015
rect 17601 4981 17635 5015
rect 19993 4981 20027 5015
rect 20453 4981 20487 5015
rect 23305 4981 23339 5015
rect 4629 4777 4663 4811
rect 5181 4777 5215 4811
rect 6653 4777 6687 4811
rect 7297 4777 7331 4811
rect 7941 4777 7975 4811
rect 10793 4777 10827 4811
rect 6101 4709 6135 4743
rect 13001 4709 13035 4743
rect 18889 4709 18923 4743
rect 19533 4709 19567 4743
rect 11253 4641 11287 4675
rect 12449 4641 12483 4675
rect 13553 4641 13587 4675
rect 17509 4641 17543 4675
rect 19717 4641 19751 4675
rect 8401 4573 8435 4607
rect 9413 4573 9447 4607
rect 14289 4573 14323 4607
rect 17765 4573 17799 4607
rect 19441 4573 19475 4607
rect 20361 4573 20395 4607
rect 21005 4573 21039 4607
rect 22845 4573 22879 4607
rect 23489 4573 23523 4607
rect 9680 4505 9714 4539
rect 13461 4505 13495 4539
rect 15209 4505 15243 4539
rect 19717 4505 19751 4539
rect 22600 4505 22634 4539
rect 8493 4437 8527 4471
rect 11805 4437 11839 4471
rect 12173 4437 12207 4471
rect 12265 4437 12299 4471
rect 13369 4437 13403 4471
rect 14473 4437 14507 4471
rect 16497 4437 16531 4471
rect 20177 4437 20211 4471
rect 20913 4437 20947 4471
rect 21465 4437 21499 4471
rect 23305 4437 23339 4471
rect 4629 4233 4663 4267
rect 17233 4233 17267 4267
rect 20453 4233 20487 4267
rect 20269 4165 20303 4199
rect 21005 4165 21039 4199
rect 22284 4165 22318 4199
rect 7757 4097 7791 4131
rect 8861 4097 8895 4131
rect 9588 4097 9622 4131
rect 11805 4097 11839 4131
rect 12705 4097 12739 4131
rect 14289 4097 14323 4131
rect 14556 4097 14590 4131
rect 16313 4097 16347 4131
rect 17325 4097 17359 4131
rect 19553 4097 19587 4131
rect 20545 4097 20579 4131
rect 22017 4097 22051 4131
rect 9321 4029 9355 4063
rect 12449 4029 12483 4063
rect 17417 4029 17451 4063
rect 19809 4029 19843 4063
rect 10701 3961 10735 3995
rect 16865 3961 16899 3995
rect 21373 3961 21407 3995
rect 23397 3961 23431 3995
rect 8677 3893 8711 3927
rect 11989 3893 12023 3927
rect 13829 3893 13863 3927
rect 15669 3893 15703 3927
rect 16129 3893 16163 3927
rect 18429 3893 18463 3927
rect 20269 3893 20303 3927
rect 21465 3893 21499 3927
rect 23949 3893 23983 3927
rect 9229 3689 9263 3723
rect 11897 3689 11931 3723
rect 15485 3689 15519 3723
rect 18521 3689 18555 3723
rect 20729 3689 20763 3723
rect 23121 3689 23155 3723
rect 23581 3689 23615 3723
rect 20177 3621 20211 3655
rect 23489 3621 23523 3655
rect 8493 3553 8527 3587
rect 10517 3553 10551 3587
rect 14841 3553 14875 3587
rect 17969 3553 18003 3587
rect 19533 3553 19567 3587
rect 22569 3553 22603 3587
rect 23397 3553 23431 3587
rect 7757 3485 7791 3519
rect 8401 3485 8435 3519
rect 9413 3485 9447 3519
rect 9873 3485 9907 3519
rect 12357 3485 12391 3519
rect 15117 3485 15151 3519
rect 15945 3485 15979 3519
rect 16212 3485 16246 3519
rect 18153 3485 18187 3519
rect 19809 3485 19843 3519
rect 22313 3485 22347 3519
rect 23949 3485 23983 3519
rect 24777 3485 24811 3519
rect 10762 3417 10796 3451
rect 12602 3417 12636 3451
rect 7941 3349 7975 3383
rect 9965 3349 9999 3383
rect 13737 3349 13771 3383
rect 15025 3349 15059 3383
rect 17325 3349 17359 3383
rect 18061 3349 18095 3383
rect 19717 3349 19751 3383
rect 21189 3349 21223 3383
rect 24593 3349 24627 3383
rect 11161 3145 11195 3179
rect 15209 3145 15243 3179
rect 15669 3145 15703 3179
rect 20177 3145 20211 3179
rect 20821 3145 20855 3179
rect 23397 3145 23431 3179
rect 25237 3145 25271 3179
rect 10037 3077 10071 3111
rect 14749 3077 14783 3111
rect 22284 3077 22318 3111
rect 1869 3009 1903 3043
rect 8493 3009 8527 3043
rect 9321 3009 9355 3043
rect 11805 3009 11839 3043
rect 12265 3009 12299 3043
rect 15577 3009 15611 3043
rect 17325 3009 17359 3043
rect 18898 3009 18932 3043
rect 19165 3009 19199 3043
rect 20361 3009 20395 3043
rect 21005 3009 21039 3043
rect 21189 3009 21223 3043
rect 21465 3009 21499 3043
rect 22017 3009 22051 3043
rect 23857 3009 23891 3043
rect 24777 3009 24811 3043
rect 8585 2941 8619 2975
rect 9781 2941 9815 2975
rect 13001 2941 13035 2975
rect 15761 2941 15795 2975
rect 28365 2941 28399 2975
rect 9137 2873 9171 2907
rect 24041 2873 24075 2907
rect 24593 2873 24627 2907
rect 1685 2805 1719 2839
rect 6561 2805 6595 2839
rect 7205 2805 7239 2839
rect 8033 2805 8067 2839
rect 12449 2805 12483 2839
rect 17141 2805 17175 2839
rect 17785 2805 17819 2839
rect 21373 2805 21407 2839
rect 8585 2601 8619 2635
rect 10333 2601 10367 2635
rect 12541 2601 12575 2635
rect 14381 2601 14415 2635
rect 16313 2601 16347 2635
rect 18337 2601 18371 2635
rect 23857 2601 23891 2635
rect 7941 2533 7975 2567
rect 20361 2533 20395 2567
rect 21373 2533 21407 2567
rect 22385 2533 22419 2567
rect 23029 2533 23063 2567
rect 24777 2533 24811 2567
rect 7297 2465 7331 2499
rect 13001 2465 13035 2499
rect 13185 2465 13219 2499
rect 14933 2465 14967 2499
rect 2053 2397 2087 2431
rect 3157 2397 3191 2431
rect 4261 2397 4295 2431
rect 5089 2397 5123 2431
rect 8401 2397 8435 2431
rect 9597 2397 9631 2431
rect 10241 2397 10275 2431
rect 11161 2397 11195 2431
rect 12081 2397 12115 2431
rect 14473 2397 14507 2431
rect 16865 2397 16899 2431
rect 17601 2397 17635 2431
rect 18521 2397 18555 2431
rect 18797 2397 18831 2431
rect 19441 2397 19475 2431
rect 20177 2397 20211 2431
rect 21005 2397 21039 2431
rect 22017 2397 22051 2431
rect 23213 2397 23247 2431
rect 23673 2397 23707 2431
rect 24593 2397 24627 2431
rect 25329 2397 25363 2431
rect 26065 2397 26099 2431
rect 27169 2397 27203 2431
rect 28181 2397 28215 2431
rect 15200 2329 15234 2363
rect 1869 2261 1903 2295
rect 2973 2261 3007 2295
rect 4077 2261 4111 2295
rect 9781 2261 9815 2295
rect 10977 2261 11011 2295
rect 11897 2261 11931 2295
rect 12909 2261 12943 2295
rect 17049 2261 17083 2295
rect 17785 2261 17819 2295
rect 18705 2261 18739 2295
rect 19625 2261 19659 2295
rect 21465 2261 21499 2295
rect 22477 2261 22511 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 3421 27591 3479 27597
rect 3421 27557 3433 27591
rect 3467 27588 3479 27591
rect 3786 27588 3792 27600
rect 3467 27560 3792 27588
rect 3467 27557 3479 27560
rect 3421 27551 3479 27557
rect 3786 27548 3792 27560
rect 3844 27548 3850 27600
rect 8570 27588 8576 27600
rect 8531 27560 8576 27588
rect 8570 27548 8576 27560
rect 8628 27548 8634 27600
rect 9309 27591 9367 27597
rect 9309 27557 9321 27591
rect 9355 27557 9367 27591
rect 9309 27551 9367 27557
rect 11885 27591 11943 27597
rect 11885 27557 11897 27591
rect 11931 27588 11943 27591
rect 17862 27588 17868 27600
rect 11931 27560 17868 27588
rect 11931 27557 11943 27560
rect 11885 27551 11943 27557
rect 3804 27452 3832 27548
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 3804 27424 3985 27452
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 6546 27452 6552 27464
rect 6507 27424 6552 27452
rect 3973 27415 4031 27421
rect 6546 27412 6552 27424
rect 6604 27452 6610 27464
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 6604 27424 7205 27452
rect 6604 27412 6610 27424
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 8588 27452 8616 27548
rect 9324 27520 9352 27551
rect 17862 27548 17868 27560
rect 17920 27548 17926 27600
rect 20809 27591 20867 27597
rect 20809 27557 20821 27591
rect 20855 27588 20867 27591
rect 21174 27588 21180 27600
rect 20855 27560 21180 27588
rect 20855 27557 20867 27560
rect 20809 27551 20867 27557
rect 21174 27548 21180 27560
rect 21232 27548 21238 27600
rect 23293 27591 23351 27597
rect 23293 27557 23305 27591
rect 23339 27588 23351 27591
rect 23658 27588 23664 27600
rect 23339 27560 23664 27588
rect 23339 27557 23351 27560
rect 23293 27551 23351 27557
rect 23658 27548 23664 27560
rect 23716 27548 23722 27600
rect 25777 27591 25835 27597
rect 25777 27557 25789 27591
rect 25823 27588 25835 27591
rect 26142 27588 26148 27600
rect 25823 27560 26148 27588
rect 25823 27557 25835 27560
rect 25777 27551 25835 27557
rect 26142 27548 26148 27560
rect 26200 27548 26206 27600
rect 17770 27520 17776 27532
rect 9324 27492 17776 27520
rect 17770 27480 17776 27492
rect 17828 27480 17834 27532
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 8588 27424 9137 27452
rect 7193 27415 7251 27421
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 10413 27455 10471 27461
rect 10413 27421 10425 27455
rect 10459 27452 10471 27455
rect 11238 27452 11244 27464
rect 10459 27424 11244 27452
rect 10459 27421 10471 27424
rect 10413 27415 10471 27421
rect 11238 27412 11244 27424
rect 11296 27452 11302 27464
rect 11701 27455 11759 27461
rect 11701 27452 11713 27455
rect 11296 27424 11713 27452
rect 11296 27412 11302 27424
rect 11701 27421 11713 27424
rect 11747 27421 11759 27455
rect 12618 27452 12624 27464
rect 12579 27424 12624 27452
rect 11701 27415 11759 27421
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 12802 27452 12808 27464
rect 12763 27424 12808 27452
rect 12802 27412 12808 27424
rect 12860 27412 12866 27464
rect 13814 27412 13820 27464
rect 13872 27452 13878 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13872 27424 14289 27452
rect 13872 27412 13878 27424
rect 14277 27421 14289 27424
rect 14323 27452 14335 27455
rect 14921 27455 14979 27461
rect 14921 27452 14933 27455
rect 14323 27424 14933 27452
rect 14323 27421 14335 27424
rect 14277 27415 14335 27421
rect 14921 27421 14933 27424
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 16206 27412 16212 27464
rect 16264 27452 16270 27464
rect 17037 27455 17095 27461
rect 17037 27452 17049 27455
rect 16264 27424 17049 27452
rect 16264 27412 16270 27424
rect 17037 27421 17049 27424
rect 17083 27452 17095 27455
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 17083 27424 17509 27452
rect 17083 27421 17095 27424
rect 17037 27415 17095 27421
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 18690 27412 18696 27464
rect 18748 27452 18754 27464
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 18748 27424 19625 27452
rect 18748 27412 18754 27424
rect 19613 27421 19625 27424
rect 19659 27452 19671 27455
rect 20073 27455 20131 27461
rect 20073 27452 20085 27455
rect 19659 27424 20085 27452
rect 19659 27421 19671 27424
rect 19613 27415 19671 27421
rect 20073 27421 20085 27424
rect 20119 27421 20131 27455
rect 21192 27452 21220 27548
rect 21453 27455 21511 27461
rect 21453 27452 21465 27455
rect 21192 27424 21465 27452
rect 20073 27415 20131 27421
rect 21453 27421 21465 27424
rect 21499 27421 21511 27455
rect 23676 27452 23704 27548
rect 23937 27455 23995 27461
rect 23937 27452 23949 27455
rect 23676 27424 23949 27452
rect 21453 27415 21511 27421
rect 23937 27421 23949 27424
rect 23983 27421 23995 27455
rect 26160 27452 26188 27548
rect 26421 27455 26479 27461
rect 26421 27452 26433 27455
rect 26160 27424 26433 27452
rect 23937 27415 23995 27421
rect 26421 27421 26433 27424
rect 26467 27421 26479 27455
rect 26421 27415 26479 27421
rect 27709 27455 27767 27461
rect 27709 27421 27721 27455
rect 27755 27452 27767 27455
rect 28350 27452 28356 27464
rect 27755 27424 28356 27452
rect 27755 27421 27767 27424
rect 27709 27415 27767 27421
rect 28350 27412 28356 27424
rect 28408 27412 28414 27464
rect 13265 27387 13323 27393
rect 13265 27384 13277 27387
rect 10152 27356 13277 27384
rect 10152 27328 10180 27356
rect 13265 27353 13277 27356
rect 13311 27353 13323 27387
rect 13265 27347 13323 27353
rect 17954 27344 17960 27396
rect 18012 27384 18018 27396
rect 18012 27356 21312 27384
rect 18012 27344 18018 27356
rect 4154 27316 4160 27328
rect 4115 27288 4160 27316
rect 4154 27276 4160 27288
rect 4212 27276 4218 27328
rect 6730 27316 6736 27328
rect 6691 27288 6736 27316
rect 6730 27276 6736 27288
rect 6788 27276 6794 27328
rect 9861 27319 9919 27325
rect 9861 27285 9873 27319
rect 9907 27316 9919 27319
rect 10134 27316 10140 27328
rect 9907 27288 10140 27316
rect 9907 27285 9919 27288
rect 9861 27279 9919 27285
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 10870 27316 10876 27328
rect 10831 27288 10876 27316
rect 10870 27276 10876 27288
rect 10928 27276 10934 27328
rect 12805 27319 12863 27325
rect 12805 27285 12817 27319
rect 12851 27316 12863 27319
rect 12986 27316 12992 27328
rect 12851 27288 12992 27316
rect 12851 27285 12863 27288
rect 12805 27279 12863 27285
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 14461 27319 14519 27325
rect 14461 27285 14473 27319
rect 14507 27316 14519 27319
rect 15194 27316 15200 27328
rect 14507 27288 15200 27316
rect 14507 27285 14519 27288
rect 14461 27279 14519 27285
rect 15194 27276 15200 27288
rect 15252 27276 15258 27328
rect 15286 27276 15292 27328
rect 15344 27316 15350 27328
rect 16853 27319 16911 27325
rect 16853 27316 16865 27319
rect 15344 27288 16865 27316
rect 15344 27276 15350 27288
rect 16853 27285 16865 27288
rect 16899 27285 16911 27319
rect 16853 27279 16911 27285
rect 17678 27276 17684 27328
rect 17736 27316 17742 27328
rect 21284 27325 21312 27356
rect 19429 27319 19487 27325
rect 19429 27316 19441 27319
rect 17736 27288 19441 27316
rect 17736 27276 17742 27288
rect 19429 27285 19441 27288
rect 19475 27285 19487 27319
rect 19429 27279 19487 27285
rect 21269 27319 21327 27325
rect 21269 27285 21281 27319
rect 21315 27285 21327 27319
rect 23750 27316 23756 27328
rect 23711 27288 23756 27316
rect 21269 27279 21327 27285
rect 23750 27276 23756 27288
rect 23808 27276 23814 27328
rect 26234 27316 26240 27328
rect 26195 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 28166 27316 28172 27328
rect 28127 27288 28172 27316
rect 28166 27276 28172 27288
rect 28224 27276 28230 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 8849 27115 8907 27121
rect 8849 27081 8861 27115
rect 8895 27112 8907 27115
rect 9858 27112 9864 27124
rect 8895 27084 9864 27112
rect 8895 27081 8907 27084
rect 8849 27075 8907 27081
rect 9858 27072 9864 27084
rect 9916 27112 9922 27124
rect 10870 27112 10876 27124
rect 9916 27084 10876 27112
rect 9916 27072 9922 27084
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 9493 27047 9551 27053
rect 9493 27044 9505 27047
rect 8996 27016 9505 27044
rect 8996 27004 9002 27016
rect 9493 27013 9505 27016
rect 9539 27013 9551 27047
rect 9493 27007 9551 27013
rect 12253 27047 12311 27053
rect 12253 27013 12265 27047
rect 12299 27044 12311 27047
rect 12710 27044 12716 27056
rect 12299 27016 12716 27044
rect 12299 27013 12311 27016
rect 12253 27007 12311 27013
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 12894 27004 12900 27056
rect 12952 27044 12958 27056
rect 13909 27047 13967 27053
rect 13909 27044 13921 27047
rect 12952 27016 13921 27044
rect 12952 27004 12958 27016
rect 13909 27013 13921 27016
rect 13955 27044 13967 27047
rect 13998 27044 14004 27056
rect 13955 27016 14004 27044
rect 13955 27013 13967 27016
rect 13909 27007 13967 27013
rect 13998 27004 14004 27016
rect 14056 27004 14062 27056
rect 8386 26936 8392 26988
rect 8444 26976 8450 26988
rect 9309 26979 9367 26985
rect 9309 26976 9321 26979
rect 8444 26948 9321 26976
rect 8444 26936 8450 26948
rect 9309 26945 9321 26948
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 9585 26979 9643 26985
rect 9585 26945 9597 26979
rect 9631 26945 9643 26979
rect 9585 26939 9643 26945
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 9600 26908 9628 26939
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10744 26948 10793 26976
rect 10744 26936 10750 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10962 26976 10968 26988
rect 10923 26948 10968 26976
rect 10781 26939 10839 26945
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 11790 26936 11796 26988
rect 11848 26976 11854 26988
rect 12069 26979 12127 26985
rect 12069 26976 12081 26979
rect 11848 26948 12081 26976
rect 11848 26936 11854 26948
rect 12069 26945 12081 26948
rect 12115 26945 12127 26979
rect 12345 26979 12403 26985
rect 12345 26976 12357 26979
rect 12069 26939 12127 26945
rect 12268 26948 12357 26976
rect 12268 26920 12296 26948
rect 12345 26945 12357 26948
rect 12391 26976 12403 26979
rect 12802 26976 12808 26988
rect 12391 26948 12808 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 12986 26976 12992 26988
rect 12947 26948 12992 26976
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 13814 26976 13820 26988
rect 13775 26948 13820 26976
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 9456 26880 9628 26908
rect 9456 26868 9462 26880
rect 12250 26868 12256 26920
rect 12308 26868 12314 26920
rect 13081 26911 13139 26917
rect 13081 26877 13093 26911
rect 13127 26908 13139 26911
rect 13170 26908 13176 26920
rect 13127 26880 13176 26908
rect 13127 26877 13139 26880
rect 13081 26871 13139 26877
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 6730 26800 6736 26852
rect 6788 26840 6794 26852
rect 12069 26843 12127 26849
rect 6788 26812 11284 26840
rect 6788 26800 6794 26812
rect 9309 26775 9367 26781
rect 9309 26741 9321 26775
rect 9355 26772 9367 26775
rect 9950 26772 9956 26784
rect 9355 26744 9956 26772
rect 9355 26741 9367 26744
rect 9309 26735 9367 26741
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 10042 26732 10048 26784
rect 10100 26772 10106 26784
rect 10965 26775 11023 26781
rect 10100 26744 10145 26772
rect 10100 26732 10106 26744
rect 10965 26741 10977 26775
rect 11011 26772 11023 26775
rect 11146 26772 11152 26784
rect 11011 26744 11152 26772
rect 11011 26741 11023 26744
rect 10965 26735 11023 26741
rect 11146 26732 11152 26744
rect 11204 26732 11210 26784
rect 11256 26772 11284 26812
rect 12069 26809 12081 26843
rect 12115 26840 12127 26843
rect 12342 26840 12348 26852
rect 12115 26812 12348 26840
rect 12115 26809 12127 26812
rect 12069 26803 12127 26809
rect 12342 26800 12348 26812
rect 12400 26840 12406 26852
rect 14108 26840 14136 26939
rect 12400 26812 14136 26840
rect 12400 26800 12406 26812
rect 13078 26772 13084 26784
rect 11256 26744 13084 26772
rect 13078 26732 13084 26744
rect 13136 26732 13142 26784
rect 13265 26775 13323 26781
rect 13265 26741 13277 26775
rect 13311 26772 13323 26775
rect 13630 26772 13636 26784
rect 13311 26744 13636 26772
rect 13311 26741 13323 26744
rect 13265 26735 13323 26741
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 14093 26775 14151 26781
rect 14093 26741 14105 26775
rect 14139 26772 14151 26775
rect 14274 26772 14280 26784
rect 14139 26744 14280 26772
rect 14139 26741 14151 26744
rect 14093 26735 14151 26741
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 15841 26775 15899 26781
rect 15841 26741 15853 26775
rect 15887 26772 15899 26775
rect 17034 26772 17040 26784
rect 15887 26744 17040 26772
rect 15887 26741 15899 26744
rect 15841 26735 15899 26741
rect 17034 26732 17040 26744
rect 17092 26732 17098 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 10597 26571 10655 26577
rect 10597 26537 10609 26571
rect 10643 26568 10655 26571
rect 10686 26568 10692 26580
rect 10643 26540 10692 26568
rect 10643 26537 10655 26540
rect 10597 26531 10655 26537
rect 10686 26528 10692 26540
rect 10744 26528 10750 26580
rect 11146 26568 11152 26580
rect 11107 26540 11152 26568
rect 11146 26528 11152 26540
rect 11204 26528 11210 26580
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12894 26568 12900 26580
rect 12391 26540 12900 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 13262 26528 13268 26580
rect 13320 26568 13326 26580
rect 17034 26568 17040 26580
rect 13320 26540 14320 26568
rect 13320 26528 13326 26540
rect 12250 26500 12256 26512
rect 11440 26472 12256 26500
rect 10428 26404 11100 26432
rect 8386 26364 8392 26376
rect 8347 26336 8392 26364
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 8570 26364 8576 26376
rect 8531 26336 8576 26364
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 9364 26336 9413 26364
rect 9364 26324 9370 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 9401 26327 9459 26333
rect 9585 26367 9643 26373
rect 9585 26333 9597 26367
rect 9631 26333 9643 26367
rect 9585 26327 9643 26333
rect 4062 26296 4068 26308
rect 4023 26268 4068 26296
rect 4062 26256 4068 26268
rect 4120 26256 4126 26308
rect 8478 26296 8484 26308
rect 8391 26268 8484 26296
rect 8478 26256 8484 26268
rect 8536 26296 8542 26308
rect 9600 26296 9628 26327
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10428 26373 10456 26404
rect 10413 26367 10471 26373
rect 10413 26364 10425 26367
rect 10008 26336 10425 26364
rect 10008 26324 10014 26336
rect 10413 26333 10425 26336
rect 10459 26333 10471 26367
rect 10413 26327 10471 26333
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 10962 26364 10968 26376
rect 10652 26336 10968 26364
rect 10652 26324 10658 26336
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 11072 26373 11100 26404
rect 11057 26367 11115 26373
rect 11057 26333 11069 26367
rect 11103 26333 11115 26367
rect 11057 26327 11115 26333
rect 11440 26296 11468 26472
rect 12250 26460 12256 26472
rect 12308 26500 12314 26512
rect 12308 26472 13032 26500
rect 12308 26460 12314 26472
rect 11517 26435 11575 26441
rect 11517 26401 11529 26435
rect 11563 26432 11575 26435
rect 12618 26432 12624 26444
rect 11563 26404 12624 26432
rect 11563 26401 11575 26404
rect 11517 26395 11575 26401
rect 12618 26392 12624 26404
rect 12676 26432 12682 26444
rect 13004 26441 13032 26472
rect 13078 26460 13084 26512
rect 13136 26500 13142 26512
rect 13136 26472 14044 26500
rect 13136 26460 13142 26472
rect 12989 26435 13047 26441
rect 12676 26404 12756 26432
rect 12676 26392 12682 26404
rect 11790 26324 11796 26376
rect 11848 26364 11854 26376
rect 12069 26367 12127 26373
rect 12069 26364 12081 26367
rect 11848 26336 12081 26364
rect 11848 26324 11854 26336
rect 12069 26333 12081 26336
rect 12115 26333 12127 26367
rect 12342 26364 12348 26376
rect 12303 26336 12348 26364
rect 12069 26327 12127 26333
rect 12342 26324 12348 26336
rect 12400 26324 12406 26376
rect 12161 26299 12219 26305
rect 12161 26296 12173 26299
rect 8536 26268 9628 26296
rect 10244 26268 12173 26296
rect 8536 26256 8542 26268
rect 2130 26228 2136 26240
rect 2091 26200 2136 26228
rect 2130 26188 2136 26200
rect 2188 26188 2194 26240
rect 2590 26228 2596 26240
rect 2551 26200 2596 26228
rect 2590 26188 2596 26200
rect 2648 26188 2654 26240
rect 3142 26188 3148 26240
rect 3200 26228 3206 26240
rect 3329 26231 3387 26237
rect 3329 26228 3341 26231
rect 3200 26200 3341 26228
rect 3200 26188 3206 26200
rect 3329 26197 3341 26200
rect 3375 26197 3387 26231
rect 3329 26191 3387 26197
rect 5353 26231 5411 26237
rect 5353 26197 5365 26231
rect 5399 26228 5411 26231
rect 6454 26228 6460 26240
rect 5399 26200 6460 26228
rect 5399 26197 5411 26200
rect 5353 26191 5411 26197
rect 6454 26188 6460 26200
rect 6512 26188 6518 26240
rect 7929 26231 7987 26237
rect 7929 26197 7941 26231
rect 7975 26228 7987 26231
rect 8294 26228 8300 26240
rect 7975 26200 8300 26228
rect 7975 26197 7987 26200
rect 7929 26191 7987 26197
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 9766 26228 9772 26240
rect 9727 26200 9772 26228
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 10244 26237 10272 26268
rect 12161 26265 12173 26268
rect 12207 26265 12219 26299
rect 12728 26296 12756 26404
rect 12989 26401 13001 26435
rect 13035 26401 13047 26435
rect 12989 26395 13047 26401
rect 13357 26435 13415 26441
rect 13357 26401 13369 26435
rect 13403 26432 13415 26435
rect 13906 26432 13912 26444
rect 13403 26404 13912 26432
rect 13403 26401 13415 26404
rect 13357 26395 13415 26401
rect 13906 26392 13912 26404
rect 13964 26392 13970 26444
rect 12894 26364 12900 26376
rect 12855 26336 12900 26364
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13096 26296 13124 26327
rect 13170 26324 13176 26376
rect 13228 26364 13234 26376
rect 13228 26336 13273 26364
rect 13228 26324 13234 26336
rect 12728 26268 13124 26296
rect 14016 26296 14044 26472
rect 14292 26373 14320 26540
rect 16776 26540 17040 26568
rect 16776 26500 16804 26540
rect 17034 26528 17040 26540
rect 17092 26568 17098 26580
rect 17092 26540 18092 26568
rect 17092 26528 17098 26540
rect 15120 26472 16804 26500
rect 15120 26441 15148 26472
rect 15105 26435 15163 26441
rect 15105 26401 15117 26435
rect 15151 26401 15163 26435
rect 15105 26395 15163 26401
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 16776 26441 16804 26472
rect 18064 26444 18092 26540
rect 23750 26500 23756 26512
rect 18524 26472 23756 26500
rect 16577 26435 16635 26441
rect 16577 26432 16589 26435
rect 15252 26404 16589 26432
rect 15252 26392 15258 26404
rect 16577 26401 16589 26404
rect 16623 26401 16635 26435
rect 16577 26395 16635 26401
rect 16761 26435 16819 26441
rect 16761 26401 16773 26435
rect 16807 26401 16819 26435
rect 17770 26432 17776 26444
rect 17731 26404 17776 26432
rect 16761 26395 16819 26401
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26432 18015 26435
rect 18046 26432 18052 26444
rect 18003 26404 18052 26432
rect 18003 26401 18015 26404
rect 17957 26395 18015 26401
rect 18046 26392 18052 26404
rect 18104 26392 18110 26444
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14458 26364 14464 26376
rect 14419 26336 14464 26364
rect 14277 26327 14335 26333
rect 14458 26324 14464 26336
rect 14516 26324 14522 26376
rect 15286 26364 15292 26376
rect 15247 26336 15292 26364
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26333 16543 26367
rect 17678 26364 17684 26376
rect 17639 26336 17684 26364
rect 16485 26327 16543 26333
rect 15197 26299 15255 26305
rect 15197 26296 15209 26299
rect 14016 26268 15209 26296
rect 12161 26259 12219 26265
rect 15197 26265 15209 26268
rect 15243 26265 15255 26299
rect 16500 26296 16528 26327
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 18524 26296 18552 26472
rect 23750 26460 23756 26472
rect 23808 26460 23814 26512
rect 28166 26432 28172 26444
rect 22066 26404 28172 26432
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26364 19671 26367
rect 22066 26364 22094 26404
rect 28166 26392 28172 26404
rect 28224 26392 28230 26444
rect 19659 26336 22094 26364
rect 25409 26367 25467 26373
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 25409 26333 25421 26367
rect 25455 26364 25467 26367
rect 26234 26364 26240 26376
rect 25455 26336 26240 26364
rect 25455 26333 25467 26336
rect 25409 26327 25467 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 19518 26296 19524 26308
rect 16500 26268 18552 26296
rect 19479 26268 19524 26296
rect 15197 26259 15255 26265
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 24946 26256 24952 26308
rect 25004 26296 25010 26308
rect 25317 26299 25375 26305
rect 25317 26296 25329 26299
rect 25004 26268 25329 26296
rect 25004 26256 25010 26268
rect 25317 26265 25329 26268
rect 25363 26265 25375 26299
rect 25317 26259 25375 26265
rect 10229 26231 10287 26237
rect 10229 26197 10241 26231
rect 10275 26197 10287 26231
rect 14366 26228 14372 26240
rect 14327 26200 14372 26228
rect 10229 26191 10287 26197
rect 14366 26188 14372 26200
rect 14424 26188 14430 26240
rect 15654 26228 15660 26240
rect 15615 26200 15660 26228
rect 15654 26188 15660 26200
rect 15712 26188 15718 26240
rect 16117 26231 16175 26237
rect 16117 26197 16129 26231
rect 16163 26228 16175 26231
rect 16206 26228 16212 26240
rect 16163 26200 16212 26228
rect 16163 26197 16175 26200
rect 16117 26191 16175 26197
rect 16206 26188 16212 26200
rect 16264 26188 16270 26240
rect 17126 26188 17132 26240
rect 17184 26228 17190 26240
rect 17313 26231 17371 26237
rect 17313 26228 17325 26231
rect 17184 26200 17325 26228
rect 17184 26188 17190 26200
rect 17313 26197 17325 26200
rect 17359 26197 17371 26231
rect 17313 26191 17371 26197
rect 18601 26231 18659 26237
rect 18601 26197 18613 26231
rect 18647 26228 18659 26231
rect 18690 26228 18696 26240
rect 18647 26200 18696 26228
rect 18647 26197 18659 26200
rect 18601 26191 18659 26197
rect 18690 26188 18696 26200
rect 18748 26188 18754 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 4062 26024 4068 26036
rect 2746 25996 4068 26024
rect 2222 25848 2228 25900
rect 2280 25888 2286 25900
rect 2746 25888 2774 25996
rect 4062 25984 4068 25996
rect 4120 26024 4126 26036
rect 4893 26027 4951 26033
rect 4893 26024 4905 26027
rect 4120 25996 4905 26024
rect 4120 25984 4126 25996
rect 4893 25993 4905 25996
rect 4939 25993 4951 26027
rect 10594 26024 10600 26036
rect 10555 25996 10600 26024
rect 4893 25987 4951 25993
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 10870 26024 10876 26036
rect 10831 25996 10876 26024
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 10965 26027 11023 26033
rect 10965 25993 10977 26027
rect 11011 26024 11023 26027
rect 11054 26024 11060 26036
rect 11011 25996 11060 26024
rect 11011 25993 11023 25996
rect 10965 25987 11023 25993
rect 11054 25984 11060 25996
rect 11112 25984 11118 26036
rect 12529 26027 12587 26033
rect 12529 25993 12541 26027
rect 12575 26024 12587 26027
rect 13170 26024 13176 26036
rect 12575 25996 13176 26024
rect 12575 25993 12587 25996
rect 12529 25987 12587 25993
rect 13170 25984 13176 25996
rect 13228 25984 13234 26036
rect 13446 26024 13452 26036
rect 13359 25996 13452 26024
rect 9306 25956 9312 25968
rect 8220 25928 9312 25956
rect 8220 25897 8248 25928
rect 9306 25916 9312 25928
rect 9364 25916 9370 25968
rect 10137 25959 10195 25965
rect 10137 25925 10149 25959
rect 10183 25956 10195 25959
rect 13081 25959 13139 25965
rect 13081 25956 13093 25959
rect 10183 25928 13093 25956
rect 10183 25925 10195 25928
rect 10137 25919 10195 25925
rect 13081 25925 13093 25928
rect 13127 25956 13139 25959
rect 13372 25956 13400 25996
rect 13446 25984 13452 25996
rect 13504 26024 13510 26036
rect 14458 26024 14464 26036
rect 13504 25996 14464 26024
rect 13504 25984 13510 25996
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 17773 26027 17831 26033
rect 17773 25993 17785 26027
rect 17819 26024 17831 26027
rect 17954 26024 17960 26036
rect 17819 25996 17960 26024
rect 17819 25993 17831 25996
rect 17773 25987 17831 25993
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 13127 25928 13400 25956
rect 13127 25925 13139 25928
rect 13081 25919 13139 25925
rect 14366 25916 14372 25968
rect 14424 25956 14430 25968
rect 14645 25959 14703 25965
rect 14645 25956 14657 25959
rect 14424 25928 14657 25956
rect 14424 25916 14430 25928
rect 14645 25925 14657 25928
rect 14691 25925 14703 25959
rect 17862 25956 17868 25968
rect 17823 25928 17868 25956
rect 14645 25919 14703 25925
rect 17862 25916 17868 25928
rect 17920 25916 17926 25968
rect 2280 25860 2774 25888
rect 8205 25891 8263 25897
rect 2280 25848 2286 25860
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25888 8447 25891
rect 8478 25888 8484 25900
rect 8435 25860 8484 25888
rect 8435 25857 8447 25860
rect 8389 25851 8447 25857
rect 8478 25848 8484 25860
rect 8536 25848 8542 25900
rect 8938 25888 8944 25900
rect 8899 25860 8944 25888
rect 8938 25848 8944 25860
rect 8996 25848 9002 25900
rect 9033 25891 9091 25897
rect 9033 25857 9045 25891
rect 9079 25888 9091 25891
rect 9122 25888 9128 25900
rect 9079 25860 9128 25888
rect 9079 25857 9091 25860
rect 9033 25851 9091 25857
rect 9122 25848 9128 25860
rect 9180 25848 9186 25900
rect 9950 25888 9956 25900
rect 9911 25860 9956 25888
rect 9950 25848 9956 25860
rect 10008 25848 10014 25900
rect 10778 25888 10784 25900
rect 10739 25860 10784 25888
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 10980 25860 11713 25888
rect 2501 25823 2559 25829
rect 2501 25789 2513 25823
rect 2547 25820 2559 25823
rect 2590 25820 2596 25832
rect 2547 25792 2596 25820
rect 2547 25789 2559 25792
rect 2501 25783 2559 25789
rect 2590 25780 2596 25792
rect 2648 25820 2654 25832
rect 6914 25820 6920 25832
rect 2648 25792 6920 25820
rect 2648 25780 2654 25792
rect 6914 25780 6920 25792
rect 6972 25820 6978 25832
rect 7101 25823 7159 25829
rect 7101 25820 7113 25823
rect 6972 25792 7113 25820
rect 6972 25780 6978 25792
rect 7101 25789 7113 25792
rect 7147 25789 7159 25823
rect 7101 25783 7159 25789
rect 9217 25823 9275 25829
rect 9217 25789 9229 25823
rect 9263 25820 9275 25823
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 9263 25792 9689 25820
rect 9263 25789 9275 25792
rect 9217 25783 9275 25789
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 1949 25755 2007 25761
rect 1949 25721 1961 25755
rect 1995 25752 2007 25755
rect 2682 25752 2688 25764
rect 1995 25724 2688 25752
rect 1995 25721 2007 25724
rect 1949 25715 2007 25721
rect 2682 25712 2688 25724
rect 2740 25712 2746 25764
rect 8389 25755 8447 25761
rect 8389 25721 8401 25755
rect 8435 25752 8447 25755
rect 10980 25752 11008 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11885 25891 11943 25897
rect 11885 25857 11897 25891
rect 11931 25857 11943 25891
rect 12802 25888 12808 25900
rect 12763 25860 12808 25888
rect 11885 25851 11943 25857
rect 11146 25752 11152 25764
rect 8435 25724 11008 25752
rect 11107 25724 11152 25752
rect 8435 25721 8447 25724
rect 8389 25715 8447 25721
rect 11146 25712 11152 25724
rect 11204 25712 11210 25764
rect 3421 25687 3479 25693
rect 3421 25653 3433 25687
rect 3467 25684 3479 25687
rect 3694 25684 3700 25696
rect 3467 25656 3700 25684
rect 3467 25653 3479 25656
rect 3421 25647 3479 25653
rect 3694 25644 3700 25656
rect 3752 25684 3758 25696
rect 3881 25687 3939 25693
rect 3881 25684 3893 25687
rect 3752 25656 3893 25684
rect 3752 25644 3758 25656
rect 3881 25653 3893 25656
rect 3927 25653 3939 25687
rect 3881 25647 3939 25653
rect 5537 25687 5595 25693
rect 5537 25653 5549 25687
rect 5583 25684 5595 25687
rect 5810 25684 5816 25696
rect 5583 25656 5816 25684
rect 5583 25653 5595 25656
rect 5537 25647 5595 25653
rect 5810 25644 5816 25656
rect 5868 25644 5874 25696
rect 7650 25684 7656 25696
rect 7611 25656 7656 25684
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 9766 25684 9772 25696
rect 9679 25656 9772 25684
rect 9766 25644 9772 25656
rect 9824 25684 9830 25696
rect 11900 25684 11928 25851
rect 12802 25848 12808 25860
rect 12860 25848 12866 25900
rect 13173 25891 13231 25897
rect 13173 25857 13185 25891
rect 13219 25888 13231 25891
rect 13262 25888 13268 25900
rect 13219 25860 13268 25888
rect 13219 25857 13231 25860
rect 13173 25851 13231 25857
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13998 25888 14004 25900
rect 13959 25860 14004 25888
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14829 25891 14887 25897
rect 14829 25888 14841 25891
rect 14148 25860 14841 25888
rect 14148 25848 14154 25860
rect 14829 25857 14841 25860
rect 14875 25857 14887 25891
rect 16206 25888 16212 25900
rect 16167 25860 16212 25888
rect 14829 25851 14887 25857
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 12710 25820 12716 25832
rect 12671 25792 12716 25820
rect 12710 25780 12716 25792
rect 12768 25780 12774 25832
rect 13906 25820 13912 25832
rect 13867 25792 13912 25820
rect 13906 25780 13912 25792
rect 13964 25780 13970 25832
rect 18046 25820 18052 25832
rect 17959 25792 18052 25820
rect 18046 25780 18052 25792
rect 18104 25820 18110 25832
rect 18690 25820 18696 25832
rect 18104 25792 18696 25820
rect 18104 25780 18110 25792
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 13170 25712 13176 25764
rect 13228 25752 13234 25764
rect 13633 25755 13691 25761
rect 13633 25752 13645 25755
rect 13228 25724 13645 25752
rect 13228 25712 13234 25724
rect 13633 25721 13645 25724
rect 13679 25721 13691 25755
rect 13633 25715 13691 25721
rect 15565 25755 15623 25761
rect 15565 25721 15577 25755
rect 15611 25752 15623 25755
rect 16850 25752 16856 25764
rect 15611 25724 16856 25752
rect 15611 25721 15623 25724
rect 15565 25715 15623 25721
rect 16850 25712 16856 25724
rect 16908 25712 16914 25764
rect 12066 25684 12072 25696
rect 9824 25656 11928 25684
rect 12027 25656 12072 25684
rect 9824 25644 9830 25656
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 13354 25644 13360 25696
rect 13412 25684 13418 25696
rect 15013 25687 15071 25693
rect 15013 25684 15025 25687
rect 13412 25656 15025 25684
rect 13412 25644 13418 25656
rect 15013 25653 15025 25656
rect 15059 25653 15071 25687
rect 15013 25647 15071 25653
rect 15746 25644 15752 25696
rect 15804 25684 15810 25696
rect 16025 25687 16083 25693
rect 16025 25684 16037 25687
rect 15804 25656 16037 25684
rect 15804 25644 15810 25656
rect 16025 25653 16037 25656
rect 16071 25653 16083 25687
rect 16025 25647 16083 25653
rect 16945 25687 17003 25693
rect 16945 25653 16957 25687
rect 16991 25684 17003 25687
rect 17218 25684 17224 25696
rect 16991 25656 17224 25684
rect 16991 25653 17003 25656
rect 16945 25647 17003 25653
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 17405 25687 17463 25693
rect 17405 25653 17417 25687
rect 17451 25684 17463 25687
rect 17586 25684 17592 25696
rect 17451 25656 17592 25684
rect 17451 25653 17463 25656
rect 17405 25647 17463 25653
rect 17586 25644 17592 25656
rect 17644 25644 17650 25696
rect 18690 25684 18696 25696
rect 18651 25656 18696 25684
rect 18690 25644 18696 25656
rect 18748 25644 18754 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25449 8447 25483
rect 8389 25443 8447 25449
rect 8404 25412 8432 25443
rect 8478 25440 8484 25492
rect 8536 25480 8542 25492
rect 8573 25483 8631 25489
rect 8573 25480 8585 25483
rect 8536 25452 8585 25480
rect 8536 25440 8542 25452
rect 8573 25449 8585 25452
rect 8619 25449 8631 25483
rect 10042 25480 10048 25492
rect 8573 25443 8631 25449
rect 9646 25452 10048 25480
rect 8938 25412 8944 25424
rect 8404 25384 8944 25412
rect 8938 25372 8944 25384
rect 8996 25372 9002 25424
rect 9646 25412 9674 25452
rect 10042 25440 10048 25452
rect 10100 25440 10106 25492
rect 11790 25480 11796 25492
rect 11751 25452 11796 25480
rect 11790 25440 11796 25452
rect 11848 25440 11854 25492
rect 12894 25440 12900 25492
rect 12952 25480 12958 25492
rect 13357 25483 13415 25489
rect 13357 25480 13369 25483
rect 12952 25452 13369 25480
rect 12952 25440 12958 25452
rect 13357 25449 13369 25452
rect 13403 25449 13415 25483
rect 13357 25443 13415 25449
rect 10870 25412 10876 25424
rect 9048 25384 9674 25412
rect 10520 25384 10876 25412
rect 5718 25304 5724 25356
rect 5776 25344 5782 25356
rect 5813 25347 5871 25353
rect 5813 25344 5825 25347
rect 5776 25316 5825 25344
rect 5776 25304 5782 25316
rect 5813 25313 5825 25316
rect 5859 25344 5871 25347
rect 7193 25347 7251 25353
rect 7193 25344 7205 25347
rect 5859 25316 7205 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 7193 25313 7205 25316
rect 7239 25344 7251 25347
rect 9048 25344 9076 25384
rect 7239 25316 9076 25344
rect 7239 25313 7251 25316
rect 7193 25307 7251 25313
rect 9398 25304 9404 25356
rect 9456 25344 9462 25356
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 9456 25316 9965 25344
rect 9456 25304 9462 25316
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 9953 25307 10011 25313
rect 3053 25279 3111 25285
rect 3053 25245 3065 25279
rect 3099 25276 3111 25279
rect 3970 25276 3976 25288
rect 3099 25248 3976 25276
rect 3099 25245 3111 25248
rect 3053 25239 3111 25245
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 7745 25279 7803 25285
rect 7745 25245 7757 25279
rect 7791 25276 7803 25279
rect 8662 25276 8668 25288
rect 7791 25248 8668 25276
rect 7791 25245 7803 25248
rect 7745 25239 7803 25245
rect 8662 25236 8668 25248
rect 8720 25236 8726 25288
rect 9214 25236 9220 25288
rect 9272 25276 9278 25288
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 9272 25248 9321 25276
rect 9272 25236 9278 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25276 9551 25279
rect 9674 25276 9680 25288
rect 9539 25248 9680 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 9674 25236 9680 25248
rect 9732 25276 9738 25288
rect 10410 25276 10416 25288
rect 9732 25248 10416 25276
rect 9732 25236 9738 25248
rect 10410 25236 10416 25248
rect 10468 25236 10474 25288
rect 10520 25276 10548 25384
rect 10870 25372 10876 25384
rect 10928 25372 10934 25424
rect 10686 25344 10692 25356
rect 10647 25316 10692 25344
rect 10686 25304 10692 25316
rect 10744 25304 10750 25356
rect 10576 25279 10634 25285
rect 10576 25276 10588 25279
rect 10520 25248 10588 25276
rect 2501 25211 2559 25217
rect 2501 25177 2513 25211
rect 2547 25208 2559 25211
rect 8205 25211 8263 25217
rect 2547 25180 3740 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 3712 25152 3740 25180
rect 8205 25177 8217 25211
rect 8251 25177 8263 25211
rect 8205 25171 8263 25177
rect 8421 25211 8479 25217
rect 8421 25177 8433 25211
rect 8467 25208 8479 25211
rect 9030 25208 9036 25220
rect 8467 25180 9036 25208
rect 8467 25177 8479 25180
rect 8421 25171 8479 25177
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2222 25140 2228 25152
rect 1995 25112 2228 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 2222 25100 2228 25112
rect 2280 25100 2286 25152
rect 3694 25100 3700 25152
rect 3752 25140 3758 25152
rect 3973 25143 4031 25149
rect 3973 25140 3985 25143
rect 3752 25112 3985 25140
rect 3752 25100 3758 25112
rect 3973 25109 3985 25112
rect 4019 25109 4031 25143
rect 3973 25103 4031 25109
rect 4617 25143 4675 25149
rect 4617 25109 4629 25143
rect 4663 25140 4675 25143
rect 4706 25140 4712 25152
rect 4663 25112 4712 25140
rect 4663 25109 4675 25112
rect 4617 25103 4675 25109
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 5074 25140 5080 25152
rect 5035 25112 5080 25140
rect 5074 25100 5080 25112
rect 5132 25100 5138 25152
rect 6454 25100 6460 25152
rect 6512 25140 6518 25152
rect 6549 25143 6607 25149
rect 6549 25140 6561 25143
rect 6512 25112 6561 25140
rect 6512 25100 6518 25112
rect 6549 25109 6561 25112
rect 6595 25109 6607 25143
rect 8220 25140 8248 25171
rect 9030 25168 9036 25180
rect 9088 25208 9094 25220
rect 9125 25211 9183 25217
rect 9125 25208 9137 25211
rect 9088 25180 9137 25208
rect 9088 25168 9094 25180
rect 9125 25177 9137 25180
rect 9171 25208 9183 25211
rect 9582 25208 9588 25220
rect 9171 25180 9588 25208
rect 9171 25177 9183 25180
rect 9125 25171 9183 25177
rect 9582 25168 9588 25180
rect 9640 25168 9646 25220
rect 9214 25140 9220 25152
rect 8220 25112 9220 25140
rect 6549 25103 6607 25109
rect 9214 25100 9220 25112
rect 9272 25100 9278 25152
rect 9398 25100 9404 25152
rect 9456 25140 9462 25152
rect 10520 25140 10548 25248
rect 10576 25245 10588 25248
rect 10622 25245 10634 25279
rect 10778 25276 10784 25288
rect 10739 25248 10784 25276
rect 10576 25239 10634 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 10888 25276 10916 25372
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12802 25344 12808 25356
rect 12667 25316 12808 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 12897 25347 12955 25353
rect 12897 25313 12909 25347
rect 12943 25344 12955 25347
rect 13262 25344 13268 25356
rect 12943 25316 13268 25344
rect 12943 25313 12955 25316
rect 12897 25307 12955 25313
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 14369 25347 14427 25353
rect 14369 25344 14381 25347
rect 13556 25316 14381 25344
rect 13556 25288 13584 25316
rect 14369 25313 14381 25316
rect 14415 25313 14427 25347
rect 14369 25307 14427 25313
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 10888 25248 11713 25276
rect 11701 25245 11713 25248
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25245 11943 25279
rect 11885 25239 11943 25245
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25276 12587 25279
rect 12710 25276 12716 25288
rect 12575 25248 12716 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 10689 25211 10747 25217
rect 10689 25177 10701 25211
rect 10735 25177 10747 25211
rect 10689 25171 10747 25177
rect 10965 25211 11023 25217
rect 10965 25177 10977 25211
rect 11011 25208 11023 25211
rect 11146 25208 11152 25220
rect 11011 25180 11152 25208
rect 11011 25177 11023 25180
rect 10965 25171 11023 25177
rect 9456 25112 10548 25140
rect 10704 25140 10732 25171
rect 11146 25168 11152 25180
rect 11204 25208 11210 25220
rect 11790 25208 11796 25220
rect 11204 25180 11796 25208
rect 11204 25168 11210 25180
rect 11790 25168 11796 25180
rect 11848 25208 11854 25220
rect 11900 25208 11928 25239
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 13538 25276 13544 25288
rect 13499 25248 13544 25276
rect 13538 25236 13544 25248
rect 13596 25236 13602 25288
rect 13630 25236 13636 25288
rect 13688 25276 13694 25288
rect 14461 25279 14519 25285
rect 14461 25276 14473 25279
rect 13688 25248 14473 25276
rect 13688 25236 13694 25248
rect 14461 25245 14473 25248
rect 14507 25245 14519 25279
rect 14461 25239 14519 25245
rect 15654 25236 15660 25288
rect 15712 25276 15718 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 15712 25248 16221 25276
rect 15712 25236 15718 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 17126 25276 17132 25288
rect 17087 25248 17132 25276
rect 16209 25239 16267 25245
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 17586 25276 17592 25288
rect 17547 25248 17592 25276
rect 17586 25236 17592 25248
rect 17644 25236 17650 25288
rect 11848 25180 11928 25208
rect 11848 25168 11854 25180
rect 11054 25140 11060 25152
rect 10704 25112 11060 25140
rect 9456 25100 9462 25112
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 14458 25100 14464 25152
rect 14516 25140 14522 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14516 25112 14841 25140
rect 14516 25100 14522 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 14829 25103 14887 25109
rect 15657 25143 15715 25149
rect 15657 25109 15669 25143
rect 15703 25140 15715 25143
rect 15930 25140 15936 25152
rect 15703 25112 15936 25140
rect 15703 25109 15715 25112
rect 15657 25103 15715 25109
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 16393 25143 16451 25149
rect 16393 25109 16405 25143
rect 16439 25140 16451 25143
rect 16482 25140 16488 25152
rect 16439 25112 16488 25140
rect 16439 25109 16451 25112
rect 16393 25103 16451 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 16942 25140 16948 25152
rect 16903 25112 16948 25140
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17770 25140 17776 25152
rect 17731 25112 17776 25140
rect 17770 25100 17776 25112
rect 17828 25100 17834 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 2130 24896 2136 24948
rect 2188 24936 2194 24948
rect 3513 24939 3571 24945
rect 3513 24936 3525 24939
rect 2188 24908 3525 24936
rect 2188 24896 2194 24908
rect 3513 24905 3525 24908
rect 3559 24936 3571 24939
rect 3786 24936 3792 24948
rect 3559 24908 3792 24936
rect 3559 24905 3571 24908
rect 3513 24899 3571 24905
rect 3786 24896 3792 24908
rect 3844 24936 3850 24948
rect 5074 24936 5080 24948
rect 3844 24908 5080 24936
rect 3844 24896 3850 24908
rect 5074 24896 5080 24908
rect 5132 24896 5138 24948
rect 8389 24939 8447 24945
rect 8389 24905 8401 24939
rect 8435 24936 8447 24939
rect 8938 24936 8944 24948
rect 8435 24908 8944 24936
rect 8435 24905 8447 24908
rect 8389 24899 8447 24905
rect 8938 24896 8944 24908
rect 8996 24936 9002 24948
rect 9398 24936 9404 24948
rect 8996 24908 9404 24936
rect 8996 24896 9002 24908
rect 9398 24896 9404 24908
rect 9456 24936 9462 24948
rect 12529 24939 12587 24945
rect 9456 24908 10180 24936
rect 9456 24896 9462 24908
rect 9122 24868 9128 24880
rect 9083 24840 9128 24868
rect 9122 24828 9128 24840
rect 9180 24828 9186 24880
rect 9232 24840 9996 24868
rect 9232 24812 9260 24840
rect 7276 24803 7334 24809
rect 7276 24769 7288 24803
rect 7322 24800 7334 24803
rect 8846 24800 8852 24812
rect 7322 24772 8852 24800
rect 7322 24769 7334 24772
rect 7276 24763 7334 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 8941 24803 8999 24809
rect 8941 24769 8953 24803
rect 8987 24769 8999 24803
rect 9214 24800 9220 24812
rect 9175 24772 9220 24800
rect 8941 24763 8999 24769
rect 1949 24735 2007 24741
rect 1949 24701 1961 24735
rect 1995 24732 2007 24735
rect 4982 24732 4988 24744
rect 1995 24704 4988 24732
rect 1995 24701 2007 24704
rect 1949 24695 2007 24701
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 7006 24732 7012 24744
rect 6967 24704 7012 24732
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 8754 24692 8760 24744
rect 8812 24732 8818 24744
rect 8956 24732 8984 24763
rect 9214 24760 9220 24772
rect 9272 24760 9278 24812
rect 9345 24803 9403 24809
rect 9345 24769 9357 24803
rect 9391 24800 9403 24803
rect 9391 24772 9536 24800
rect 9391 24769 9403 24772
rect 9345 24763 9403 24769
rect 8812 24704 8984 24732
rect 9508 24732 9536 24772
rect 9582 24760 9588 24812
rect 9640 24800 9646 24812
rect 9861 24803 9919 24809
rect 9861 24800 9873 24803
rect 9640 24772 9873 24800
rect 9640 24760 9646 24772
rect 9861 24769 9873 24772
rect 9907 24769 9919 24803
rect 9968 24800 9996 24840
rect 10152 24809 10180 24908
rect 12529 24905 12541 24939
rect 12575 24936 12587 24939
rect 12710 24936 12716 24948
rect 12575 24908 12716 24936
rect 12575 24905 12587 24908
rect 12529 24899 12587 24905
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 22465 24939 22523 24945
rect 22465 24905 22477 24939
rect 22511 24936 22523 24939
rect 22511 24908 23336 24936
rect 22511 24905 22523 24908
rect 22465 24899 22523 24905
rect 11054 24828 11060 24880
rect 11112 24868 11118 24880
rect 22480 24868 22508 24899
rect 11112 24840 12572 24868
rect 11112 24828 11118 24840
rect 10045 24803 10103 24809
rect 10045 24800 10057 24803
rect 9968 24772 10057 24800
rect 9861 24763 9919 24769
rect 10045 24769 10057 24772
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10594 24800 10600 24812
rect 10555 24772 10600 24800
rect 10137 24763 10195 24769
rect 9674 24732 9680 24744
rect 9508 24704 9680 24732
rect 8812 24692 8818 24704
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 9876 24732 9904 24763
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10796 24732 10824 24763
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11020 24772 11713 24800
rect 11020 24760 11026 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 11790 24760 11796 24812
rect 11848 24800 11854 24812
rect 12544 24809 12572 24840
rect 22388 24840 22508 24868
rect 11885 24803 11943 24809
rect 11885 24800 11897 24803
rect 11848 24772 11897 24800
rect 11848 24760 11854 24772
rect 11885 24769 11897 24772
rect 11931 24769 11943 24803
rect 11885 24763 11943 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24769 12403 24803
rect 12345 24763 12403 24769
rect 12529 24803 12587 24809
rect 12529 24769 12541 24803
rect 12575 24769 12587 24803
rect 13262 24800 13268 24812
rect 13223 24772 13268 24800
rect 12529 24763 12587 24769
rect 9876 24704 10824 24732
rect 10870 24692 10876 24744
rect 10928 24732 10934 24744
rect 12360 24732 12388 24763
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 13446 24800 13452 24812
rect 13407 24772 13452 24800
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14090 24800 14096 24812
rect 13679 24772 14096 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 15188 24803 15246 24809
rect 15188 24769 15200 24803
rect 15234 24800 15246 24803
rect 17034 24800 17040 24812
rect 15234 24772 17040 24800
rect 15234 24769 15246 24772
rect 15188 24763 15246 24769
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24769 17831 24803
rect 17954 24800 17960 24812
rect 17915 24772 17960 24800
rect 17773 24763 17831 24769
rect 10928 24704 12388 24732
rect 14921 24735 14979 24741
rect 10928 24692 10934 24704
rect 14921 24701 14933 24735
rect 14967 24701 14979 24735
rect 17788 24732 17816 24763
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 18690 24800 18696 24812
rect 18651 24772 18696 24800
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 18046 24732 18052 24744
rect 17788 24704 18052 24732
rect 14921 24695 14979 24701
rect 4157 24667 4215 24673
rect 4157 24633 4169 24667
rect 4203 24664 4215 24667
rect 5718 24664 5724 24676
rect 4203 24636 5724 24664
rect 4203 24633 4215 24636
rect 4157 24627 4215 24633
rect 5718 24624 5724 24636
rect 5776 24624 5782 24676
rect 8570 24624 8576 24676
rect 8628 24664 8634 24676
rect 9861 24667 9919 24673
rect 9861 24664 9873 24667
rect 8628 24636 9873 24664
rect 8628 24624 8634 24636
rect 9861 24633 9873 24636
rect 9907 24633 9919 24667
rect 9861 24627 9919 24633
rect 2498 24596 2504 24608
rect 2459 24568 2504 24596
rect 2498 24556 2504 24568
rect 2556 24556 2562 24608
rect 2682 24556 2688 24608
rect 2740 24596 2746 24608
rect 2961 24599 3019 24605
rect 2961 24596 2973 24599
rect 2740 24568 2973 24596
rect 2740 24556 2746 24568
rect 2961 24565 2973 24568
rect 3007 24565 3019 24599
rect 2961 24559 3019 24565
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 4617 24599 4675 24605
rect 4617 24596 4629 24599
rect 4028 24568 4629 24596
rect 4028 24556 4034 24568
rect 4617 24565 4629 24568
rect 4663 24596 4675 24599
rect 5537 24599 5595 24605
rect 5537 24596 5549 24599
rect 4663 24568 5549 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 5537 24565 5549 24568
rect 5583 24565 5595 24599
rect 5537 24559 5595 24565
rect 8941 24599 8999 24605
rect 8941 24565 8953 24599
rect 8987 24596 8999 24599
rect 9766 24596 9772 24608
rect 8987 24568 9772 24596
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 10686 24596 10692 24608
rect 10647 24568 10692 24596
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 11793 24599 11851 24605
rect 11793 24565 11805 24599
rect 11839 24596 11851 24599
rect 12802 24596 12808 24608
rect 11839 24568 12808 24596
rect 11839 24565 11851 24568
rect 11793 24559 11851 24565
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 13998 24556 14004 24608
rect 14056 24596 14062 24608
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 14056 24568 14381 24596
rect 14056 24556 14062 24568
rect 14369 24565 14381 24568
rect 14415 24565 14427 24599
rect 14936 24596 14964 24695
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18892 24732 18920 24763
rect 19242 24760 19248 24812
rect 19300 24800 19306 24812
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 19300 24772 19349 24800
rect 19300 24760 19306 24772
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 19337 24763 19395 24769
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19610 24800 19616 24812
rect 19484 24772 19529 24800
rect 19571 24772 19616 24800
rect 19484 24760 19490 24772
rect 19610 24760 19616 24772
rect 19668 24760 19674 24812
rect 21266 24800 21272 24812
rect 21227 24772 21272 24800
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 21453 24803 21511 24809
rect 21453 24769 21465 24803
rect 21499 24769 21511 24803
rect 21453 24763 21511 24769
rect 21468 24732 21496 24763
rect 21542 24732 21548 24744
rect 18892 24704 19472 24732
rect 19444 24676 19472 24704
rect 19628 24704 21548 24732
rect 16301 24667 16359 24673
rect 16301 24633 16313 24667
rect 16347 24664 16359 24667
rect 17402 24664 17408 24676
rect 16347 24636 17408 24664
rect 16347 24633 16359 24636
rect 16301 24627 16359 24633
rect 17402 24624 17408 24636
rect 17460 24624 17466 24676
rect 17865 24667 17923 24673
rect 17865 24633 17877 24667
rect 17911 24664 17923 24667
rect 18230 24664 18236 24676
rect 17911 24636 18236 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 18230 24624 18236 24636
rect 18288 24664 18294 24676
rect 18874 24664 18880 24676
rect 18288 24636 18880 24664
rect 18288 24624 18294 24636
rect 18874 24624 18880 24636
rect 18932 24624 18938 24676
rect 19426 24624 19432 24676
rect 19484 24624 19490 24676
rect 19628 24673 19656 24704
rect 21542 24692 21548 24704
rect 21600 24692 21606 24744
rect 22005 24735 22063 24741
rect 22005 24701 22017 24735
rect 22051 24732 22063 24735
rect 22278 24732 22284 24744
rect 22051 24704 22284 24732
rect 22051 24701 22063 24704
rect 22005 24695 22063 24701
rect 22278 24692 22284 24704
rect 22336 24692 22342 24744
rect 19613 24667 19671 24673
rect 19613 24633 19625 24667
rect 19659 24633 19671 24667
rect 22388 24664 22416 24840
rect 23308 24812 23336 24908
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 23290 24800 23296 24812
rect 22520 24772 22565 24800
rect 23251 24772 23296 24800
rect 22520 24760 22526 24772
rect 23290 24760 23296 24772
rect 23348 24760 23354 24812
rect 23106 24692 23112 24744
rect 23164 24732 23170 24744
rect 23201 24735 23259 24741
rect 23201 24732 23213 24735
rect 23164 24704 23213 24732
rect 23164 24692 23170 24704
rect 23201 24701 23213 24704
rect 23247 24701 23259 24735
rect 23201 24695 23259 24701
rect 19613 24627 19671 24633
rect 19720 24636 22416 24664
rect 15194 24596 15200 24608
rect 14936 24568 15200 24596
rect 14369 24559 14427 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 16850 24596 16856 24608
rect 16811 24568 16856 24596
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 18782 24596 18788 24608
rect 18743 24568 18788 24596
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 18966 24556 18972 24608
rect 19024 24596 19030 24608
rect 19720 24596 19748 24636
rect 22462 24624 22468 24676
rect 22520 24664 22526 24676
rect 24486 24664 24492 24676
rect 22520 24636 24492 24664
rect 22520 24624 22526 24636
rect 24486 24624 24492 24636
rect 24544 24624 24550 24676
rect 21450 24596 21456 24608
rect 19024 24568 19748 24596
rect 21411 24568 21456 24596
rect 19024 24556 19030 24568
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 22094 24556 22100 24608
rect 22152 24596 22158 24608
rect 22649 24599 22707 24605
rect 22152 24568 22197 24596
rect 22152 24556 22158 24568
rect 22649 24565 22661 24599
rect 22695 24596 22707 24599
rect 22738 24596 22744 24608
rect 22695 24568 22744 24596
rect 22695 24565 22707 24568
rect 22649 24559 22707 24565
rect 22738 24556 22744 24568
rect 22796 24556 22802 24608
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24596 23719 24599
rect 24670 24596 24676 24608
rect 23707 24568 24676 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 5718 24392 5724 24404
rect 5679 24364 5724 24392
rect 5718 24352 5724 24364
rect 5776 24352 5782 24404
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 16574 24392 16580 24404
rect 8628 24364 11008 24392
rect 16487 24364 16580 24392
rect 8628 24352 8634 24364
rect 3421 24327 3479 24333
rect 3421 24293 3433 24327
rect 3467 24324 3479 24327
rect 4890 24324 4896 24336
rect 3467 24296 4896 24324
rect 3467 24293 3479 24296
rect 3421 24287 3479 24293
rect 4890 24284 4896 24296
rect 4948 24284 4954 24336
rect 4982 24284 4988 24336
rect 5040 24324 5046 24336
rect 6454 24324 6460 24336
rect 5040 24296 6460 24324
rect 5040 24284 5046 24296
rect 6454 24284 6460 24296
rect 6512 24284 6518 24336
rect 8754 24284 8760 24336
rect 8812 24324 8818 24336
rect 10870 24324 10876 24336
rect 8812 24296 10876 24324
rect 8812 24284 8818 24296
rect 2976 24228 5212 24256
rect 2976 24197 3004 24228
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24157 3019 24191
rect 2961 24151 3019 24157
rect 3142 24148 3148 24200
rect 3200 24188 3206 24200
rect 3237 24191 3295 24197
rect 3237 24188 3249 24191
rect 3200 24160 3249 24188
rect 3200 24148 3206 24160
rect 3237 24157 3249 24160
rect 3283 24157 3295 24191
rect 3237 24151 3295 24157
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 4982 24188 4988 24200
rect 4939 24160 4988 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 5184 24197 5212 24228
rect 9030 24216 9036 24268
rect 9088 24256 9094 24268
rect 9508 24265 9536 24296
rect 10870 24284 10876 24296
rect 10928 24284 10934 24336
rect 9309 24259 9367 24265
rect 9309 24256 9321 24259
rect 9088 24228 9321 24256
rect 9088 24216 9094 24228
rect 9309 24225 9321 24228
rect 9355 24225 9367 24259
rect 9309 24219 9367 24225
rect 9493 24259 9551 24265
rect 9493 24225 9505 24259
rect 9539 24225 9551 24259
rect 10594 24256 10600 24268
rect 9493 24219 9551 24225
rect 9692 24228 10600 24256
rect 5169 24191 5227 24197
rect 5169 24157 5181 24191
rect 5215 24188 5227 24191
rect 5350 24188 5356 24200
rect 5215 24160 5356 24188
rect 5215 24157 5227 24160
rect 5169 24151 5227 24157
rect 5350 24148 5356 24160
rect 5408 24188 5414 24200
rect 6181 24191 6239 24197
rect 6181 24188 6193 24191
rect 5408 24160 6193 24188
rect 5408 24148 5414 24160
rect 6181 24157 6193 24160
rect 6227 24157 6239 24191
rect 6454 24188 6460 24200
rect 6415 24160 6460 24188
rect 6181 24151 6239 24157
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 7064 24160 7113 24188
rect 7064 24148 7070 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9401 24191 9459 24197
rect 9401 24188 9413 24191
rect 9272 24160 9413 24188
rect 9272 24148 9278 24160
rect 9401 24157 9413 24160
rect 9447 24157 9459 24191
rect 9401 24151 9459 24157
rect 9582 24148 9588 24200
rect 9640 24188 9646 24200
rect 9692 24188 9720 24228
rect 10594 24216 10600 24228
rect 10652 24216 10658 24268
rect 9640 24160 9720 24188
rect 9640 24148 9646 24160
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 10980 24197 11008 24364
rect 16574 24352 16580 24364
rect 16632 24392 16638 24404
rect 17586 24392 17592 24404
rect 16632 24364 17592 24392
rect 16632 24352 16638 24364
rect 17586 24352 17592 24364
rect 17644 24352 17650 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 19705 24395 19763 24401
rect 19705 24392 19717 24395
rect 19668 24364 19717 24392
rect 19668 24352 19674 24364
rect 19705 24361 19717 24364
rect 19751 24392 19763 24395
rect 20441 24395 20499 24401
rect 20441 24392 20453 24395
rect 19751 24364 20453 24392
rect 19751 24361 19763 24364
rect 19705 24355 19763 24361
rect 20441 24361 20453 24364
rect 20487 24361 20499 24395
rect 23106 24392 23112 24404
rect 23067 24364 23112 24392
rect 20441 24355 20499 24361
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23569 24395 23627 24401
rect 23569 24361 23581 24395
rect 23615 24361 23627 24395
rect 23569 24355 23627 24361
rect 12802 24324 12808 24336
rect 11900 24296 12808 24324
rect 10137 24191 10195 24197
rect 10137 24188 10149 24191
rect 9824 24160 10149 24188
rect 9824 24148 9830 24160
rect 10137 24157 10149 24160
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 10965 24191 11023 24197
rect 10965 24157 10977 24191
rect 11011 24157 11023 24191
rect 11146 24188 11152 24200
rect 11107 24160 11152 24188
rect 10965 24151 11023 24157
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 11900 24197 11928 24296
rect 12802 24284 12808 24296
rect 12860 24284 12866 24336
rect 19889 24327 19947 24333
rect 19889 24293 19901 24327
rect 19935 24293 19947 24327
rect 19889 24287 19947 24293
rect 22005 24327 22063 24333
rect 22005 24293 22017 24327
rect 22051 24324 22063 24327
rect 22094 24324 22100 24336
rect 22051 24296 22100 24324
rect 22051 24293 22063 24296
rect 22005 24287 22063 24293
rect 11977 24259 12035 24265
rect 11977 24225 11989 24259
rect 12023 24225 12035 24259
rect 11977 24219 12035 24225
rect 13081 24259 13139 24265
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 13906 24256 13912 24268
rect 13127 24228 13912 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 3053 24123 3111 24129
rect 3053 24089 3065 24123
rect 3099 24120 3111 24123
rect 4246 24120 4252 24132
rect 3099 24092 4252 24120
rect 3099 24089 3111 24092
rect 3053 24083 3111 24089
rect 4246 24080 4252 24092
rect 4304 24080 4310 24132
rect 6270 24120 6276 24132
rect 6231 24092 6276 24120
rect 6270 24080 6276 24092
rect 6328 24080 6334 24132
rect 7368 24123 7426 24129
rect 7368 24089 7380 24123
rect 7414 24120 7426 24123
rect 9030 24120 9036 24132
rect 7414 24092 9036 24120
rect 7414 24089 7426 24092
rect 7368 24083 7426 24089
rect 9030 24080 9036 24092
rect 9088 24080 9094 24132
rect 9306 24120 9312 24132
rect 9140 24092 9312 24120
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 2222 24052 2228 24064
rect 2183 24024 2228 24052
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 4157 24055 4215 24061
rect 4157 24052 4169 24055
rect 4028 24024 4169 24052
rect 4028 24012 4034 24024
rect 4157 24021 4169 24024
rect 4203 24021 4215 24055
rect 4157 24015 4215 24021
rect 4709 24055 4767 24061
rect 4709 24021 4721 24055
rect 4755 24052 4767 24055
rect 4798 24052 4804 24064
rect 4755 24024 4804 24052
rect 4755 24021 4767 24024
rect 4709 24015 4767 24021
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 5077 24055 5135 24061
rect 5077 24021 5089 24055
rect 5123 24052 5135 24055
rect 5442 24052 5448 24064
rect 5123 24024 5448 24052
rect 5123 24021 5135 24024
rect 5077 24015 5135 24021
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 6638 24052 6644 24064
rect 6599 24024 6644 24052
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 8478 24052 8484 24064
rect 8439 24024 8484 24052
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 9140 24061 9168 24092
rect 9306 24080 9312 24092
rect 9364 24120 9370 24132
rect 10321 24123 10379 24129
rect 10321 24120 10333 24123
rect 9364 24092 10333 24120
rect 9364 24080 9370 24092
rect 10321 24089 10333 24092
rect 10367 24089 10379 24123
rect 10321 24083 10379 24089
rect 9125 24055 9183 24061
rect 9125 24021 9137 24055
rect 9171 24021 9183 24055
rect 9125 24015 9183 24021
rect 10505 24055 10563 24061
rect 10505 24021 10517 24055
rect 10551 24052 10563 24055
rect 10594 24052 10600 24064
rect 10551 24024 10600 24052
rect 10551 24021 10563 24024
rect 10505 24015 10563 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 10962 24052 10968 24064
rect 10923 24024 10968 24052
rect 10962 24012 10968 24024
rect 11020 24052 11026 24064
rect 11992 24052 12020 24219
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 19904 24256 19932 24287
rect 22094 24284 22100 24296
rect 22152 24324 22158 24336
rect 23584 24324 23612 24355
rect 22152 24296 23612 24324
rect 22152 24284 22158 24296
rect 21266 24256 21272 24268
rect 19904 24228 21272 24256
rect 21266 24216 21272 24228
rect 21324 24256 21330 24268
rect 22738 24256 22744 24268
rect 21324 24228 21404 24256
rect 22699 24228 22744 24256
rect 21324 24216 21330 24228
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 12124 24160 12173 24188
rect 12124 24148 12130 24160
rect 12161 24157 12173 24160
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 13541 24191 13599 24197
rect 12308 24160 12353 24188
rect 12308 24148 12314 24160
rect 13541 24157 13553 24191
rect 13587 24157 13599 24191
rect 13722 24188 13728 24200
rect 13683 24160 13728 24188
rect 13541 24151 13599 24157
rect 13556 24120 13584 24151
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 15194 24188 15200 24200
rect 15155 24160 15200 24188
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 18046 24188 18052 24200
rect 17359 24160 18052 24188
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 18690 24188 18696 24200
rect 18647 24160 18696 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 18874 24188 18880 24200
rect 18835 24160 18880 24188
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 19242 24148 19248 24200
rect 19300 24188 19306 24200
rect 19300 24160 19656 24188
rect 19300 24148 19306 24160
rect 14642 24120 14648 24132
rect 13556 24092 14648 24120
rect 14642 24080 14648 24092
rect 14700 24080 14706 24132
rect 15464 24123 15522 24129
rect 15464 24089 15476 24123
rect 15510 24120 15522 24123
rect 15746 24120 15752 24132
rect 15510 24092 15752 24120
rect 15510 24089 15522 24092
rect 15464 24083 15522 24089
rect 15746 24080 15752 24092
rect 15804 24080 15810 24132
rect 19518 24120 19524 24132
rect 19479 24092 19524 24120
rect 19518 24080 19524 24092
rect 19576 24080 19582 24132
rect 19628 24120 19656 24160
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 21376 24197 21404 24228
rect 22738 24216 22744 24228
rect 22796 24216 22802 24268
rect 22833 24259 22891 24265
rect 22833 24225 22845 24259
rect 22879 24256 22891 24259
rect 23198 24256 23204 24268
rect 22879 24228 23204 24256
rect 22879 24225 22891 24228
rect 22833 24219 22891 24225
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 24670 24256 24676 24268
rect 24631 24228 24676 24256
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 20128 24160 20361 24188
rect 20128 24148 20134 24160
rect 20349 24157 20361 24160
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21542 24188 21548 24200
rect 21503 24160 21548 24188
rect 21361 24151 21419 24157
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24157 21879 24191
rect 22462 24188 22468 24200
rect 22423 24160 22468 24188
rect 21821 24151 21879 24157
rect 19721 24123 19779 24129
rect 19721 24120 19733 24123
rect 19628 24092 19733 24120
rect 19721 24089 19733 24092
rect 19767 24089 19779 24123
rect 19721 24083 19779 24089
rect 11020 24024 12020 24052
rect 12437 24055 12495 24061
rect 11020 24012 11026 24024
rect 12437 24021 12449 24055
rect 12483 24052 12495 24055
rect 12894 24052 12900 24064
rect 12483 24024 12900 24052
rect 12483 24021 12495 24024
rect 12437 24015 12495 24021
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 13630 24052 13636 24064
rect 13591 24024 13636 24052
rect 13630 24012 13636 24024
rect 13688 24012 13694 24064
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 13872 24024 14289 24052
rect 13872 24012 13878 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 17773 24055 17831 24061
rect 17773 24021 17785 24055
rect 17819 24052 17831 24055
rect 17862 24052 17868 24064
rect 17819 24024 17868 24052
rect 17819 24021 17831 24024
rect 17773 24015 17831 24021
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 18417 24055 18475 24061
rect 18417 24021 18429 24055
rect 18463 24052 18475 24055
rect 18506 24052 18512 24064
rect 18463 24024 18512 24052
rect 18463 24021 18475 24024
rect 18417 24015 18475 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 18785 24055 18843 24061
rect 18785 24021 18797 24055
rect 18831 24052 18843 24055
rect 19426 24052 19432 24064
rect 18831 24024 19432 24052
rect 18831 24021 18843 24024
rect 18785 24015 18843 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 21266 24012 21272 24064
rect 21324 24052 21330 24064
rect 21836 24052 21864 24151
rect 22462 24148 22468 24160
rect 22520 24148 22526 24200
rect 22646 24188 22652 24200
rect 22607 24160 22652 24188
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 22925 24191 22983 24197
rect 22925 24157 22937 24191
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 22186 24080 22192 24132
rect 22244 24120 22250 24132
rect 22940 24120 22968 24151
rect 23474 24148 23480 24200
rect 23532 24188 23538 24200
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 23532 24160 23581 24188
rect 23532 24148 23538 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 24765 24191 24823 24197
rect 24765 24188 24777 24191
rect 23661 24151 23719 24157
rect 23952 24160 24777 24188
rect 22244 24092 22968 24120
rect 22244 24080 22250 24092
rect 23382 24080 23388 24132
rect 23440 24120 23446 24132
rect 23676 24120 23704 24151
rect 23750 24120 23756 24132
rect 23440 24092 23756 24120
rect 23440 24080 23446 24092
rect 23750 24080 23756 24092
rect 23808 24080 23814 24132
rect 23566 24052 23572 24064
rect 21324 24024 23572 24052
rect 21324 24012 21330 24024
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 23952 24061 23980 24160
rect 24765 24157 24777 24160
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 23937 24055 23995 24061
rect 23937 24021 23949 24055
rect 23983 24021 23995 24055
rect 23937 24015 23995 24021
rect 24854 24012 24860 24064
rect 24912 24052 24918 24064
rect 25133 24055 25191 24061
rect 25133 24052 25145 24055
rect 24912 24024 25145 24052
rect 24912 24012 24918 24024
rect 25133 24021 25145 24024
rect 25179 24021 25191 24055
rect 25133 24015 25191 24021
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 2682 23848 2688 23860
rect 1688 23820 2688 23848
rect 1688 23789 1716 23820
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 5629 23851 5687 23857
rect 5629 23817 5641 23851
rect 5675 23848 5687 23851
rect 8754 23848 8760 23860
rect 5675 23820 8760 23848
rect 5675 23817 5687 23820
rect 5629 23811 5687 23817
rect 8754 23808 8760 23820
rect 8812 23808 8818 23860
rect 9030 23848 9036 23860
rect 8991 23820 9036 23848
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10686 23848 10692 23860
rect 10192 23820 10692 23848
rect 10192 23808 10198 23820
rect 10686 23808 10692 23820
rect 10744 23848 10750 23860
rect 10781 23851 10839 23857
rect 10781 23848 10793 23851
rect 10744 23820 10793 23848
rect 10744 23808 10750 23820
rect 10781 23817 10793 23820
rect 10827 23817 10839 23851
rect 15746 23848 15752 23860
rect 15707 23820 15752 23848
rect 10781 23811 10839 23817
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 16117 23851 16175 23857
rect 16117 23817 16129 23851
rect 16163 23848 16175 23851
rect 16574 23848 16580 23860
rect 16163 23820 16580 23848
rect 16163 23817 16175 23820
rect 16117 23811 16175 23817
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 17402 23808 17408 23820
rect 17460 23848 17466 23860
rect 18506 23848 18512 23860
rect 17460 23820 17908 23848
rect 18467 23820 18512 23848
rect 17460 23808 17466 23820
rect 1673 23783 1731 23789
rect 1673 23749 1685 23783
rect 1719 23749 1731 23783
rect 1854 23780 1860 23792
rect 1815 23752 1860 23780
rect 1673 23743 1731 23749
rect 1854 23740 1860 23752
rect 1912 23740 1918 23792
rect 8478 23740 8484 23792
rect 8536 23780 8542 23792
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 8536 23752 9413 23780
rect 8536 23740 8542 23752
rect 9401 23749 9413 23752
rect 9447 23780 9459 23783
rect 9674 23780 9680 23792
rect 9447 23752 9680 23780
rect 9447 23749 9459 23752
rect 9401 23743 9459 23749
rect 9674 23740 9680 23752
rect 9732 23740 9738 23792
rect 14737 23783 14795 23789
rect 14737 23749 14749 23783
rect 14783 23780 14795 23783
rect 15194 23780 15200 23792
rect 14783 23752 15200 23780
rect 14783 23749 14795 23752
rect 14737 23743 14795 23749
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 4338 23712 4344 23724
rect 4299 23684 4344 23712
rect 2133 23675 2191 23681
rect 2148 23644 2176 23675
rect 4338 23672 4344 23684
rect 4396 23672 4402 23724
rect 5350 23672 5356 23724
rect 5408 23712 5414 23724
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 5408 23684 5549 23712
rect 5408 23672 5414 23684
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 5810 23712 5816 23724
rect 5723 23684 5816 23712
rect 5537 23675 5595 23681
rect 5810 23672 5816 23684
rect 5868 23712 5874 23724
rect 6362 23712 6368 23724
rect 5868 23684 6368 23712
rect 5868 23672 5874 23684
rect 6362 23672 6368 23684
rect 6420 23672 6426 23724
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23712 6883 23715
rect 7466 23712 7472 23724
rect 6871 23684 7472 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 7282 23644 7288 23656
rect 2148 23616 7288 23644
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 9232 23644 9260 23675
rect 9490 23672 9496 23724
rect 9548 23712 9554 23724
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 9548 23684 9593 23712
rect 9968 23684 10149 23712
rect 9548 23672 9554 23684
rect 9858 23644 9864 23656
rect 9232 23616 9864 23644
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 3970 23536 3976 23588
rect 4028 23576 4034 23588
rect 4985 23579 5043 23585
rect 4985 23576 4997 23579
rect 4028 23548 4997 23576
rect 4028 23536 4034 23548
rect 4985 23545 4997 23548
rect 5031 23545 5043 23579
rect 4985 23539 5043 23545
rect 5258 23536 5264 23588
rect 5316 23576 5322 23588
rect 8113 23579 8171 23585
rect 8113 23576 8125 23579
rect 5316 23548 8125 23576
rect 5316 23536 5322 23548
rect 8113 23545 8125 23548
rect 8159 23545 8171 23579
rect 8113 23539 8171 23545
rect 9582 23536 9588 23588
rect 9640 23576 9646 23588
rect 9968 23576 9996 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 10594 23672 10600 23724
rect 10652 23712 10658 23724
rect 10689 23715 10747 23721
rect 10689 23712 10701 23715
rect 10652 23684 10701 23712
rect 10652 23672 10658 23684
rect 10689 23681 10701 23684
rect 10735 23681 10747 23715
rect 10962 23712 10968 23724
rect 10875 23684 10968 23712
rect 10689 23675 10747 23681
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 11698 23672 11704 23724
rect 11756 23712 11762 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 11756 23684 12081 23712
rect 11756 23672 11762 23684
rect 12069 23681 12081 23684
rect 12115 23712 12127 23715
rect 12250 23712 12256 23724
rect 12115 23684 12256 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 12529 23715 12587 23721
rect 12529 23681 12541 23715
rect 12575 23712 12587 23715
rect 12802 23712 12808 23724
rect 12575 23684 12808 23712
rect 12575 23681 12587 23684
rect 12529 23675 12587 23681
rect 10226 23604 10232 23656
rect 10284 23644 10290 23656
rect 10980 23644 11008 23672
rect 12360 23644 12388 23675
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 12989 23715 13047 23721
rect 12989 23681 13001 23715
rect 13035 23712 13047 23715
rect 15838 23712 15844 23724
rect 13035 23684 15844 23712
rect 13035 23681 13047 23684
rect 12989 23675 13047 23681
rect 15212 23656 15240 23684
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 15930 23672 15936 23724
rect 15988 23712 15994 23724
rect 16209 23715 16267 23721
rect 15988 23684 16033 23712
rect 15988 23672 15994 23684
rect 16209 23681 16221 23715
rect 16255 23712 16267 23715
rect 16850 23712 16856 23724
rect 16255 23684 16856 23712
rect 16255 23681 16267 23684
rect 16209 23675 16267 23681
rect 10284 23616 12388 23644
rect 10284 23604 10290 23616
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 16022 23576 16028 23588
rect 9640 23548 9996 23576
rect 15212 23548 16028 23576
rect 9640 23536 9646 23548
rect 1857 23511 1915 23517
rect 1857 23477 1869 23511
rect 1903 23508 1915 23511
rect 2130 23508 2136 23520
rect 1903 23480 2136 23508
rect 1903 23477 1915 23480
rect 1857 23471 1915 23477
rect 2130 23468 2136 23480
rect 2188 23468 2194 23520
rect 2866 23468 2872 23520
rect 2924 23508 2930 23520
rect 3053 23511 3111 23517
rect 3053 23508 3065 23511
rect 2924 23480 3065 23508
rect 2924 23468 2930 23480
rect 3053 23477 3065 23480
rect 3099 23508 3111 23511
rect 4062 23508 4068 23520
rect 3099 23480 4068 23508
rect 3099 23477 3111 23480
rect 3053 23471 3111 23477
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 5997 23511 6055 23517
rect 5997 23477 6009 23511
rect 6043 23508 6055 23511
rect 6730 23508 6736 23520
rect 6043 23480 6736 23508
rect 6043 23477 6055 23480
rect 5997 23471 6055 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 9548 23480 10057 23508
rect 9548 23468 9554 23480
rect 10045 23477 10057 23480
rect 10091 23477 10103 23511
rect 10045 23471 10103 23477
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 11238 23508 11244 23520
rect 11195 23480 11244 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 11238 23468 11244 23480
rect 11296 23468 11302 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12066 23508 12072 23520
rect 11931 23480 12072 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 13998 23468 14004 23520
rect 14056 23508 14062 23520
rect 15212 23517 15240 23548
rect 16022 23536 16028 23548
rect 16080 23576 16086 23588
rect 16224 23576 16252 23675
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23681 17555 23715
rect 17880 23712 17908 23820
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 18690 23808 18696 23860
rect 18748 23848 18754 23860
rect 20165 23851 20223 23857
rect 20165 23848 20177 23851
rect 18748 23820 20177 23848
rect 18748 23808 18754 23820
rect 20165 23817 20177 23820
rect 20211 23817 20223 23851
rect 20165 23811 20223 23817
rect 21177 23851 21235 23857
rect 21177 23817 21189 23851
rect 21223 23848 21235 23851
rect 22278 23848 22284 23860
rect 21223 23820 22284 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22370 23808 22376 23860
rect 22428 23848 22434 23860
rect 23198 23848 23204 23860
rect 22428 23820 23204 23848
rect 22428 23808 22434 23820
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23348 23820 24348 23848
rect 23348 23808 23354 23820
rect 17954 23740 17960 23792
rect 18012 23780 18018 23792
rect 18601 23783 18659 23789
rect 18601 23780 18613 23783
rect 18012 23752 18613 23780
rect 18012 23740 18018 23752
rect 18601 23749 18613 23752
rect 18647 23749 18659 23783
rect 21450 23780 21456 23792
rect 21411 23752 21456 23780
rect 18601 23743 18659 23749
rect 21450 23740 21456 23752
rect 21508 23780 21514 23792
rect 21508 23752 23428 23780
rect 21508 23740 21514 23752
rect 19429 23715 19487 23721
rect 19429 23712 19441 23715
rect 17880 23684 19441 23712
rect 17497 23675 17555 23681
rect 19429 23681 19441 23684
rect 19475 23681 19487 23715
rect 20070 23712 20076 23724
rect 19983 23684 20076 23712
rect 19429 23675 19487 23681
rect 16868 23644 16896 23672
rect 17512 23644 17540 23675
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 20254 23712 20260 23724
rect 20215 23684 20260 23712
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 21085 23715 21143 23721
rect 21085 23712 21097 23715
rect 20496 23684 21097 23712
rect 20496 23672 20502 23684
rect 21085 23681 21097 23684
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 21361 23715 21419 23721
rect 21361 23681 21373 23715
rect 21407 23712 21419 23715
rect 21407 23684 22094 23712
rect 21407 23681 21419 23684
rect 21361 23675 21419 23681
rect 16868 23616 17540 23644
rect 18046 23604 18052 23656
rect 18104 23644 18110 23656
rect 18325 23647 18383 23653
rect 18325 23644 18337 23647
rect 18104 23616 18337 23644
rect 18104 23604 18110 23616
rect 18325 23613 18337 23616
rect 18371 23644 18383 23647
rect 19242 23644 19248 23656
rect 18371 23616 19248 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 20088 23644 20116 23672
rect 19352 23616 20116 23644
rect 18966 23576 18972 23588
rect 16080 23548 16252 23576
rect 18927 23548 18972 23576
rect 16080 23536 16086 23548
rect 18966 23536 18972 23548
rect 19024 23536 19030 23588
rect 15197 23511 15255 23517
rect 15197 23508 15209 23511
rect 14056 23480 15209 23508
rect 14056 23468 14062 23480
rect 15197 23477 15209 23480
rect 15243 23477 15255 23511
rect 15197 23471 15255 23477
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 19352 23508 19380 23616
rect 21100 23576 21128 23675
rect 22066 23644 22094 23684
rect 22186 23672 22192 23724
rect 22244 23712 22250 23724
rect 22244 23684 22289 23712
rect 22244 23672 22250 23684
rect 22370 23672 22376 23724
rect 22428 23712 22434 23724
rect 22557 23715 22615 23721
rect 22428 23684 22473 23712
rect 22428 23672 22434 23684
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22738 23712 22744 23724
rect 22603 23684 22744 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23400 23721 23428 23752
rect 22833 23715 22891 23721
rect 22833 23681 22845 23715
rect 22879 23681 22891 23715
rect 22833 23675 22891 23681
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23566 23712 23572 23724
rect 23527 23684 23572 23712
rect 23385 23675 23443 23681
rect 22066 23616 22232 23644
rect 22204 23576 22232 23616
rect 22278 23604 22284 23656
rect 22336 23644 22342 23656
rect 22646 23644 22652 23656
rect 22336 23616 22652 23644
rect 22336 23604 22342 23616
rect 22646 23604 22652 23616
rect 22704 23644 22710 23656
rect 22848 23644 22876 23675
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23712 23719 23715
rect 23750 23712 23756 23724
rect 23707 23684 23756 23712
rect 23707 23681 23719 23684
rect 23661 23675 23719 23681
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 24320 23721 24348 23820
rect 24305 23715 24363 23721
rect 24305 23681 24317 23715
rect 24351 23681 24363 23715
rect 24486 23712 24492 23724
rect 24447 23684 24492 23712
rect 24305 23675 24363 23681
rect 24486 23672 24492 23684
rect 24544 23672 24550 23724
rect 24578 23672 24584 23724
rect 24636 23712 24642 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 24636 23684 25053 23712
rect 24636 23672 24642 23684
rect 25041 23681 25053 23684
rect 25087 23681 25099 23715
rect 25041 23675 25099 23681
rect 25225 23715 25283 23721
rect 25225 23681 25237 23715
rect 25271 23712 25283 23715
rect 25590 23712 25596 23724
rect 25271 23684 25596 23712
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 23474 23644 23480 23656
rect 22704 23616 22876 23644
rect 23435 23616 23480 23644
rect 22704 23604 22710 23616
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 22462 23576 22468 23588
rect 21100 23548 22094 23576
rect 22204 23548 22468 23576
rect 19518 23508 19524 23520
rect 16448 23480 19380 23508
rect 19479 23480 19524 23508
rect 16448 23468 16454 23480
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 21266 23508 21272 23520
rect 21227 23480 21272 23508
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 22066 23508 22094 23548
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 22833 23579 22891 23585
rect 22833 23545 22845 23579
rect 22879 23576 22891 23579
rect 23492 23576 23520 23604
rect 24305 23579 24363 23585
rect 24305 23576 24317 23579
rect 22879 23548 23520 23576
rect 23584 23548 24317 23576
rect 22879 23545 22891 23548
rect 22833 23539 22891 23545
rect 22848 23508 22876 23539
rect 22066 23480 22876 23508
rect 23198 23468 23204 23520
rect 23256 23508 23262 23520
rect 23584 23508 23612 23548
rect 24305 23545 24317 23548
rect 24351 23545 24363 23579
rect 24305 23539 24363 23545
rect 23842 23508 23848 23520
rect 23256 23480 23612 23508
rect 23803 23480 23848 23508
rect 23256 23468 23262 23480
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 25130 23508 25136 23520
rect 25091 23480 25136 23508
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 7466 23304 7472 23316
rect 7427 23276 7472 23304
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 8846 23264 8852 23316
rect 8904 23304 8910 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 8904 23276 9137 23304
rect 8904 23264 8910 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 15838 23264 15844 23316
rect 15896 23304 15902 23316
rect 16393 23307 16451 23313
rect 16393 23304 16405 23307
rect 15896 23276 16405 23304
rect 15896 23264 15902 23276
rect 16393 23273 16405 23276
rect 16439 23273 16451 23307
rect 16393 23267 16451 23273
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 17313 23307 17371 23313
rect 17313 23304 17325 23307
rect 16908 23276 17325 23304
rect 16908 23264 16914 23276
rect 17313 23273 17325 23276
rect 17359 23273 17371 23307
rect 17313 23267 17371 23273
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 18049 23307 18107 23313
rect 18049 23304 18061 23307
rect 18012 23276 18061 23304
rect 18012 23264 18018 23276
rect 18049 23273 18061 23276
rect 18095 23273 18107 23307
rect 18049 23267 18107 23273
rect 18138 23264 18144 23316
rect 18196 23264 18202 23316
rect 19426 23304 19432 23316
rect 19387 23276 19432 23304
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 22738 23304 22744 23316
rect 22112 23276 22744 23304
rect 12437 23239 12495 23245
rect 12437 23236 12449 23239
rect 11440 23208 12449 23236
rect 2590 23168 2596 23180
rect 2240 23140 2596 23168
rect 2130 23060 2136 23112
rect 2188 23100 2194 23112
rect 2240 23109 2268 23140
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 3050 23168 3056 23180
rect 2700 23140 3056 23168
rect 2225 23103 2283 23109
rect 2225 23100 2237 23103
rect 2188 23072 2237 23100
rect 2188 23060 2194 23072
rect 2225 23069 2237 23072
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23100 2559 23103
rect 2700 23100 2728 23140
rect 3050 23128 3056 23140
rect 3108 23168 3114 23180
rect 5074 23168 5080 23180
rect 3108 23140 5080 23168
rect 3108 23128 3114 23140
rect 2547 23072 2728 23100
rect 3145 23103 3203 23109
rect 2547 23069 2559 23072
rect 2501 23063 2559 23069
rect 3145 23069 3157 23103
rect 3191 23069 3203 23103
rect 3145 23063 3203 23069
rect 3421 23103 3479 23109
rect 3421 23069 3433 23103
rect 3467 23100 3479 23103
rect 3694 23100 3700 23112
rect 3467 23072 3700 23100
rect 3467 23069 3479 23072
rect 3421 23063 3479 23069
rect 3160 23032 3188 23063
rect 3694 23060 3700 23072
rect 3752 23060 3758 23112
rect 4356 23109 4384 23140
rect 5074 23128 5080 23140
rect 5132 23168 5138 23180
rect 5350 23168 5356 23180
rect 5132 23140 5356 23168
rect 5132 23128 5138 23140
rect 5350 23128 5356 23140
rect 5408 23128 5414 23180
rect 7006 23168 7012 23180
rect 6967 23140 7012 23168
rect 7006 23128 7012 23140
rect 7064 23128 7070 23180
rect 9398 23168 9404 23180
rect 8588 23140 9404 23168
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23069 4675 23103
rect 5258 23100 5264 23112
rect 5219 23072 5264 23100
rect 4617 23063 4675 23069
rect 4632 23032 4660 23063
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 7650 23100 7656 23112
rect 7611 23072 7656 23100
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 8294 23100 8300 23112
rect 8255 23072 8300 23100
rect 8294 23060 8300 23072
rect 8352 23060 8358 23112
rect 8478 23060 8484 23112
rect 8536 23100 8542 23112
rect 8588 23109 8616 23140
rect 9398 23128 9404 23140
rect 9456 23168 9462 23180
rect 11330 23168 11336 23180
rect 9456 23140 11336 23168
rect 9456 23128 9462 23140
rect 8573 23103 8631 23109
rect 8573 23100 8585 23103
rect 8536 23072 8585 23100
rect 8536 23060 8542 23072
rect 8573 23069 8585 23072
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9600 23109 9628 23140
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9088 23072 9321 23100
rect 9088 23060 9094 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 5350 23032 5356 23044
rect 2240 23004 4660 23032
rect 4724 23004 5356 23032
rect 2240 22976 2268 23004
rect 2038 22964 2044 22976
rect 1999 22936 2044 22964
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 2222 22924 2228 22976
rect 2280 22924 2286 22976
rect 2406 22964 2412 22976
rect 2367 22936 2412 22964
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 2958 22964 2964 22976
rect 2919 22936 2964 22964
rect 2958 22924 2964 22936
rect 3016 22924 3022 22976
rect 3234 22924 3240 22976
rect 3292 22964 3298 22976
rect 3329 22967 3387 22973
rect 3329 22964 3341 22967
rect 3292 22936 3341 22964
rect 3292 22924 3298 22936
rect 3329 22933 3341 22936
rect 3375 22933 3387 22967
rect 3329 22927 3387 22933
rect 4433 22967 4491 22973
rect 4433 22933 4445 22967
rect 4479 22964 4491 22967
rect 4724 22964 4752 23004
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 9324 23032 9352 23063
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 10410 23100 10416 23112
rect 9916 23072 10416 23100
rect 9916 23060 9922 23072
rect 10410 23060 10416 23072
rect 10468 23100 10474 23112
rect 10796 23109 10824 23140
rect 11330 23128 11336 23140
rect 11388 23128 11394 23180
rect 10505 23103 10563 23109
rect 10505 23100 10517 23103
rect 10468 23072 10517 23100
rect 10468 23060 10474 23072
rect 10505 23069 10517 23072
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 11238 23100 11244 23112
rect 11199 23072 11244 23100
rect 10781 23063 10839 23069
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11440 23109 11468 23208
rect 12437 23205 12449 23208
rect 12483 23236 12495 23239
rect 18156 23236 18184 23264
rect 19242 23236 19248 23248
rect 12483 23208 14504 23236
rect 18156 23208 19248 23236
rect 12483 23205 12495 23208
rect 12437 23199 12495 23205
rect 12158 23168 12164 23180
rect 12119 23140 12164 23168
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 12894 23128 12900 23180
rect 12952 23168 12958 23180
rect 13262 23168 13268 23180
rect 12952 23140 13268 23168
rect 12952 23128 12958 23140
rect 13262 23128 13268 23140
rect 13320 23128 13326 23180
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23069 11483 23103
rect 12066 23100 12072 23112
rect 12027 23072 12072 23100
rect 11425 23063 11483 23069
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 13354 23100 13360 23112
rect 13315 23072 13360 23100
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 14476 23109 14504 23208
rect 19242 23196 19248 23208
rect 19300 23236 19306 23248
rect 21082 23236 21088 23248
rect 19300 23208 21088 23236
rect 19300 23196 19306 23208
rect 18138 23128 18144 23180
rect 18196 23168 18202 23180
rect 18417 23171 18475 23177
rect 18417 23168 18429 23171
rect 18196 23140 18429 23168
rect 18196 23128 18202 23140
rect 18417 23137 18429 23140
rect 18463 23137 18475 23171
rect 18417 23131 18475 23137
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23168 18567 23171
rect 19518 23168 19524 23180
rect 18555 23140 19524 23168
rect 18555 23137 18567 23140
rect 18509 23131 18567 23137
rect 19518 23128 19524 23140
rect 19576 23168 19582 23180
rect 19576 23140 19932 23168
rect 19576 23128 19582 23140
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 18233 23103 18291 23109
rect 18233 23100 18245 23103
rect 17920 23072 18245 23100
rect 17920 23060 17926 23072
rect 18233 23069 18245 23072
rect 18279 23069 18291 23103
rect 18233 23063 18291 23069
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23100 18383 23103
rect 19334 23100 19340 23112
rect 18371 23072 19340 23100
rect 18371 23069 18383 23072
rect 18325 23063 18383 23069
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 19392 23072 19625 23100
rect 19392 23060 19398 23072
rect 19613 23069 19625 23072
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 19702 23060 19708 23112
rect 19760 23100 19766 23112
rect 19904 23109 19932 23140
rect 19996 23109 20024 23208
rect 21082 23196 21088 23208
rect 21140 23196 21146 23248
rect 22112 23245 22140 23276
rect 22738 23264 22744 23276
rect 22796 23304 22802 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22796 23276 22937 23304
rect 22796 23264 22802 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 22925 23267 22983 23273
rect 22097 23239 22155 23245
rect 22097 23205 22109 23239
rect 22143 23205 22155 23239
rect 22097 23199 22155 23205
rect 23385 23239 23443 23245
rect 23385 23205 23397 23239
rect 23431 23236 23443 23239
rect 23431 23208 25176 23236
rect 23431 23205 23443 23208
rect 23385 23199 23443 23205
rect 20530 23128 20536 23180
rect 20588 23168 20594 23180
rect 24578 23168 24584 23180
rect 20588 23140 22416 23168
rect 20588 23128 20594 23140
rect 19889 23103 19947 23109
rect 19760 23072 19805 23100
rect 19760 23060 19766 23072
rect 19889 23069 19901 23103
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 20901 23103 20959 23109
rect 20901 23069 20913 23103
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 10042 23032 10048 23044
rect 9324 23004 10048 23032
rect 10042 22992 10048 23004
rect 10100 23032 10106 23044
rect 10870 23032 10876 23044
rect 10100 23004 10876 23032
rect 10100 22992 10106 23004
rect 10870 22992 10876 23004
rect 10928 22992 10934 23044
rect 11256 23032 11284 23060
rect 11882 23032 11888 23044
rect 11256 23004 11888 23032
rect 11882 22992 11888 23004
rect 11940 23032 11946 23044
rect 14277 23035 14335 23041
rect 14277 23032 14289 23035
rect 11940 23004 14289 23032
rect 11940 22992 11946 23004
rect 14277 23001 14289 23004
rect 14323 23001 14335 23035
rect 14277 22995 14335 23001
rect 14550 22992 14556 23044
rect 14608 23032 14614 23044
rect 15105 23035 15163 23041
rect 15105 23032 15117 23035
rect 14608 23004 15117 23032
rect 14608 22992 14614 23004
rect 15105 23001 15117 23004
rect 15151 23001 15163 23035
rect 15105 22995 15163 23001
rect 18690 22992 18696 23044
rect 18748 23032 18754 23044
rect 20916 23032 20944 23063
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21085 23103 21143 23109
rect 21085 23100 21097 23103
rect 21048 23072 21097 23100
rect 21048 23060 21054 23072
rect 21085 23069 21097 23072
rect 21131 23069 21143 23103
rect 21085 23063 21143 23069
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23100 21327 23103
rect 21910 23100 21916 23112
rect 21315 23072 21916 23100
rect 21315 23069 21327 23072
rect 21269 23063 21327 23069
rect 18748 23004 20944 23032
rect 21100 23032 21128 23063
rect 21910 23060 21916 23072
rect 21968 23060 21974 23112
rect 22005 23103 22063 23109
rect 22005 23069 22017 23103
rect 22051 23069 22063 23103
rect 22005 23063 22063 23069
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23100 22247 23103
rect 22278 23100 22284 23112
rect 22235 23072 22284 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22020 23032 22048 23063
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22388 23109 22416 23140
rect 22848 23140 24584 23168
rect 22848 23109 22876 23140
rect 24578 23128 24584 23140
rect 24636 23128 24642 23180
rect 25148 23177 25176 23208
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 22373 23103 22431 23109
rect 22373 23069 22385 23103
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23069 22891 23103
rect 23198 23100 23204 23112
rect 23159 23072 23204 23100
rect 22833 23063 22891 23069
rect 22462 23032 22468 23044
rect 21100 23004 21864 23032
rect 22020 23004 22468 23032
rect 18748 22992 18754 23004
rect 4479 22936 4752 22964
rect 4801 22967 4859 22973
rect 4479 22933 4491 22936
rect 4433 22927 4491 22933
rect 4801 22933 4813 22967
rect 4847 22964 4859 22967
rect 4982 22964 4988 22976
rect 4847 22936 4988 22964
rect 4847 22933 4859 22936
rect 4801 22927 4859 22933
rect 4982 22924 4988 22936
rect 5040 22924 5046 22976
rect 7742 22924 7748 22976
rect 7800 22964 7806 22976
rect 8113 22967 8171 22973
rect 8113 22964 8125 22967
rect 7800 22936 8125 22964
rect 7800 22924 7806 22936
rect 8113 22933 8125 22936
rect 8159 22933 8171 22967
rect 8113 22927 8171 22933
rect 8481 22967 8539 22973
rect 8481 22933 8493 22967
rect 8527 22964 8539 22967
rect 9122 22964 9128 22976
rect 8527 22936 9128 22964
rect 8527 22933 8539 22936
rect 8481 22927 8539 22933
rect 9122 22924 9128 22936
rect 9180 22964 9186 22976
rect 9306 22964 9312 22976
rect 9180 22936 9312 22964
rect 9180 22924 9186 22936
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 9493 22967 9551 22973
rect 9493 22964 9505 22967
rect 9456 22936 9505 22964
rect 9456 22924 9462 22936
rect 9493 22933 9505 22936
rect 9539 22933 9551 22967
rect 10318 22964 10324 22976
rect 10279 22936 10324 22964
rect 9493 22927 9551 22933
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 10689 22967 10747 22973
rect 10689 22933 10701 22967
rect 10735 22964 10747 22967
rect 10778 22964 10784 22976
rect 10735 22936 10784 22964
rect 10735 22933 10747 22936
rect 10689 22927 10747 22933
rect 10778 22924 10784 22936
rect 10836 22964 10842 22976
rect 11146 22964 11152 22976
rect 10836 22936 11152 22964
rect 10836 22924 10842 22936
rect 11146 22924 11152 22936
rect 11204 22924 11210 22976
rect 11425 22967 11483 22973
rect 11425 22933 11437 22967
rect 11471 22964 11483 22967
rect 13446 22964 13452 22976
rect 11471 22936 13452 22964
rect 11471 22933 11483 22936
rect 11425 22927 11483 22933
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 13722 22964 13728 22976
rect 13683 22936 13728 22964
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 17678 22924 17684 22976
rect 17736 22964 17742 22976
rect 20254 22964 20260 22976
rect 17736 22936 20260 22964
rect 17736 22924 17742 22936
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 20916 22964 20944 23004
rect 21174 22964 21180 22976
rect 20916 22936 21180 22964
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 21634 22924 21640 22976
rect 21692 22964 21698 22976
rect 21729 22967 21787 22973
rect 21729 22964 21741 22967
rect 21692 22936 21741 22964
rect 21692 22924 21698 22936
rect 21729 22933 21741 22936
rect 21775 22933 21787 22967
rect 21836 22964 21864 23004
rect 22462 22992 22468 23004
rect 22520 22992 22526 23044
rect 22848 22964 22876 23063
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 23842 23100 23848 23112
rect 23803 23072 23848 23100
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23069 24087 23103
rect 24029 23063 24087 23069
rect 23658 22992 23664 23044
rect 23716 23032 23722 23044
rect 24044 23032 24072 23063
rect 24854 23060 24860 23112
rect 24912 23100 24918 23112
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 24912 23072 26249 23100
rect 24912 23060 24918 23072
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 26237 23063 26295 23069
rect 23716 23004 24072 23032
rect 23716 22992 23722 23004
rect 25130 22992 25136 23044
rect 25188 23032 25194 23044
rect 25317 23035 25375 23041
rect 25317 23032 25329 23035
rect 25188 23004 25329 23032
rect 25188 22992 25194 23004
rect 25317 23001 25329 23004
rect 25363 23001 25375 23035
rect 25317 22995 25375 23001
rect 21836 22936 22876 22964
rect 23937 22967 23995 22973
rect 21729 22927 21787 22933
rect 23937 22933 23949 22967
rect 23983 22964 23995 22967
rect 25038 22964 25044 22976
rect 23983 22936 25044 22964
rect 23983 22933 23995 22936
rect 23937 22927 23995 22933
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 25406 22964 25412 22976
rect 25367 22936 25412 22964
rect 25406 22924 25412 22936
rect 25464 22924 25470 22976
rect 25774 22964 25780 22976
rect 25735 22936 25780 22964
rect 25774 22924 25780 22936
rect 25832 22924 25838 22976
rect 26326 22964 26332 22976
rect 26287 22936 26332 22964
rect 26326 22924 26332 22936
rect 26384 22924 26390 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 2406 22720 2412 22772
rect 2464 22760 2470 22772
rect 5718 22760 5724 22772
rect 2464 22732 5724 22760
rect 2464 22720 2470 22732
rect 5718 22720 5724 22732
rect 5776 22720 5782 22772
rect 6270 22720 6276 22772
rect 6328 22760 6334 22772
rect 7466 22760 7472 22772
rect 6328 22732 7472 22760
rect 6328 22720 6334 22732
rect 7466 22720 7472 22732
rect 7524 22760 7530 22772
rect 7929 22763 7987 22769
rect 7929 22760 7941 22763
rect 7524 22732 7941 22760
rect 7524 22720 7530 22732
rect 7929 22729 7941 22732
rect 7975 22729 7987 22763
rect 7929 22723 7987 22729
rect 8481 22763 8539 22769
rect 8481 22729 8493 22763
rect 8527 22760 8539 22763
rect 9030 22760 9036 22772
rect 8527 22732 9036 22760
rect 8527 22729 8539 22732
rect 8481 22723 8539 22729
rect 2038 22652 2044 22704
rect 2096 22692 2102 22704
rect 4310 22695 4368 22701
rect 4310 22692 4322 22695
rect 2096 22664 4322 22692
rect 2096 22652 2102 22664
rect 4310 22661 4322 22664
rect 4356 22661 4368 22695
rect 4310 22655 4368 22661
rect 6638 22652 6644 22704
rect 6696 22692 6702 22704
rect 6794 22695 6852 22701
rect 6794 22692 6806 22695
rect 6696 22664 6806 22692
rect 6696 22652 6702 22664
rect 6794 22661 6806 22664
rect 6840 22661 6852 22695
rect 7944 22692 7972 22723
rect 9030 22720 9036 22732
rect 9088 22720 9094 22772
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9398 22760 9404 22772
rect 9180 22732 9404 22760
rect 9180 22720 9186 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 9493 22763 9551 22769
rect 9493 22729 9505 22763
rect 9539 22760 9551 22763
rect 9582 22760 9588 22772
rect 9539 22732 9588 22760
rect 9539 22729 9551 22732
rect 9493 22723 9551 22729
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 13357 22763 13415 22769
rect 9876 22732 11192 22760
rect 8570 22692 8576 22704
rect 7944 22664 8576 22692
rect 6794 22655 6852 22661
rect 8570 22652 8576 22664
rect 8628 22692 8634 22704
rect 8941 22695 8999 22701
rect 8941 22692 8953 22695
rect 8628 22664 8953 22692
rect 8628 22652 8634 22664
rect 8941 22661 8953 22664
rect 8987 22692 8999 22695
rect 9876 22692 9904 22732
rect 8987 22664 9904 22692
rect 9953 22695 10011 22701
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9953 22661 9965 22695
rect 9999 22692 10011 22695
rect 10594 22692 10600 22704
rect 9999 22664 10600 22692
rect 9999 22661 10011 22664
rect 9953 22655 10011 22661
rect 10594 22652 10600 22664
rect 10652 22652 10658 22704
rect 10962 22652 10968 22704
rect 11020 22692 11026 22704
rect 11020 22664 11065 22692
rect 11020 22652 11026 22664
rect 2222 22584 2228 22636
rect 2280 22624 2286 22636
rect 2409 22627 2467 22633
rect 2409 22624 2421 22627
rect 2280 22596 2421 22624
rect 2280 22584 2286 22596
rect 2409 22593 2421 22596
rect 2455 22593 2467 22627
rect 2409 22587 2467 22593
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22593 2651 22627
rect 2593 22587 2651 22593
rect 2685 22627 2743 22633
rect 2685 22593 2697 22627
rect 2731 22624 2743 22627
rect 3050 22624 3056 22636
rect 2731 22596 3056 22624
rect 2731 22593 2743 22596
rect 2685 22587 2743 22593
rect 2608 22556 2636 22587
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 3510 22624 3516 22636
rect 3471 22596 3516 22624
rect 3329 22587 3387 22593
rect 2774 22556 2780 22568
rect 2608 22528 2780 22556
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 3344 22556 3372 22587
rect 3510 22584 3516 22596
rect 3568 22584 3574 22636
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 3694 22624 3700 22636
rect 3651 22596 3700 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 3694 22584 3700 22596
rect 3752 22584 3758 22636
rect 4062 22624 4068 22636
rect 4023 22596 4068 22624
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 6454 22624 6460 22636
rect 4172 22596 6460 22624
rect 4172 22556 4200 22596
rect 6454 22584 6460 22596
rect 6512 22584 6518 22636
rect 9214 22624 9220 22636
rect 9175 22596 9220 22624
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 9306 22584 9312 22636
rect 9364 22624 9370 22636
rect 10134 22624 10140 22636
rect 9364 22596 9409 22624
rect 10095 22596 10140 22624
rect 9364 22584 9370 22596
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 10226 22584 10232 22636
rect 10284 22624 10290 22636
rect 10689 22627 10747 22633
rect 10284 22596 10329 22624
rect 10284 22584 10290 22596
rect 10689 22593 10701 22627
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 6546 22556 6552 22568
rect 3344 22528 4200 22556
rect 6507 22528 6552 22556
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 9398 22516 9404 22568
rect 9456 22556 9462 22568
rect 10704 22556 10732 22587
rect 10778 22584 10784 22636
rect 10836 22614 10842 22636
rect 10873 22627 10931 22633
rect 10873 22614 10885 22627
rect 10836 22593 10885 22614
rect 10919 22593 10931 22627
rect 10836 22587 10931 22593
rect 11077 22627 11135 22633
rect 11077 22593 11089 22627
rect 11123 22624 11135 22627
rect 11164 22624 11192 22732
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 13538 22760 13544 22772
rect 13403 22732 13544 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 14093 22763 14151 22769
rect 14093 22729 14105 22763
rect 14139 22760 14151 22763
rect 16390 22760 16396 22772
rect 14139 22732 16396 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 18230 22720 18236 22772
rect 18288 22760 18294 22772
rect 18782 22760 18788 22772
rect 18288 22732 18368 22760
rect 18288 22720 18294 22732
rect 13906 22652 13912 22704
rect 13964 22692 13970 22704
rect 16114 22692 16120 22704
rect 13964 22664 16120 22692
rect 13964 22652 13970 22664
rect 11123 22596 11192 22624
rect 11123 22593 11135 22596
rect 11077 22587 11135 22593
rect 10836 22586 10916 22587
rect 10836 22584 10842 22586
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 11698 22624 11704 22636
rect 11388 22596 11704 22624
rect 11388 22584 11394 22596
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 11790 22584 11796 22636
rect 11848 22624 11854 22636
rect 11848 22596 11893 22624
rect 11848 22584 11854 22596
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 13081 22627 13139 22633
rect 12032 22596 12077 22624
rect 12032 22584 12038 22596
rect 13081 22593 13093 22627
rect 13127 22593 13139 22627
rect 13262 22624 13268 22636
rect 13223 22596 13268 22624
rect 13081 22587 13139 22593
rect 9456 22528 10732 22556
rect 10965 22559 11023 22565
rect 9456 22516 9462 22528
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11606 22556 11612 22568
rect 11011 22528 11612 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 13096 22556 13124 22587
rect 13262 22584 13268 22596
rect 13320 22584 13326 22636
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 13630 22624 13636 22636
rect 13587 22596 13636 22624
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 13630 22584 13636 22596
rect 13688 22584 13694 22636
rect 13998 22624 14004 22636
rect 13959 22596 14004 22624
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 14292 22633 14320 22664
rect 16114 22652 16120 22664
rect 16172 22652 16178 22704
rect 18340 22701 18368 22732
rect 18432 22732 18788 22760
rect 18432 22701 18460 22732
rect 18782 22720 18788 22732
rect 18840 22760 18846 22772
rect 20165 22763 20223 22769
rect 18840 22732 19564 22760
rect 18840 22720 18846 22732
rect 18325 22695 18383 22701
rect 18325 22661 18337 22695
rect 18371 22661 18383 22695
rect 18325 22655 18383 22661
rect 18417 22695 18475 22701
rect 18417 22661 18429 22695
rect 18463 22661 18475 22695
rect 18417 22655 18475 22661
rect 18555 22695 18613 22701
rect 18555 22661 18567 22695
rect 18601 22692 18613 22695
rect 19426 22692 19432 22704
rect 18601 22664 19432 22692
rect 18601 22661 18613 22664
rect 18555 22655 18613 22661
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 14277 22627 14335 22633
rect 14277 22593 14289 22627
rect 14323 22593 14335 22627
rect 14277 22587 14335 22593
rect 15188 22627 15246 22633
rect 15188 22593 15200 22627
rect 15234 22624 15246 22627
rect 15562 22624 15568 22636
rect 15234 22596 15568 22624
rect 15234 22593 15246 22596
rect 15188 22587 15246 22593
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 17313 22627 17371 22633
rect 17313 22593 17325 22627
rect 17359 22624 17371 22627
rect 17862 22624 17868 22636
rect 17359 22596 17868 22624
rect 17359 22593 17371 22596
rect 17313 22587 17371 22593
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 19150 22624 19156 22636
rect 18279 22596 19156 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19536 22633 19564 22732
rect 20165 22729 20177 22763
rect 20211 22760 20223 22763
rect 20990 22760 20996 22772
rect 20211 22732 20996 22760
rect 20211 22729 20223 22732
rect 20165 22723 20223 22729
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 21266 22720 21272 22772
rect 21324 22760 21330 22772
rect 22005 22763 22063 22769
rect 22005 22760 22017 22763
rect 21324 22732 22017 22760
rect 21324 22720 21330 22732
rect 22005 22729 22017 22732
rect 22051 22729 22063 22763
rect 22005 22723 22063 22729
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 22925 22763 22983 22769
rect 22925 22760 22937 22763
rect 22612 22732 22937 22760
rect 22612 22720 22618 22732
rect 22925 22729 22937 22732
rect 22971 22760 22983 22763
rect 23382 22760 23388 22772
rect 22971 22732 23388 22760
rect 22971 22729 22983 22732
rect 22925 22723 22983 22729
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 19702 22652 19708 22704
rect 19760 22692 19766 22704
rect 20530 22692 20536 22704
rect 19760 22664 20536 22692
rect 19760 22652 19766 22664
rect 20530 22652 20536 22664
rect 20588 22652 20594 22704
rect 20622 22652 20628 22704
rect 20680 22692 20686 22704
rect 21085 22695 21143 22701
rect 21085 22692 21097 22695
rect 20680 22664 21097 22692
rect 20680 22652 20686 22664
rect 21085 22661 21097 22664
rect 21131 22661 21143 22695
rect 21085 22655 21143 22661
rect 21174 22652 21180 22704
rect 21232 22692 21238 22704
rect 25406 22692 25412 22704
rect 21232 22664 25412 22692
rect 21232 22652 21238 22664
rect 25406 22652 25412 22664
rect 25464 22692 25470 22704
rect 26050 22692 26056 22704
rect 25464 22664 26056 22692
rect 25464 22652 25470 22664
rect 26050 22652 26056 22664
rect 26108 22692 26114 22704
rect 26108 22664 26188 22692
rect 26108 22652 26114 22664
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 19260 22596 19349 22624
rect 13354 22556 13360 22568
rect 13096 22528 13360 22556
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 14918 22556 14924 22568
rect 14879 22528 14924 22556
rect 14918 22516 14924 22528
rect 14976 22516 14982 22568
rect 17402 22516 17408 22568
rect 17460 22556 17466 22568
rect 17497 22559 17555 22565
rect 17497 22556 17509 22559
rect 17460 22528 17509 22556
rect 17460 22516 17466 22528
rect 17497 22525 17509 22528
rect 17543 22525 17555 22559
rect 17497 22519 17555 22525
rect 17589 22559 17647 22565
rect 17589 22525 17601 22559
rect 17635 22556 17647 22559
rect 17678 22556 17684 22568
rect 17635 22528 17684 22556
rect 17635 22525 17647 22528
rect 17589 22519 17647 22525
rect 17678 22516 17684 22528
rect 17736 22516 17742 22568
rect 18690 22556 18696 22568
rect 18651 22528 18696 22556
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 1762 22488 1768 22500
rect 1675 22460 1768 22488
rect 1762 22448 1768 22460
rect 1820 22488 1826 22500
rect 3050 22488 3056 22500
rect 1820 22460 3056 22488
rect 1820 22448 1826 22460
rect 3050 22448 3056 22460
rect 3108 22448 3114 22500
rect 10229 22491 10287 22497
rect 10229 22457 10241 22491
rect 10275 22488 10287 22491
rect 11238 22488 11244 22500
rect 10275 22460 11244 22488
rect 10275 22457 10287 22460
rect 10229 22451 10287 22457
rect 11238 22448 11244 22460
rect 11296 22448 11302 22500
rect 11348 22460 12434 22488
rect 2225 22423 2283 22429
rect 2225 22389 2237 22423
rect 2271 22420 2283 22423
rect 2406 22420 2412 22432
rect 2271 22392 2412 22420
rect 2271 22389 2283 22392
rect 2225 22383 2283 22389
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 3142 22420 3148 22432
rect 3103 22392 3148 22420
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 5445 22423 5503 22429
rect 5445 22389 5457 22423
rect 5491 22420 5503 22423
rect 5718 22420 5724 22432
rect 5491 22392 5724 22420
rect 5491 22389 5503 22392
rect 5445 22383 5503 22389
rect 5718 22380 5724 22392
rect 5776 22380 5782 22432
rect 5902 22420 5908 22432
rect 5863 22392 5908 22420
rect 5902 22380 5908 22392
rect 5960 22380 5966 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 11348 22420 11376 22460
rect 12158 22420 12164 22432
rect 8352 22392 11376 22420
rect 12119 22392 12164 22420
rect 8352 22380 8358 22392
rect 12158 22380 12164 22392
rect 12216 22380 12222 22432
rect 12406 22420 12434 22460
rect 18230 22448 18236 22500
rect 18288 22488 18294 22500
rect 19260 22488 19288 22596
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22593 19579 22627
rect 19521 22587 19579 22593
rect 19889 22627 19947 22633
rect 19889 22593 19901 22627
rect 19935 22624 19947 22627
rect 22186 22624 22192 22636
rect 19935 22596 20668 22624
rect 22147 22596 22192 22624
rect 19935 22593 19947 22596
rect 19889 22587 19947 22593
rect 20162 22556 20168 22568
rect 20123 22528 20168 22556
rect 20162 22516 20168 22528
rect 20220 22516 20226 22568
rect 20640 22565 20668 22596
rect 22186 22584 22192 22596
rect 22244 22624 22250 22636
rect 22833 22627 22891 22633
rect 22833 22624 22845 22627
rect 22244 22596 22845 22624
rect 22244 22584 22250 22596
rect 22833 22593 22845 22596
rect 22879 22593 22891 22627
rect 22833 22587 22891 22593
rect 23017 22627 23075 22633
rect 23017 22593 23029 22627
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22624 23627 22627
rect 23750 22624 23756 22636
rect 23615 22596 23756 22624
rect 23615 22593 23627 22596
rect 23569 22587 23627 22593
rect 20625 22559 20683 22565
rect 20625 22525 20637 22559
rect 20671 22525 20683 22559
rect 20625 22519 20683 22525
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 22373 22559 22431 22565
rect 22373 22556 22385 22559
rect 21140 22528 22385 22556
rect 21140 22516 21146 22528
rect 22373 22525 22385 22528
rect 22419 22556 22431 22559
rect 23032 22556 23060 22587
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22624 23903 22627
rect 23934 22624 23940 22636
rect 23891 22596 23940 22624
rect 23891 22593 23903 22596
rect 23845 22587 23903 22593
rect 23934 22584 23940 22596
rect 23992 22624 23998 22636
rect 24486 22624 24492 22636
rect 23992 22596 24492 22624
rect 23992 22584 23998 22596
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 25225 22627 25283 22633
rect 25225 22593 25237 22627
rect 25271 22624 25283 22627
rect 25774 22624 25780 22636
rect 25271 22596 25780 22624
rect 25271 22593 25283 22596
rect 25225 22587 25283 22593
rect 25774 22584 25780 22596
rect 25832 22584 25838 22636
rect 26160 22633 26188 22664
rect 26145 22627 26203 22633
rect 26145 22593 26157 22627
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 23658 22556 23664 22568
rect 22419 22528 23060 22556
rect 23619 22528 23664 22556
rect 22419 22525 22431 22528
rect 22373 22519 22431 22525
rect 23658 22516 23664 22528
rect 23716 22516 23722 22568
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25409 22559 25467 22565
rect 25409 22556 25421 22559
rect 24912 22528 25421 22556
rect 24912 22516 24918 22528
rect 25409 22525 25421 22528
rect 25455 22525 25467 22559
rect 25409 22519 25467 22525
rect 25501 22559 25559 22565
rect 25501 22525 25513 22559
rect 25547 22556 25559 22559
rect 25590 22556 25596 22568
rect 25547 22528 25596 22556
rect 25547 22525 25559 22528
rect 25501 22519 25559 22525
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 26053 22559 26111 22565
rect 26053 22525 26065 22559
rect 26099 22556 26111 22559
rect 26234 22556 26240 22568
rect 26099 22528 26240 22556
rect 26099 22525 26111 22528
rect 26053 22519 26111 22525
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 18288 22460 19288 22488
rect 20717 22491 20775 22497
rect 18288 22448 18294 22460
rect 20717 22457 20729 22491
rect 20763 22457 20775 22491
rect 20717 22451 20775 22457
rect 13906 22420 13912 22432
rect 12406 22392 13912 22420
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 14461 22423 14519 22429
rect 14461 22389 14473 22423
rect 14507 22420 14519 22423
rect 15286 22420 15292 22432
rect 14507 22392 15292 22420
rect 14507 22389 14519 22392
rect 14461 22383 14519 22389
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 16298 22420 16304 22432
rect 16259 22392 16304 22420
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17129 22423 17187 22429
rect 17129 22420 17141 22423
rect 16816 22392 17141 22420
rect 16816 22380 16822 22392
rect 17129 22389 17141 22392
rect 17175 22389 17187 22423
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 17129 22383 17187 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 20732 22420 20760 22451
rect 19392 22392 20760 22420
rect 24029 22423 24087 22429
rect 19392 22380 19398 22392
rect 24029 22389 24041 22423
rect 24075 22420 24087 22423
rect 24578 22420 24584 22432
rect 24075 22392 24584 22420
rect 24075 22389 24087 22392
rect 24029 22383 24087 22389
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 24670 22380 24676 22432
rect 24728 22420 24734 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24728 22392 25053 22420
rect 24728 22380 24734 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 26418 22420 26424 22432
rect 26379 22392 26424 22420
rect 25041 22383 25099 22389
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 5997 22219 6055 22225
rect 5997 22185 6009 22219
rect 6043 22216 6055 22219
rect 6043 22188 9674 22216
rect 6043 22185 6055 22188
rect 5997 22179 6055 22185
rect 8386 22040 8392 22092
rect 8444 22080 8450 22092
rect 9214 22080 9220 22092
rect 8444 22052 9220 22080
rect 8444 22040 8450 22052
rect 9214 22040 9220 22052
rect 9272 22080 9278 22092
rect 9272 22052 9536 22080
rect 9272 22040 9278 22052
rect 2041 22015 2099 22021
rect 2041 21981 2053 22015
rect 2087 21981 2099 22015
rect 4062 22012 4068 22024
rect 4023 21984 4068 22012
rect 2041 21975 2099 21981
rect 2056 21876 2084 21975
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4332 22015 4390 22021
rect 4332 21981 4344 22015
rect 4378 22012 4390 22015
rect 4798 22012 4804 22024
rect 4378 21984 4804 22012
rect 4378 21981 4390 21984
rect 4332 21975 4390 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 22012 6515 22015
rect 6546 22012 6552 22024
rect 6503 21984 6552 22012
rect 6503 21981 6515 21984
rect 6457 21975 6515 21981
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 6730 22021 6736 22024
rect 6724 21975 6736 22021
rect 6788 22012 6794 22024
rect 6788 21984 6824 22012
rect 6730 21972 6736 21975
rect 6788 21972 6794 21984
rect 8570 21972 8576 22024
rect 8628 22012 8634 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8628 21984 9137 22012
rect 8628 21972 8634 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9306 22012 9312 22024
rect 9267 21984 9312 22012
rect 9125 21975 9183 21981
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 9508 22021 9536 22052
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 2308 21947 2366 21953
rect 2308 21913 2320 21947
rect 2354 21944 2366 21947
rect 2406 21944 2412 21956
rect 2354 21916 2412 21944
rect 2354 21913 2366 21916
rect 2308 21907 2366 21913
rect 2406 21904 2412 21916
rect 2464 21904 2470 21956
rect 2866 21944 2872 21956
rect 2700 21916 2872 21944
rect 2700 21876 2728 21916
rect 2866 21904 2872 21916
rect 2924 21904 2930 21956
rect 9398 21944 9404 21956
rect 7852 21916 9404 21944
rect 2056 21848 2728 21876
rect 2774 21836 2780 21888
rect 2832 21876 2838 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 2832 21848 3433 21876
rect 2832 21836 2838 21848
rect 3421 21845 3433 21848
rect 3467 21876 3479 21879
rect 5166 21876 5172 21888
rect 3467 21848 5172 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 5442 21876 5448 21888
rect 5403 21848 5448 21876
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 7852 21885 7880 21916
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 9646 21944 9674 22188
rect 11238 22176 11244 22228
rect 11296 22216 11302 22228
rect 12066 22216 12072 22228
rect 11296 22188 12072 22216
rect 11296 22176 11302 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 12710 22216 12716 22228
rect 12671 22188 12716 22216
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 13725 22219 13783 22225
rect 13725 22185 13737 22219
rect 13771 22216 13783 22219
rect 14550 22216 14556 22228
rect 13771 22188 14556 22216
rect 13771 22185 13783 22188
rect 13725 22179 13783 22185
rect 14550 22176 14556 22188
rect 14608 22176 14614 22228
rect 16114 22176 16120 22228
rect 16172 22216 16178 22228
rect 16172 22188 16574 22216
rect 16172 22176 16178 22188
rect 11698 22108 11704 22160
rect 11756 22148 11762 22160
rect 13998 22148 14004 22160
rect 11756 22120 14004 22148
rect 11756 22108 11762 22120
rect 13998 22108 14004 22120
rect 14056 22108 14062 22160
rect 16390 22148 16396 22160
rect 16351 22120 16396 22148
rect 16390 22108 16396 22120
rect 16448 22108 16454 22160
rect 10962 22040 10968 22092
rect 11020 22080 11026 22092
rect 11790 22080 11796 22092
rect 11020 22052 11796 22080
rect 11020 22040 11026 22052
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12434 22040 12440 22092
rect 12492 22080 12498 22092
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 12492 22052 12725 22080
rect 12492 22040 12498 22052
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 12802 22040 12808 22092
rect 12860 22080 12866 22092
rect 14642 22080 14648 22092
rect 12860 22052 14648 22080
rect 12860 22040 12866 22052
rect 12618 22012 12624 22024
rect 12579 21984 12624 22012
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 13446 21972 13452 22024
rect 13504 22012 13510 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 13504 21984 13553 22012
rect 13504 21972 13510 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 14384 22021 14412 22052
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 16546 22080 16574 22188
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18233 22219 18291 22225
rect 18233 22216 18245 22219
rect 18196 22188 18245 22216
rect 18196 22176 18202 22188
rect 18233 22185 18245 22188
rect 18279 22185 18291 22219
rect 19426 22216 19432 22228
rect 19387 22188 19432 22216
rect 18233 22179 18291 22185
rect 19426 22176 19432 22188
rect 19484 22176 19490 22228
rect 20622 22216 20628 22228
rect 19720 22188 20628 22216
rect 19150 22108 19156 22160
rect 19208 22148 19214 22160
rect 19518 22148 19524 22160
rect 19208 22120 19524 22148
rect 19208 22108 19214 22120
rect 19518 22108 19524 22120
rect 19576 22108 19582 22160
rect 19610 22108 19616 22160
rect 19668 22108 19674 22160
rect 19720 22157 19748 22188
rect 20622 22176 20628 22188
rect 20680 22216 20686 22228
rect 20717 22219 20775 22225
rect 20717 22216 20729 22219
rect 20680 22188 20729 22216
rect 20680 22176 20686 22188
rect 20717 22185 20729 22188
rect 20763 22185 20775 22219
rect 20717 22179 20775 22185
rect 21269 22219 21327 22225
rect 21269 22185 21281 22219
rect 21315 22216 21327 22219
rect 21910 22216 21916 22228
rect 21315 22188 21916 22216
rect 21315 22185 21327 22188
rect 21269 22179 21327 22185
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 22005 22219 22063 22225
rect 22005 22185 22017 22219
rect 22051 22216 22063 22219
rect 22186 22216 22192 22228
rect 22051 22188 22192 22216
rect 22051 22185 22063 22188
rect 22005 22179 22063 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 23750 22216 23756 22228
rect 23711 22188 23756 22216
rect 23750 22176 23756 22188
rect 23808 22176 23814 22228
rect 24854 22176 24860 22228
rect 24912 22216 24918 22228
rect 25038 22216 25044 22228
rect 24912 22188 25044 22216
rect 24912 22176 24918 22188
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 19705 22151 19763 22157
rect 19705 22117 19717 22151
rect 19751 22117 19763 22151
rect 19705 22111 19763 22117
rect 20254 22108 20260 22160
rect 20312 22148 20318 22160
rect 22094 22148 22100 22160
rect 20312 22120 22100 22148
rect 20312 22108 20318 22120
rect 16546 22052 16988 22080
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 13780 21984 14289 22012
rect 13780 21972 13786 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 14918 22012 14924 22024
rect 14792 21984 14924 22012
rect 14792 21972 14798 21984
rect 14918 21972 14924 21984
rect 14976 22012 14982 22024
rect 15286 22021 15292 22024
rect 15013 22015 15071 22021
rect 15013 22012 15025 22015
rect 14976 21984 15025 22012
rect 14976 21972 14982 21984
rect 15013 21981 15025 21984
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 15280 21975 15292 22021
rect 15344 22012 15350 22024
rect 16850 22012 16856 22024
rect 15344 21984 15380 22012
rect 16811 21984 16856 22012
rect 15286 21972 15292 21975
rect 15344 21972 15350 21984
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 16960 22012 16988 22052
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 19628 22080 19656 22108
rect 19392 22052 19656 22080
rect 19392 22040 19398 22052
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 20220 22052 21220 22080
rect 20220 22040 20226 22052
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 16960 21984 18705 22012
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 18693 21975 18751 21981
rect 19352 21984 19625 22012
rect 19352 21956 19380 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19794 22012 19800 22024
rect 19755 21984 19800 22012
rect 19613 21975 19671 21981
rect 19794 21972 19800 21984
rect 19852 21972 19858 22024
rect 19886 21972 19892 22024
rect 19944 22012 19950 22024
rect 20073 22015 20131 22021
rect 19944 21984 19989 22012
rect 19944 21972 19950 21984
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20530 22012 20536 22024
rect 20491 21984 20536 22012
rect 20073 21975 20131 21981
rect 10410 21944 10416 21956
rect 9646 21916 10416 21944
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 12161 21947 12219 21953
rect 12161 21913 12173 21947
rect 12207 21944 12219 21947
rect 12526 21944 12532 21956
rect 12207 21916 12532 21944
rect 12207 21913 12219 21916
rect 12161 21907 12219 21913
rect 12526 21904 12532 21916
rect 12584 21904 12590 21956
rect 14090 21904 14096 21956
rect 14148 21944 14154 21956
rect 14553 21947 14611 21953
rect 14553 21944 14565 21947
rect 14148 21916 14565 21944
rect 14148 21904 14154 21916
rect 14553 21913 14565 21916
rect 14599 21913 14611 21947
rect 14553 21907 14611 21913
rect 17120 21947 17178 21953
rect 17120 21913 17132 21947
rect 17166 21944 17178 21947
rect 17862 21944 17868 21956
rect 17166 21916 17868 21944
rect 17166 21913 17178 21916
rect 17120 21907 17178 21913
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 19334 21904 19340 21956
rect 19392 21904 19398 21956
rect 7837 21879 7895 21885
rect 7837 21845 7849 21879
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21876 8631 21879
rect 8846 21876 8852 21888
rect 8619 21848 8852 21876
rect 8619 21845 8631 21848
rect 8573 21839 8631 21845
rect 8846 21836 8852 21848
rect 8904 21836 8910 21888
rect 9674 21876 9680 21888
rect 9635 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 11054 21876 11060 21888
rect 10919 21848 11060 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 12986 21876 12992 21888
rect 12947 21848 12992 21876
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 14458 21885 14464 21888
rect 14454 21839 14464 21885
rect 14516 21876 14522 21888
rect 14516 21848 14554 21876
rect 14458 21836 14464 21839
rect 14516 21836 14522 21848
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 20088 21876 20116 21975
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20622 21972 20628 22024
rect 20680 21972 20686 22024
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 20806 22012 20812 22024
rect 20763 21984 20812 22012
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 20806 21972 20812 21984
rect 20864 22012 20870 22024
rect 21082 22012 21088 22024
rect 20864 21984 21088 22012
rect 20864 21972 20870 21984
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 21192 22021 21220 22052
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 21981 21235 22015
rect 21358 22012 21364 22024
rect 21319 21984 21364 22012
rect 21177 21975 21235 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 21836 22021 21864 22120
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 26418 22108 26424 22160
rect 26476 22148 26482 22160
rect 26476 22120 26556 22148
rect 26476 22108 26482 22120
rect 23566 22040 23572 22092
rect 23624 22080 23630 22092
rect 23753 22083 23811 22089
rect 23753 22080 23765 22083
rect 23624 22052 23765 22080
rect 23624 22040 23630 22052
rect 23753 22049 23765 22052
rect 23799 22080 23811 22083
rect 23934 22080 23940 22092
rect 23799 22052 23940 22080
rect 23799 22049 23811 22052
rect 23753 22043 23811 22049
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 26528 22089 26556 22120
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22080 26571 22083
rect 26559 22052 26593 22080
rect 26559 22049 26571 22052
rect 26513 22043 26571 22049
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 21981 21879 22015
rect 21821 21975 21879 21981
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 21981 22063 22015
rect 23658 22012 23664 22024
rect 23619 21984 23664 22012
rect 22005 21975 22063 21981
rect 20346 21904 20352 21956
rect 20404 21944 20410 21956
rect 20640 21944 20668 21972
rect 20404 21916 20668 21944
rect 20404 21904 20410 21916
rect 21910 21904 21916 21956
rect 21968 21944 21974 21956
rect 22014 21944 22042 21975
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24674 22015 24732 22021
rect 24674 21981 24686 22015
rect 24720 21981 24732 22015
rect 24674 21975 24732 21981
rect 21968 21916 22042 21944
rect 21968 21904 21974 21916
rect 20622 21876 20628 21888
rect 17644 21848 20628 21876
rect 17644 21836 17650 21848
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 22462 21876 22468 21888
rect 22423 21848 22468 21876
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 24029 21879 24087 21885
rect 24029 21845 24041 21879
rect 24075 21876 24087 21879
rect 24688 21876 24716 21975
rect 25038 21972 25044 22024
rect 25096 22021 25102 22024
rect 25096 22012 25104 22021
rect 25685 22015 25743 22021
rect 25096 21984 25141 22012
rect 25096 21975 25104 21984
rect 25685 21981 25697 22015
rect 25731 22012 25743 22015
rect 25774 22012 25780 22024
rect 25731 21984 25780 22012
rect 25731 21981 25743 21984
rect 25685 21975 25743 21981
rect 25096 21972 25102 21975
rect 25774 21972 25780 21984
rect 25832 21972 25838 22024
rect 25869 22015 25927 22021
rect 25869 21981 25881 22015
rect 25915 22012 25927 22015
rect 26326 22012 26332 22024
rect 25915 21984 26332 22012
rect 25915 21981 25927 21984
rect 25869 21975 25927 21981
rect 26326 21972 26332 21984
rect 26384 22012 26390 22024
rect 26697 22015 26755 22021
rect 26697 22012 26709 22015
rect 26384 21984 26709 22012
rect 26384 21972 26390 21984
rect 26697 21981 26709 21984
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 24854 21944 24860 21956
rect 24815 21916 24860 21944
rect 24854 21904 24860 21916
rect 24912 21904 24918 21956
rect 24949 21947 25007 21953
rect 24949 21913 24961 21947
rect 24995 21944 25007 21947
rect 25590 21944 25596 21956
rect 24995 21916 25596 21944
rect 24995 21913 25007 21916
rect 24949 21907 25007 21913
rect 25590 21904 25596 21916
rect 25648 21904 25654 21956
rect 24075 21848 24716 21876
rect 24075 21845 24087 21848
rect 24029 21839 24087 21845
rect 24762 21836 24768 21888
rect 24820 21876 24826 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 24820 21848 25237 21876
rect 24820 21836 24826 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 25777 21879 25835 21885
rect 25777 21845 25789 21879
rect 25823 21876 25835 21879
rect 26605 21879 26663 21885
rect 26605 21876 26617 21879
rect 25823 21848 26617 21876
rect 25823 21845 25835 21848
rect 25777 21839 25835 21845
rect 26605 21845 26617 21848
rect 26651 21845 26663 21879
rect 26605 21839 26663 21845
rect 27065 21879 27123 21885
rect 27065 21845 27077 21879
rect 27111 21876 27123 21879
rect 27154 21876 27160 21888
rect 27111 21848 27160 21876
rect 27111 21845 27123 21848
rect 27065 21839 27123 21845
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 3418 21672 3424 21684
rect 2271 21644 3424 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 9306 21672 9312 21684
rect 9267 21644 9312 21672
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 11146 21672 11152 21684
rect 11107 21644 11152 21672
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 11790 21632 11796 21684
rect 11848 21672 11854 21684
rect 13081 21675 13139 21681
rect 13081 21672 13093 21675
rect 11848 21644 13093 21672
rect 11848 21632 11854 21644
rect 13081 21641 13093 21644
rect 13127 21641 13139 21675
rect 14090 21672 14096 21684
rect 14051 21644 14096 21672
rect 13081 21635 13139 21641
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 15562 21672 15568 21684
rect 15523 21644 15568 21672
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 15933 21675 15991 21681
rect 15933 21641 15945 21675
rect 15979 21672 15991 21675
rect 16298 21672 16304 21684
rect 15979 21644 16304 21672
rect 15979 21641 15991 21644
rect 15933 21635 15991 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 18230 21632 18236 21684
rect 18288 21672 18294 21684
rect 19061 21675 19119 21681
rect 19061 21672 19073 21675
rect 18288 21644 19073 21672
rect 18288 21632 18294 21644
rect 19061 21641 19073 21644
rect 19107 21641 19119 21675
rect 19061 21635 19119 21641
rect 19245 21675 19303 21681
rect 19245 21641 19257 21675
rect 19291 21672 19303 21675
rect 19794 21672 19800 21684
rect 19291 21644 19800 21672
rect 19291 21641 19303 21644
rect 19245 21635 19303 21641
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 19886 21632 19892 21684
rect 19944 21672 19950 21684
rect 23474 21672 23480 21684
rect 19944 21644 22876 21672
rect 19944 21632 19950 21644
rect 3145 21607 3203 21613
rect 3145 21573 3157 21607
rect 3191 21604 3203 21607
rect 3510 21604 3516 21616
rect 3191 21576 3516 21604
rect 3191 21573 3203 21576
rect 3145 21567 3203 21573
rect 3510 21564 3516 21576
rect 3568 21564 3574 21616
rect 5074 21564 5080 21616
rect 5132 21604 5138 21616
rect 10036 21607 10094 21613
rect 5132 21576 7512 21604
rect 5132 21564 5138 21576
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21536 2099 21539
rect 2130 21536 2136 21548
rect 2087 21508 2136 21536
rect 2087 21505 2099 21508
rect 2041 21499 2099 21505
rect 2130 21496 2136 21508
rect 2188 21496 2194 21548
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21536 3019 21539
rect 3050 21536 3056 21548
rect 3007 21508 3056 21536
rect 3007 21505 3019 21508
rect 2961 21499 3019 21505
rect 2332 21468 2360 21499
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3237 21539 3295 21545
rect 3237 21505 3249 21539
rect 3283 21536 3295 21539
rect 3694 21536 3700 21548
rect 3283 21508 3700 21536
rect 3283 21505 3295 21508
rect 3237 21499 3295 21505
rect 3252 21468 3280 21499
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 7098 21536 7104 21548
rect 5859 21508 7104 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 7193 21539 7251 21545
rect 7193 21505 7205 21539
rect 7239 21505 7251 21539
rect 7374 21536 7380 21548
rect 7335 21508 7380 21536
rect 7193 21499 7251 21505
rect 2332 21440 3280 21468
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 7208 21468 7236 21499
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 7484 21545 7512 21576
rect 7944 21576 9812 21604
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 7558 21536 7564 21548
rect 7515 21508 7564 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 7064 21440 7236 21468
rect 7064 21428 7070 21440
rect 1857 21335 1915 21341
rect 1857 21301 1869 21335
rect 1903 21332 1915 21335
rect 2314 21332 2320 21344
rect 1903 21304 2320 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 4338 21332 4344 21344
rect 2832 21304 2877 21332
rect 4299 21304 4344 21332
rect 2832 21292 2838 21304
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 7006 21332 7012 21344
rect 6967 21304 7012 21332
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7208 21332 7236 21440
rect 7742 21428 7748 21480
rect 7800 21468 7806 21480
rect 7944 21477 7972 21576
rect 8018 21496 8024 21548
rect 8076 21536 8082 21548
rect 9784 21545 9812 21576
rect 10036 21573 10048 21607
rect 10082 21604 10094 21607
rect 10318 21604 10324 21616
rect 10082 21576 10324 21604
rect 10082 21573 10094 21576
rect 10036 21567 10094 21573
rect 10318 21564 10324 21576
rect 10376 21564 10382 21616
rect 11968 21607 12026 21613
rect 11968 21573 11980 21607
rect 12014 21604 12026 21607
rect 12158 21604 12164 21616
rect 12014 21576 12164 21604
rect 12014 21573 12026 21576
rect 11968 21567 12026 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 13630 21564 13636 21616
rect 13688 21604 13694 21616
rect 13725 21607 13783 21613
rect 13725 21604 13737 21607
rect 13688 21576 13737 21604
rect 13688 21564 13694 21576
rect 13725 21573 13737 21576
rect 13771 21573 13783 21607
rect 16942 21604 16948 21616
rect 13725 21567 13783 21573
rect 14844 21576 16948 21604
rect 8185 21539 8243 21545
rect 8185 21536 8197 21539
rect 8076 21508 8197 21536
rect 8076 21496 8082 21508
rect 8185 21505 8197 21508
rect 8231 21505 8243 21539
rect 8185 21499 8243 21505
rect 9769 21539 9827 21545
rect 9769 21505 9781 21539
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 14182 21536 14188 21548
rect 13955 21508 14188 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 14844 21545 14872 21576
rect 16942 21564 16948 21576
rect 17000 21564 17006 21616
rect 17120 21607 17178 21613
rect 17120 21573 17132 21607
rect 17166 21604 17178 21607
rect 17954 21604 17960 21616
rect 17166 21576 17960 21604
rect 17166 21573 17178 21576
rect 17120 21567 17178 21573
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 19518 21564 19524 21616
rect 19576 21604 19582 21616
rect 19705 21607 19763 21613
rect 19705 21604 19717 21607
rect 19576 21576 19717 21604
rect 19576 21564 19582 21576
rect 19705 21573 19717 21576
rect 19751 21573 19763 21607
rect 20162 21604 20168 21616
rect 20123 21576 20168 21604
rect 19705 21567 19763 21573
rect 20162 21564 20168 21576
rect 20220 21604 20226 21616
rect 20714 21604 20720 21616
rect 20220 21576 20720 21604
rect 20220 21564 20226 21576
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 21358 21564 21364 21616
rect 21416 21604 21422 21616
rect 21416 21576 22784 21604
rect 21416 21564 21422 21576
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 15562 21536 15568 21548
rect 15059 21508 15568 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7800 21440 7941 21468
rect 7800 21428 7806 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 11701 21471 11759 21477
rect 11701 21468 11713 21471
rect 11020 21440 11713 21468
rect 11020 21428 11026 21440
rect 11701 21437 11713 21440
rect 11747 21437 11759 21471
rect 11701 21431 11759 21437
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 14844 21468 14872 21499
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 15746 21536 15752 21548
rect 15707 21508 15752 21536
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16022 21536 16028 21548
rect 15896 21508 16028 21536
rect 15896 21496 15902 21508
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 17460 21508 18705 21536
rect 17460 21496 17466 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19889 21539 19947 21545
rect 19889 21536 19901 21539
rect 19484 21508 19901 21536
rect 19484 21496 19490 21508
rect 19889 21505 19901 21508
rect 19935 21505 19947 21539
rect 19889 21499 19947 21505
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21505 20039 21539
rect 20622 21536 20628 21548
rect 20583 21508 20628 21536
rect 19981 21499 20039 21505
rect 13596 21440 14872 21468
rect 15105 21471 15163 21477
rect 13596 21428 13602 21440
rect 15105 21437 15117 21471
rect 15151 21468 15163 21471
rect 16666 21468 16672 21480
rect 15151 21440 16672 21468
rect 15151 21437 15163 21440
rect 15105 21431 15163 21437
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 16850 21468 16856 21480
rect 16811 21440 16856 21468
rect 16850 21428 16856 21440
rect 16908 21428 16914 21480
rect 19242 21468 19248 21480
rect 18248 21440 19248 21468
rect 18248 21409 18276 21440
rect 19242 21428 19248 21440
rect 19300 21468 19306 21480
rect 19797 21471 19855 21477
rect 19797 21468 19809 21471
rect 19300 21440 19809 21468
rect 19300 21428 19306 21440
rect 19797 21437 19809 21440
rect 19843 21437 19855 21471
rect 19797 21431 19855 21437
rect 18233 21403 18291 21409
rect 18233 21369 18245 21403
rect 18279 21369 18291 21403
rect 18233 21363 18291 21369
rect 18340 21372 19288 21400
rect 10042 21332 10048 21344
rect 7208 21304 10048 21332
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 12986 21292 12992 21344
rect 13044 21332 13050 21344
rect 18340 21332 18368 21372
rect 13044 21304 18368 21332
rect 19061 21335 19119 21341
rect 13044 21292 13050 21304
rect 19061 21301 19073 21335
rect 19107 21332 19119 21335
rect 19150 21332 19156 21344
rect 19107 21304 19156 21332
rect 19107 21301 19119 21304
rect 19061 21295 19119 21301
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 19260 21332 19288 21372
rect 19334 21360 19340 21412
rect 19392 21400 19398 21412
rect 19996 21400 20024 21499
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 19392 21372 20024 21400
rect 19392 21360 19398 21372
rect 20070 21360 20076 21412
rect 20128 21400 20134 21412
rect 22462 21400 22468 21412
rect 20128 21372 22468 21400
rect 20128 21360 20134 21372
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 19978 21332 19984 21344
rect 19260 21304 19984 21332
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 21269 21335 21327 21341
rect 21269 21332 21281 21335
rect 20680 21304 21281 21332
rect 20680 21292 20686 21304
rect 21269 21301 21281 21304
rect 21315 21332 21327 21335
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21315 21304 22017 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22756 21332 22784 21576
rect 22848 21545 22876 21644
rect 22940 21644 23480 21672
rect 22940 21545 22968 21644
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24762 21672 24768 21684
rect 24443 21644 24768 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 25130 21632 25136 21684
rect 25188 21672 25194 21684
rect 26421 21675 26479 21681
rect 26421 21672 26433 21675
rect 25188 21644 26433 21672
rect 25188 21632 25194 21644
rect 26421 21641 26433 21644
rect 26467 21641 26479 21675
rect 26421 21635 26479 21641
rect 23385 21607 23443 21613
rect 23385 21573 23397 21607
rect 23431 21604 23443 21607
rect 23431 21576 26556 21604
rect 23431 21573 23443 21576
rect 23385 21567 23443 21573
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 23106 21536 23112 21548
rect 23067 21508 23112 21536
rect 22925 21499 22983 21505
rect 22848 21468 22876 21499
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21536 23259 21539
rect 23842 21536 23848 21548
rect 23247 21508 23848 21536
rect 23247 21505 23259 21508
rect 23201 21499 23259 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 26528 21545 26556 21576
rect 25409 21539 25467 21545
rect 25409 21536 25421 21539
rect 25188 21508 25421 21536
rect 25188 21496 25194 21508
rect 25409 21505 25421 21508
rect 25455 21505 25467 21539
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 25409 21499 25467 21505
rect 25516 21508 26249 21536
rect 23014 21468 23020 21480
rect 22848 21440 23020 21468
rect 23014 21428 23020 21440
rect 23072 21428 23078 21480
rect 24670 21468 24676 21480
rect 24631 21440 24676 21468
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 24765 21471 24823 21477
rect 24765 21437 24777 21471
rect 24811 21468 24823 21471
rect 25317 21471 25375 21477
rect 25317 21468 25329 21471
rect 24811 21440 25329 21468
rect 24811 21437 24823 21440
rect 24765 21431 24823 21437
rect 25317 21437 25329 21440
rect 25363 21437 25375 21471
rect 25317 21431 25375 21437
rect 23658 21360 23664 21412
rect 23716 21400 23722 21412
rect 24581 21403 24639 21409
rect 24581 21400 24593 21403
rect 23716 21372 24593 21400
rect 23716 21360 23722 21372
rect 24581 21369 24593 21372
rect 24627 21400 24639 21403
rect 25516 21400 25544 21508
rect 26237 21505 26249 21508
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 26513 21539 26571 21545
rect 26513 21505 26525 21539
rect 26559 21505 26571 21539
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 26513 21499 26571 21505
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27246 21496 27252 21548
rect 27304 21536 27310 21548
rect 27341 21539 27399 21545
rect 27341 21536 27353 21539
rect 27304 21508 27353 21536
rect 27304 21496 27310 21508
rect 27341 21505 27353 21508
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 26234 21400 26240 21412
rect 24627 21372 25544 21400
rect 26195 21372 26240 21400
rect 24627 21369 24639 21372
rect 24581 21363 24639 21369
rect 26234 21360 26240 21372
rect 26292 21360 26298 21412
rect 25590 21332 25596 21344
rect 22756 21304 25596 21332
rect 22005 21295 22063 21301
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 25685 21335 25743 21341
rect 25685 21301 25697 21335
rect 25731 21332 25743 21335
rect 26326 21332 26332 21344
rect 25731 21304 26332 21332
rect 25731 21301 25743 21304
rect 25685 21295 25743 21301
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 27249 21335 27307 21341
rect 27249 21301 27261 21335
rect 27295 21332 27307 21335
rect 27706 21332 27712 21344
rect 27295 21304 27712 21332
rect 27295 21301 27307 21304
rect 27249 21295 27307 21301
rect 27706 21292 27712 21304
rect 27764 21292 27770 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 6546 21128 6552 21140
rect 6507 21100 6552 21128
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 7098 21088 7104 21140
rect 7156 21128 7162 21140
rect 7469 21131 7527 21137
rect 7469 21128 7481 21131
rect 7156 21100 7481 21128
rect 7156 21088 7162 21100
rect 7469 21097 7481 21100
rect 7515 21097 7527 21131
rect 7469 21091 7527 21097
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 13265 21131 13323 21137
rect 13265 21128 13277 21131
rect 13044 21100 13277 21128
rect 13044 21088 13050 21100
rect 13265 21097 13277 21100
rect 13311 21097 13323 21131
rect 13446 21128 13452 21140
rect 13407 21100 13452 21128
rect 13265 21091 13323 21097
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 8662 21060 8668 21072
rect 7248 21032 8668 21060
rect 7248 21020 7254 21032
rect 8662 21020 8668 21032
rect 8720 21020 8726 21072
rect 13280 21060 13308 21091
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 16850 21088 16856 21140
rect 16908 21128 16914 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 16908 21100 16957 21128
rect 16908 21088 16914 21100
rect 16945 21097 16957 21100
rect 16991 21097 17003 21131
rect 16945 21091 17003 21097
rect 17034 21088 17040 21140
rect 17092 21128 17098 21140
rect 19886 21128 19892 21140
rect 17092 21100 19892 21128
rect 17092 21088 17098 21100
rect 19886 21088 19892 21100
rect 19944 21088 19950 21140
rect 23658 21128 23664 21140
rect 23619 21100 23664 21128
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 24670 21088 24676 21140
rect 24728 21128 24734 21140
rect 24949 21131 25007 21137
rect 24949 21128 24961 21131
rect 24728 21100 24961 21128
rect 24728 21088 24734 21100
rect 24949 21097 24961 21100
rect 24995 21097 25007 21131
rect 26973 21131 27031 21137
rect 24949 21091 25007 21097
rect 25332 21100 25544 21128
rect 13814 21060 13820 21072
rect 13280 21032 13820 21060
rect 13814 21020 13820 21032
rect 13872 21020 13878 21072
rect 15746 21060 15752 21072
rect 14568 21032 15752 21060
rect 8478 20992 8484 21004
rect 8128 20964 8484 20992
rect 5258 20924 5264 20936
rect 5219 20896 5264 20924
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 8128 20933 8156 20964
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 8573 20995 8631 21001
rect 8573 20961 8585 20995
rect 8619 20992 8631 20995
rect 10226 20992 10232 21004
rect 8619 20964 10232 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 14568 20992 14596 21032
rect 15746 21020 15752 21032
rect 15804 21060 15810 21072
rect 16206 21060 16212 21072
rect 15804 21032 16212 21060
rect 15804 21020 15810 21032
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 21542 21060 21548 21072
rect 16356 21032 21548 21060
rect 16356 21020 16362 21032
rect 21542 21020 21548 21032
rect 21600 21060 21606 21072
rect 25332 21060 25360 21100
rect 21600 21032 21772 21060
rect 21600 21020 21606 21032
rect 12406 20964 14596 20992
rect 7653 20927 7711 20933
rect 7653 20924 7665 20927
rect 7340 20896 7665 20924
rect 7340 20884 7346 20896
rect 7653 20893 7665 20896
rect 7699 20893 7711 20927
rect 7653 20887 7711 20893
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20920 8447 20927
rect 8435 20893 8464 20920
rect 8389 20887 8464 20893
rect 1581 20859 1639 20865
rect 1581 20825 1593 20859
rect 1627 20856 1639 20859
rect 2958 20856 2964 20868
rect 1627 20828 2964 20856
rect 1627 20825 1639 20828
rect 1581 20819 1639 20825
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 4706 20856 4712 20868
rect 4667 20828 4712 20856
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 8436 20856 8464 20887
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 8720 20896 10425 20924
rect 8720 20884 8726 20896
rect 10413 20893 10425 20896
rect 10459 20924 10471 20927
rect 11054 20924 11060 20936
rect 10459 20896 11060 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 8570 20856 8576 20868
rect 8436 20828 8576 20856
rect 8570 20816 8576 20828
rect 8628 20856 8634 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 8628 20828 9229 20856
rect 8628 20816 8634 20828
rect 9217 20825 9229 20828
rect 9263 20856 9275 20859
rect 12406 20856 12434 20964
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 14921 20995 14979 21001
rect 14921 20992 14933 20995
rect 14700 20964 14933 20992
rect 14700 20952 14706 20964
rect 14921 20961 14933 20964
rect 14967 20961 14979 20995
rect 14921 20955 14979 20961
rect 17218 20952 17224 21004
rect 17276 20992 17282 21004
rect 20070 20992 20076 21004
rect 17276 20964 20076 20992
rect 17276 20952 17282 20964
rect 20070 20952 20076 20964
rect 20128 20952 20134 21004
rect 21744 21001 21772 21032
rect 23216 21032 25360 21060
rect 25409 21063 25467 21069
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20961 21787 20995
rect 21729 20955 21787 20961
rect 21640 20936 21692 20942
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 14240 20896 14473 20924
rect 14240 20884 14246 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 14829 20927 14887 20933
rect 14608 20896 14653 20924
rect 14608 20884 14614 20896
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 18138 20924 18144 20936
rect 14875 20896 18144 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 18138 20884 18144 20896
rect 18196 20884 18202 20936
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 18288 20896 18337 20924
rect 18288 20884 18294 20896
rect 18325 20893 18337 20896
rect 18371 20924 18383 20927
rect 20349 20927 20407 20933
rect 20349 20924 20361 20927
rect 18371 20896 20361 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 20349 20893 20361 20896
rect 20395 20924 20407 20927
rect 20530 20924 20536 20936
rect 20395 20896 20536 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 23014 20924 23020 20936
rect 22975 20896 23020 20924
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 23216 20933 23244 21032
rect 25409 21029 25421 21063
rect 25455 21029 25467 21063
rect 25409 21023 25467 21029
rect 23382 20992 23388 21004
rect 23343 20964 23388 20992
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23566 20952 23572 21004
rect 23624 20992 23630 21004
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 23624 20964 24593 20992
rect 23624 20952 23630 20964
rect 24581 20961 24593 20964
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 23164 20896 23213 20924
rect 23164 20884 23170 20896
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 23290 20884 23296 20936
rect 23348 20924 23354 20936
rect 23348 20896 23393 20924
rect 23348 20884 23354 20896
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 24765 20927 24823 20933
rect 23532 20896 23577 20924
rect 23532 20884 23538 20896
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24854 20924 24860 20936
rect 24811 20896 24860 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 24854 20884 24860 20896
rect 24912 20924 24918 20936
rect 25424 20924 25452 21023
rect 25516 20924 25544 21100
rect 26973 21097 26985 21131
rect 27019 21128 27031 21131
rect 27154 21128 27160 21140
rect 27019 21100 27160 21128
rect 27019 21097 27031 21100
rect 26973 21091 27031 21097
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 25590 21020 25596 21072
rect 25648 21060 25654 21072
rect 25648 21032 27476 21060
rect 25648 21020 25654 21032
rect 25590 20924 25596 20936
rect 24912 20896 25452 20924
rect 25503 20896 25596 20924
rect 24912 20884 24918 20896
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20893 25743 20927
rect 26326 20924 26332 20936
rect 26287 20896 26332 20924
rect 25685 20887 25743 20893
rect 21640 20878 21692 20884
rect 13078 20856 13084 20868
rect 9263 20828 12434 20856
rect 13039 20828 13084 20856
rect 9263 20825 9275 20828
rect 9217 20819 9275 20825
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 13265 20859 13323 20865
rect 13265 20825 13277 20859
rect 13311 20856 13323 20859
rect 13814 20856 13820 20868
rect 13311 20828 13820 20856
rect 13311 20825 13323 20828
rect 13265 20819 13323 20825
rect 13814 20816 13820 20828
rect 13872 20816 13878 20868
rect 15657 20859 15715 20865
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 18046 20856 18052 20868
rect 15703 20828 18052 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 18046 20816 18052 20828
rect 18104 20816 18110 20868
rect 19242 20816 19248 20868
rect 19300 20856 19306 20868
rect 19521 20859 19579 20865
rect 19521 20856 19533 20859
rect 19300 20828 19533 20856
rect 19300 20816 19306 20828
rect 19521 20825 19533 20828
rect 19567 20825 19579 20859
rect 21358 20856 21364 20868
rect 19521 20819 19579 20825
rect 19812 20828 21364 20856
rect 19812 20800 19840 20828
rect 21358 20816 21364 20828
rect 21416 20816 21422 20868
rect 22557 20859 22615 20865
rect 22557 20825 22569 20859
rect 22603 20825 22615 20859
rect 22557 20819 22615 20825
rect 2038 20748 2044 20800
rect 2096 20788 2102 20800
rect 2869 20791 2927 20797
rect 2869 20788 2881 20791
rect 2096 20760 2881 20788
rect 2096 20748 2102 20760
rect 2869 20757 2881 20760
rect 2915 20757 2927 20791
rect 2869 20751 2927 20757
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 4617 20791 4675 20797
rect 4617 20788 4629 20791
rect 3108 20760 4629 20788
rect 3108 20748 3114 20760
rect 4617 20757 4629 20760
rect 4663 20788 4675 20791
rect 4798 20788 4804 20800
rect 4663 20760 4804 20788
rect 4663 20757 4675 20760
rect 4617 20751 4675 20757
rect 4798 20748 4804 20760
rect 4856 20748 4862 20800
rect 5258 20748 5264 20800
rect 5316 20788 5322 20800
rect 5442 20788 5448 20800
rect 5316 20760 5448 20788
rect 5316 20748 5322 20760
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 8205 20791 8263 20797
rect 8205 20757 8217 20791
rect 8251 20788 8263 20791
rect 8386 20788 8392 20800
rect 8251 20760 8392 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 9309 20791 9367 20797
rect 9309 20788 9321 20791
rect 8996 20760 9321 20788
rect 8996 20748 9002 20760
rect 9309 20757 9321 20760
rect 9355 20757 9367 20791
rect 9309 20751 9367 20757
rect 10502 20748 10508 20800
rect 10560 20788 10566 20800
rect 10962 20788 10968 20800
rect 10560 20760 10968 20788
rect 10560 20748 10566 20760
rect 10962 20748 10968 20760
rect 11020 20788 11026 20800
rect 11701 20791 11759 20797
rect 11701 20788 11713 20791
rect 11020 20760 11713 20788
rect 11020 20748 11026 20760
rect 11701 20757 11713 20760
rect 11747 20757 11759 20791
rect 11701 20751 11759 20757
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13504 20760 14289 20788
rect 13504 20748 13510 20760
rect 14277 20757 14289 20760
rect 14323 20757 14335 20791
rect 14277 20751 14335 20757
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 18230 20788 18236 20800
rect 17736 20760 18236 20788
rect 17736 20748 17742 20760
rect 18230 20748 18236 20760
rect 18288 20788 18294 20800
rect 18509 20791 18567 20797
rect 18509 20788 18521 20791
rect 18288 20760 18521 20788
rect 18288 20748 18294 20760
rect 18509 20757 18521 20760
rect 18555 20757 18567 20791
rect 19794 20788 19800 20800
rect 19755 20760 19800 20788
rect 18509 20751 18567 20757
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 20530 20788 20536 20800
rect 20404 20760 20536 20788
rect 20404 20748 20410 20760
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 22572 20788 22600 20819
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 25409 20859 25467 20865
rect 25409 20856 25421 20859
rect 23440 20828 25421 20856
rect 23440 20816 23446 20828
rect 25409 20825 25421 20828
rect 25455 20825 25467 20859
rect 25700 20856 25728 20887
rect 26326 20884 26332 20896
rect 26384 20884 26390 20936
rect 26528 20933 26556 21032
rect 27448 20936 27476 21032
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20893 26571 20927
rect 26513 20887 26571 20893
rect 26602 20884 26608 20936
rect 26660 20924 26666 20936
rect 27246 20926 27252 20936
rect 27172 20924 27252 20926
rect 26660 20896 27252 20924
rect 26660 20884 26666 20896
rect 27246 20884 27252 20896
rect 27304 20884 27310 20936
rect 27430 20924 27436 20936
rect 27391 20896 27436 20924
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27522 20884 27528 20936
rect 27580 20924 27586 20936
rect 27893 20927 27951 20933
rect 27893 20924 27905 20927
rect 27580 20896 27905 20924
rect 27580 20884 27586 20896
rect 27893 20893 27905 20896
rect 27939 20893 27951 20927
rect 28074 20924 28080 20936
rect 28035 20896 28080 20924
rect 27893 20887 27951 20893
rect 28074 20884 28080 20896
rect 28132 20884 28138 20936
rect 25409 20819 25467 20825
rect 25516 20828 25728 20856
rect 26421 20859 26479 20865
rect 23842 20788 23848 20800
rect 22572 20760 23848 20788
rect 23842 20748 23848 20760
rect 23900 20788 23906 20800
rect 25516 20788 25544 20828
rect 26421 20825 26433 20859
rect 26467 20856 26479 20859
rect 26467 20828 27292 20856
rect 26467 20825 26479 20828
rect 26421 20819 26479 20825
rect 27264 20800 27292 20828
rect 27154 20788 27160 20800
rect 23900 20760 25544 20788
rect 27115 20760 27160 20788
rect 23900 20748 23906 20760
rect 27154 20748 27160 20760
rect 27212 20748 27218 20800
rect 27246 20748 27252 20800
rect 27304 20748 27310 20800
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 27985 20791 28043 20797
rect 27985 20788 27997 20791
rect 27672 20760 27997 20788
rect 27672 20748 27678 20760
rect 27985 20757 27997 20760
rect 28031 20757 28043 20791
rect 27985 20751 28043 20757
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 3237 20587 3295 20593
rect 3237 20553 3249 20587
rect 3283 20584 3295 20587
rect 7650 20584 7656 20596
rect 3283 20556 7656 20584
rect 3283 20553 3295 20556
rect 3237 20547 3295 20553
rect 7650 20544 7656 20556
rect 7708 20544 7714 20596
rect 7834 20544 7840 20596
rect 7892 20584 7898 20596
rect 8478 20584 8484 20596
rect 7892 20556 8340 20584
rect 7892 20544 7898 20556
rect 2501 20519 2559 20525
rect 2501 20485 2513 20519
rect 2547 20516 2559 20519
rect 2547 20488 2636 20516
rect 2547 20485 2559 20488
rect 2501 20479 2559 20485
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 1811 20420 2237 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 2608 20312 2636 20488
rect 2682 20476 2688 20528
rect 2740 20516 2746 20528
rect 2740 20488 2833 20516
rect 2740 20476 2746 20488
rect 3326 20476 3332 20528
rect 3384 20516 3390 20528
rect 3421 20519 3479 20525
rect 3421 20516 3433 20519
rect 3384 20488 3433 20516
rect 3384 20476 3390 20488
rect 3421 20485 3433 20488
rect 3467 20485 3479 20519
rect 3421 20479 3479 20485
rect 3605 20519 3663 20525
rect 3605 20485 3617 20519
rect 3651 20516 3663 20519
rect 4154 20516 4160 20528
rect 3651 20488 4160 20516
rect 3651 20485 3663 20488
rect 3605 20479 3663 20485
rect 4154 20476 4160 20488
rect 4212 20476 4218 20528
rect 5534 20516 5540 20528
rect 4264 20488 5540 20516
rect 2700 20448 2728 20476
rect 4264 20448 4292 20488
rect 5534 20476 5540 20488
rect 5592 20476 5598 20528
rect 5718 20476 5724 20528
rect 5776 20516 5782 20528
rect 8312 20525 8340 20556
rect 8404 20556 8484 20584
rect 8404 20525 8432 20556
rect 8478 20544 8484 20556
rect 8536 20544 8542 20596
rect 8665 20587 8723 20593
rect 8665 20553 8677 20587
rect 8711 20584 8723 20587
rect 12253 20587 12311 20593
rect 8711 20556 10640 20584
rect 8711 20553 8723 20556
rect 8665 20547 8723 20553
rect 8297 20519 8355 20525
rect 5776 20488 8228 20516
rect 5776 20476 5782 20488
rect 2700 20420 4292 20448
rect 4332 20451 4390 20457
rect 4332 20417 4344 20451
rect 4378 20448 4390 20451
rect 4890 20448 4896 20460
rect 4378 20420 4896 20448
rect 4378 20417 4390 20420
rect 4332 20411 4390 20417
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 6512 20420 7297 20448
rect 6512 20408 6518 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 4062 20380 4068 20392
rect 3108 20352 4068 20380
rect 3108 20340 3114 20352
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 7300 20312 7328 20411
rect 7484 20380 7512 20411
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 7926 20448 7932 20460
rect 7616 20420 7932 20448
rect 7616 20408 7622 20420
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 8200 20457 8228 20488
rect 8297 20485 8309 20519
rect 8343 20485 8355 20519
rect 8297 20479 8355 20485
rect 8389 20519 8447 20525
rect 8389 20485 8401 20519
rect 8435 20485 8447 20519
rect 9582 20516 9588 20528
rect 8389 20479 8447 20485
rect 8542 20488 9588 20516
rect 8542 20457 8570 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 10226 20476 10232 20528
rect 10284 20525 10290 20528
rect 10284 20516 10296 20525
rect 10284 20488 10329 20516
rect 10284 20479 10296 20488
rect 10284 20476 10290 20479
rect 8169 20451 8228 20457
rect 8076 20420 8121 20448
rect 8076 20408 8082 20420
rect 8169 20417 8181 20451
rect 8215 20420 8228 20451
rect 8527 20451 8585 20457
rect 8215 20417 8227 20420
rect 8169 20411 8227 20417
rect 8527 20417 8539 20451
rect 8573 20417 8585 20451
rect 10502 20448 10508 20460
rect 10463 20420 10508 20448
rect 8527 20411 8585 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 7650 20380 7656 20392
rect 7484 20352 7656 20380
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 8938 20380 8944 20392
rect 7760 20352 8944 20380
rect 7760 20312 7788 20352
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 10612 20380 10640 20556
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 12618 20584 12624 20596
rect 12299 20556 12624 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 13170 20584 13176 20596
rect 12728 20556 13176 20584
rect 12728 20516 12756 20556
rect 13170 20544 13176 20556
rect 13228 20544 13234 20596
rect 22465 20587 22523 20593
rect 14660 20556 22094 20584
rect 13354 20516 13360 20528
rect 11164 20488 12756 20516
rect 13188 20488 13360 20516
rect 10962 20448 10968 20460
rect 10923 20420 10968 20448
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11164 20457 11192 20488
rect 13188 20470 13216 20488
rect 13354 20476 13360 20488
rect 13412 20476 13418 20528
rect 14660 20525 14688 20556
rect 14645 20519 14703 20525
rect 14645 20485 14657 20519
rect 14691 20485 14703 20519
rect 14645 20479 14703 20485
rect 15657 20519 15715 20525
rect 15657 20485 15669 20519
rect 15703 20516 15715 20519
rect 16574 20516 16580 20528
rect 15703 20488 16580 20516
rect 15703 20485 15715 20488
rect 15657 20479 15715 20485
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 16666 20476 16672 20528
rect 16724 20516 16730 20528
rect 16853 20519 16911 20525
rect 16853 20516 16865 20519
rect 16724 20488 16865 20516
rect 16724 20476 16730 20488
rect 16853 20485 16865 20488
rect 16899 20485 16911 20519
rect 19150 20516 19156 20528
rect 16853 20479 16911 20485
rect 19076 20488 19156 20516
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20417 11207 20451
rect 11882 20448 11888 20460
rect 11843 20420 11888 20448
rect 11149 20411 11207 20417
rect 11882 20408 11888 20420
rect 11940 20408 11946 20460
rect 12066 20448 12072 20460
rect 12027 20420 12072 20448
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 13003 20457 13216 20470
rect 12804 20451 12862 20457
rect 12804 20448 12816 20451
rect 12768 20420 12816 20448
rect 12768 20408 12774 20420
rect 12804 20417 12816 20420
rect 12850 20417 12862 20451
rect 12804 20411 12862 20417
rect 12988 20451 13216 20457
rect 12988 20417 13000 20451
rect 13034 20442 13216 20451
rect 14274 20448 14280 20460
rect 13034 20417 13046 20442
rect 14235 20420 14280 20448
rect 12988 20411 13046 20417
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15436 20420 15577 20448
rect 15436 20408 15442 20420
rect 15565 20417 15577 20420
rect 15611 20448 15623 20451
rect 15746 20448 15752 20460
rect 15611 20420 15752 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16114 20448 16120 20460
rect 15887 20420 16120 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 19076 20457 19104 20488
rect 19150 20476 19156 20488
rect 19208 20516 19214 20528
rect 22066 20516 22094 20556
rect 22465 20553 22477 20587
rect 22511 20584 22523 20587
rect 23474 20584 23480 20596
rect 22511 20556 23480 20584
rect 22511 20553 22523 20556
rect 22465 20547 22523 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23658 20544 23664 20596
rect 23716 20584 23722 20596
rect 24762 20584 24768 20596
rect 23716 20556 24768 20584
rect 23716 20544 23722 20556
rect 24762 20544 24768 20556
rect 24820 20584 24826 20596
rect 27525 20587 27583 20593
rect 24820 20556 25360 20584
rect 24820 20544 24826 20556
rect 25225 20519 25283 20525
rect 25225 20516 25237 20519
rect 19208 20488 21220 20516
rect 22066 20488 25237 20516
rect 19208 20476 19214 20488
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19334 20448 19340 20460
rect 19295 20420 19340 20448
rect 19061 20411 19119 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19610 20448 19616 20460
rect 19484 20420 19616 20448
rect 19484 20408 19490 20420
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19886 20448 19892 20460
rect 19847 20420 19892 20448
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20438 20448 20444 20460
rect 20119 20420 20444 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20714 20448 20720 20460
rect 20588 20420 20633 20448
rect 20675 20420 20720 20448
rect 20588 20408 20594 20420
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 21192 20457 21220 20488
rect 25225 20485 25237 20488
rect 25271 20485 25283 20519
rect 25225 20479 25283 20485
rect 21177 20451 21235 20457
rect 21177 20417 21189 20451
rect 21223 20417 21235 20451
rect 21177 20411 21235 20417
rect 21542 20408 21548 20460
rect 21600 20448 21606 20460
rect 22002 20448 22008 20460
rect 21600 20420 22008 20448
rect 21600 20408 21606 20420
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20448 22983 20451
rect 23566 20448 23572 20460
rect 22971 20420 23572 20448
rect 22971 20417 22983 20420
rect 22925 20411 22983 20417
rect 11793 20383 11851 20389
rect 11793 20380 11805 20383
rect 10612 20352 11805 20380
rect 11793 20349 11805 20352
rect 11839 20349 11851 20383
rect 11974 20380 11980 20392
rect 11935 20352 11980 20380
rect 11793 20343 11851 20349
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 12896 20383 12954 20389
rect 12896 20349 12908 20383
rect 12942 20349 12954 20383
rect 12896 20343 12954 20349
rect 13081 20383 13139 20389
rect 13081 20349 13093 20383
rect 13127 20380 13139 20383
rect 13170 20380 13176 20392
rect 13127 20352 13176 20380
rect 13127 20349 13139 20352
rect 13081 20343 13139 20349
rect 2608 20284 4108 20312
rect 7300 20284 7788 20312
rect 11149 20315 11207 20321
rect 4080 20256 4108 20284
rect 11149 20281 11161 20315
rect 11195 20312 11207 20315
rect 12434 20312 12440 20324
rect 11195 20284 12440 20312
rect 11195 20281 11207 20284
rect 11149 20275 11207 20281
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 12802 20272 12808 20324
rect 12860 20312 12866 20324
rect 12912 20312 12940 20343
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 14182 20380 14188 20392
rect 14143 20352 14188 20380
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 14366 20340 14372 20392
rect 14424 20380 14430 20392
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 14424 20352 14565 20380
rect 14424 20340 14430 20352
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 14918 20340 14924 20392
rect 14976 20380 14982 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 14976 20352 20637 20380
rect 14976 20340 14982 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 22940 20380 22968 20411
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 25332 20457 25360 20556
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 27706 20584 27712 20596
rect 27571 20556 27712 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 27706 20544 27712 20556
rect 27764 20544 27770 20596
rect 27338 20476 27344 20528
rect 27396 20516 27402 20528
rect 27617 20519 27675 20525
rect 27617 20516 27629 20519
rect 27396 20488 27629 20516
rect 27396 20476 27402 20488
rect 27617 20485 27629 20488
rect 27663 20485 27675 20519
rect 27617 20479 27675 20485
rect 25133 20451 25191 20457
rect 25133 20448 25145 20451
rect 24636 20420 25145 20448
rect 24636 20408 24642 20420
rect 25133 20417 25145 20420
rect 25179 20417 25191 20451
rect 25133 20411 25191 20417
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20417 26295 20451
rect 26237 20411 26295 20417
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20448 26479 20451
rect 26510 20448 26516 20460
rect 26467 20420 26516 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 23842 20380 23848 20392
rect 20956 20352 22968 20380
rect 23803 20352 23848 20380
rect 20956 20340 20962 20352
rect 23842 20340 23848 20352
rect 23900 20340 23906 20392
rect 24673 20383 24731 20389
rect 24673 20349 24685 20383
rect 24719 20380 24731 20383
rect 26252 20380 26280 20411
rect 26510 20408 26516 20420
rect 26568 20408 26574 20460
rect 26326 20380 26332 20392
rect 24719 20352 26332 20380
rect 24719 20349 24731 20352
rect 24673 20343 24731 20349
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20349 27491 20383
rect 27433 20343 27491 20349
rect 12860 20284 12940 20312
rect 12860 20272 12866 20284
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 14384 20312 14412 20340
rect 13872 20284 14412 20312
rect 13872 20272 13878 20284
rect 15470 20272 15476 20324
rect 15528 20312 15534 20324
rect 17218 20312 17224 20324
rect 15528 20284 17224 20312
rect 15528 20272 15534 20284
rect 17218 20272 17224 20284
rect 17276 20272 17282 20324
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 21450 20312 21456 20324
rect 20588 20284 21456 20312
rect 20588 20272 20594 20284
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 21634 20272 21640 20324
rect 21692 20312 21698 20324
rect 22281 20315 22339 20321
rect 22281 20312 22293 20315
rect 21692 20284 22293 20312
rect 21692 20272 21698 20284
rect 22281 20281 22293 20284
rect 22327 20281 22339 20315
rect 27448 20312 27476 20343
rect 27614 20312 27620 20324
rect 27448 20284 27620 20312
rect 22281 20275 22339 20281
rect 27614 20272 27620 20284
rect 27672 20272 27678 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2498 20244 2504 20256
rect 2459 20216 2504 20244
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 3421 20247 3479 20253
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 3786 20244 3792 20256
rect 3467 20216 3792 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 4062 20204 4068 20256
rect 4120 20204 4126 20256
rect 4246 20204 4252 20256
rect 4304 20244 4310 20256
rect 5445 20247 5503 20253
rect 5445 20244 5457 20247
rect 4304 20216 5457 20244
rect 4304 20204 4310 20216
rect 5445 20213 5457 20216
rect 5491 20244 5503 20247
rect 5810 20244 5816 20256
rect 5491 20216 5816 20244
rect 5491 20213 5503 20216
rect 5445 20207 5503 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6362 20244 6368 20256
rect 6043 20216 6368 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 6546 20244 6552 20256
rect 6507 20216 6552 20244
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 7098 20244 7104 20256
rect 7059 20216 7104 20244
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 7834 20244 7840 20256
rect 7524 20216 7840 20244
rect 7524 20204 7530 20216
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8444 20216 9137 20244
rect 8444 20204 8450 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 13170 20244 13176 20256
rect 9364 20216 13176 20244
rect 9364 20204 9370 20216
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 13265 20247 13323 20253
rect 13265 20213 13277 20247
rect 13311 20244 13323 20247
rect 13354 20244 13360 20256
rect 13311 20216 13360 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 13998 20244 14004 20256
rect 13959 20216 14004 20244
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 16022 20244 16028 20256
rect 15983 20216 16028 20244
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18141 20247 18199 20253
rect 18141 20244 18153 20247
rect 18104 20216 18153 20244
rect 18104 20204 18110 20216
rect 18141 20213 18153 20216
rect 18187 20213 18199 20247
rect 18141 20207 18199 20213
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 19576 20216 19901 20244
rect 19576 20204 19582 20216
rect 19889 20213 19901 20216
rect 19935 20213 19947 20247
rect 19889 20207 19947 20213
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 22554 20244 22560 20256
rect 21315 20216 22560 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 22554 20204 22560 20216
rect 22612 20204 22618 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 26329 20247 26387 20253
rect 26329 20213 26341 20247
rect 26375 20244 26387 20247
rect 27062 20244 27068 20256
rect 26375 20216 27068 20244
rect 26375 20213 26387 20216
rect 26329 20207 26387 20213
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 27982 20244 27988 20256
rect 27943 20216 27988 20244
rect 27982 20204 27988 20216
rect 28040 20204 28046 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 4525 20043 4583 20049
rect 4525 20040 4537 20043
rect 3844 20012 4537 20040
rect 3844 20000 3850 20012
rect 4525 20009 4537 20012
rect 4571 20040 4583 20043
rect 4706 20040 4712 20052
rect 4571 20012 4712 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 5721 20043 5779 20049
rect 5721 20009 5733 20043
rect 5767 20040 5779 20043
rect 7742 20040 7748 20052
rect 5767 20012 7748 20040
rect 5767 20009 5779 20012
rect 5721 20003 5779 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 7834 20000 7840 20052
rect 7892 20000 7898 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8662 20040 8668 20052
rect 7984 20012 8668 20040
rect 7984 20000 7990 20012
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 11112 20012 11713 20040
rect 11112 20000 11118 20012
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 12069 20043 12127 20049
rect 12069 20009 12081 20043
rect 12115 20040 12127 20043
rect 12710 20040 12716 20052
rect 12115 20012 12716 20040
rect 12115 20009 12127 20012
rect 12069 20003 12127 20009
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 13354 20040 13360 20052
rect 13315 20012 13360 20040
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 15470 20040 15476 20052
rect 15431 20012 15476 20040
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 17862 20040 17868 20052
rect 16264 20012 16988 20040
rect 17823 20012 17868 20040
rect 16264 20000 16270 20012
rect 3421 19975 3479 19981
rect 3421 19941 3433 19975
rect 3467 19941 3479 19975
rect 3421 19935 3479 19941
rect 2038 19904 2044 19916
rect 1999 19876 2044 19904
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 3436 19904 3464 19935
rect 7282 19932 7288 19984
rect 7340 19972 7346 19984
rect 7340 19944 7788 19972
rect 7340 19932 7346 19944
rect 7760 19916 7788 19944
rect 3602 19904 3608 19916
rect 3436 19876 3608 19904
rect 3602 19864 3608 19876
rect 3660 19904 3666 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 3660 19876 7573 19904
rect 3660 19864 3666 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 7561 19867 7619 19873
rect 7742 19864 7748 19916
rect 7800 19864 7806 19916
rect 2308 19839 2366 19845
rect 2308 19805 2320 19839
rect 2354 19836 2366 19839
rect 3142 19836 3148 19848
rect 2354 19808 3148 19836
rect 2354 19805 2366 19808
rect 2308 19799 2366 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 6546 19836 6552 19848
rect 4080 19808 6552 19836
rect 4080 19768 4108 19808
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19836 7067 19839
rect 7190 19836 7196 19848
rect 7055 19808 7196 19836
rect 7055 19805 7067 19808
rect 7009 19799 7067 19805
rect 7190 19796 7196 19808
rect 7248 19796 7254 19848
rect 7852 19845 7880 20000
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 8168 19944 9812 19972
rect 8168 19932 8174 19944
rect 8128 19904 8156 19932
rect 9490 19904 9496 19916
rect 8036 19876 8156 19904
rect 9451 19876 9496 19904
rect 8036 19845 8064 19876
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 9674 19904 9680 19916
rect 9635 19876 9680 19904
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 7837 19839 7895 19845
rect 7837 19805 7849 19839
rect 7883 19805 7895 19839
rect 7837 19799 7895 19805
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8168 19808 9413 19836
rect 8168 19796 8174 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19836 9643 19839
rect 9784 19836 9812 19944
rect 10962 19932 10968 19984
rect 11020 19972 11026 19984
rect 14182 19972 14188 19984
rect 11020 19944 14188 19972
rect 11020 19932 11026 19944
rect 11974 19904 11980 19916
rect 10704 19876 11980 19904
rect 10704 19836 10732 19876
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12526 19904 12532 19916
rect 12487 19876 12532 19904
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 10870 19836 10876 19848
rect 9631 19808 10732 19836
rect 10831 19808 10876 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 2746 19740 4108 19768
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 2746 19700 2774 19740
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 4341 19771 4399 19777
rect 4341 19768 4353 19771
rect 4212 19740 4353 19768
rect 4212 19728 4218 19740
rect 4341 19737 4353 19740
rect 4387 19737 4399 19771
rect 4890 19768 4896 19780
rect 4341 19731 4399 19737
rect 4540 19740 4896 19768
rect 4540 19709 4568 19740
rect 4890 19728 4896 19740
rect 4948 19768 4954 19780
rect 5626 19768 5632 19780
rect 4948 19740 5632 19768
rect 4948 19728 4954 19740
rect 5626 19728 5632 19740
rect 5684 19768 5690 19780
rect 6822 19768 6828 19780
rect 5684 19740 6828 19768
rect 5684 19728 5690 19740
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7742 19777 7748 19780
rect 7719 19771 7748 19777
rect 7719 19737 7731 19771
rect 7719 19731 7748 19737
rect 7742 19728 7748 19731
rect 7800 19728 7806 19780
rect 7928 19771 7986 19777
rect 7928 19737 7940 19771
rect 7974 19768 7986 19771
rect 8386 19768 8392 19780
rect 7974 19740 8392 19768
rect 7974 19737 7986 19740
rect 7928 19731 7986 19737
rect 8386 19728 8392 19740
rect 8444 19728 8450 19780
rect 8478 19728 8484 19780
rect 8536 19768 8542 19780
rect 11238 19768 11244 19780
rect 8536 19740 11244 19768
rect 8536 19728 8542 19740
rect 11238 19728 11244 19740
rect 11296 19728 11302 19780
rect 11716 19768 11744 19799
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12618 19836 12624 19848
rect 11848 19808 11893 19836
rect 12579 19808 12624 19836
rect 11848 19796 11854 19808
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13280 19836 13308 19944
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 13998 19904 14004 19916
rect 13372 19876 14004 19904
rect 13372 19845 13400 19876
rect 13998 19864 14004 19876
rect 14056 19864 14062 19916
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 14918 19904 14924 19916
rect 14700 19876 14780 19904
rect 14879 19876 14924 19904
rect 14700 19864 14706 19876
rect 12943 19808 13308 19836
rect 13357 19839 13415 19845
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13630 19836 13636 19848
rect 13587 19808 13636 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 13780 19808 14473 19836
rect 13780 19796 13786 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 14752 19836 14780 19876
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 14829 19839 14887 19845
rect 14829 19836 14841 19839
rect 14608 19808 14653 19836
rect 14752 19808 14841 19836
rect 14608 19796 14614 19808
rect 14829 19805 14841 19808
rect 14875 19805 14887 19839
rect 15930 19836 15936 19848
rect 15891 19808 15936 19836
rect 14829 19799 14887 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16022 19796 16028 19848
rect 16080 19836 16086 19848
rect 16189 19839 16247 19845
rect 16189 19836 16201 19839
rect 16080 19808 16201 19836
rect 16080 19796 16086 19808
rect 16189 19805 16201 19808
rect 16235 19805 16247 19839
rect 16960 19836 16988 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 19610 20000 19616 20052
rect 19668 20040 19674 20052
rect 20070 20040 20076 20052
rect 19668 20012 20076 20040
rect 19668 20000 19674 20012
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 22189 20043 22247 20049
rect 22189 20009 22201 20043
rect 22235 20040 22247 20043
rect 23290 20040 23296 20052
rect 22235 20012 23296 20040
rect 22235 20009 22247 20012
rect 22189 20003 22247 20009
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 23842 20040 23848 20052
rect 23400 20012 23848 20040
rect 17313 19975 17371 19981
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 20806 19972 20812 19984
rect 17359 19944 20812 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 20806 19932 20812 19944
rect 20864 19972 20870 19984
rect 21174 19972 21180 19984
rect 20864 19944 21180 19972
rect 20864 19932 20870 19944
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 22002 19972 22008 19984
rect 21963 19944 22008 19972
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 20530 19904 20536 19916
rect 18156 19876 20536 19904
rect 18049 19839 18107 19845
rect 18049 19836 18061 19839
rect 16960 19808 18061 19836
rect 16189 19799 16247 19805
rect 18049 19805 18061 19808
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 14277 19771 14335 19777
rect 14277 19768 14289 19771
rect 11716 19740 14289 19768
rect 14277 19737 14289 19740
rect 14323 19737 14335 19771
rect 14277 19731 14335 19737
rect 2280 19672 2774 19700
rect 4525 19703 4583 19709
rect 2280 19660 2286 19672
rect 4525 19669 4537 19703
rect 4571 19669 4583 19703
rect 4525 19663 4583 19669
rect 4709 19703 4767 19709
rect 4709 19669 4721 19703
rect 4755 19700 4767 19703
rect 7466 19700 7472 19712
rect 4755 19672 7472 19700
rect 4755 19669 4767 19672
rect 4709 19663 4767 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7616 19672 8217 19700
rect 7616 19660 7622 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 8205 19663 8263 19669
rect 9861 19703 9919 19709
rect 9861 19669 9873 19703
rect 9907 19700 9919 19703
rect 10134 19700 10140 19712
rect 9907 19672 10140 19700
rect 9907 19669 9919 19672
rect 9861 19663 9919 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 13725 19703 13783 19709
rect 13725 19700 13737 19703
rect 13688 19672 13737 19700
rect 13688 19660 13694 19672
rect 13725 19669 13737 19672
rect 13771 19669 13783 19703
rect 13725 19663 13783 19669
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 14737 19703 14795 19709
rect 14737 19700 14749 19703
rect 14056 19672 14749 19700
rect 14056 19660 14062 19672
rect 14737 19669 14749 19672
rect 14783 19700 14795 19703
rect 14826 19700 14832 19712
rect 14783 19672 14832 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 18156 19700 18184 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21692 19876 21741 19904
rect 21692 19864 21698 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 23400 19904 23428 20012
rect 23842 20000 23848 20012
rect 23900 20000 23906 20052
rect 24026 20040 24032 20052
rect 23987 20012 24032 20040
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 25317 20043 25375 20049
rect 25317 20009 25329 20043
rect 25363 20040 25375 20043
rect 25590 20040 25596 20052
rect 25363 20012 25596 20040
rect 25363 20009 25375 20012
rect 25317 20003 25375 20009
rect 25590 20000 25596 20012
rect 25648 20000 25654 20052
rect 27893 20043 27951 20049
rect 27893 20009 27905 20043
rect 27939 20040 27951 20043
rect 28074 20040 28080 20052
rect 27939 20012 28080 20040
rect 27939 20009 27951 20012
rect 27893 20003 27951 20009
rect 28074 20000 28080 20012
rect 28132 20000 28138 20052
rect 25961 19907 26019 19913
rect 25961 19904 25973 19907
rect 21729 19867 21787 19873
rect 23032 19876 23428 19904
rect 23584 19876 25973 19904
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19830 18383 19839
rect 18414 19830 18420 19848
rect 18371 19805 18420 19830
rect 18325 19802 18420 19805
rect 18325 19799 18383 19802
rect 18414 19796 18420 19802
rect 18472 19796 18478 19848
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 19426 19836 19432 19848
rect 18564 19808 19432 19836
rect 18564 19796 18570 19808
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19610 19836 19616 19848
rect 19571 19808 19616 19836
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 19886 19836 19892 19848
rect 19847 19808 19892 19836
rect 19886 19796 19892 19808
rect 19944 19836 19950 19848
rect 20622 19836 20628 19848
rect 19944 19808 20628 19836
rect 19944 19796 19950 19808
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22738 19836 22744 19848
rect 22244 19808 22744 19836
rect 22244 19796 22250 19808
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23032 19845 23060 19876
rect 23017 19839 23075 19845
rect 23017 19805 23029 19839
rect 23063 19805 23075 19839
rect 23474 19836 23480 19848
rect 23435 19808 23480 19836
rect 23017 19799 23075 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 23584 19845 23612 19876
rect 25961 19873 25973 19876
rect 26007 19873 26019 19907
rect 27338 19904 27344 19916
rect 25961 19867 26019 19873
rect 27080 19876 27344 19904
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 19058 19728 19064 19780
rect 19116 19768 19122 19780
rect 20441 19771 20499 19777
rect 20441 19768 20453 19771
rect 19116 19740 20453 19768
rect 19116 19728 19122 19740
rect 20441 19737 20453 19740
rect 20487 19768 20499 19771
rect 20898 19768 20904 19780
rect 20487 19740 20904 19768
rect 20487 19737 20499 19740
rect 20441 19731 20499 19737
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 22925 19771 22983 19777
rect 22925 19737 22937 19771
rect 22971 19768 22983 19771
rect 23658 19768 23664 19780
rect 22971 19740 23664 19768
rect 22971 19737 22983 19740
rect 22925 19731 22983 19737
rect 23658 19728 23664 19740
rect 23716 19768 23722 19780
rect 23768 19768 23796 19799
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 24394 19836 24400 19848
rect 23900 19808 24400 19836
rect 23900 19796 23906 19808
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 25225 19839 25283 19845
rect 25225 19836 25237 19839
rect 24811 19808 25237 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 25225 19805 25237 19808
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 23716 19740 23796 19768
rect 23716 19728 23722 19740
rect 24302 19728 24308 19780
rect 24360 19768 24366 19780
rect 24780 19768 24808 19799
rect 24360 19740 24808 19768
rect 24360 19728 24366 19740
rect 24854 19728 24860 19780
rect 24912 19768 24918 19780
rect 25424 19768 25452 19799
rect 25590 19796 25596 19848
rect 25648 19836 25654 19848
rect 27080 19845 27108 19876
rect 27338 19864 27344 19876
rect 27396 19904 27402 19916
rect 27396 19876 28212 19904
rect 27396 19864 27402 19876
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25648 19808 25881 19836
rect 25648 19796 25654 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 27065 19839 27123 19845
rect 27065 19805 27077 19839
rect 27111 19805 27123 19839
rect 27065 19799 27123 19805
rect 27154 19796 27160 19848
rect 27212 19836 27218 19848
rect 28184 19845 28212 19876
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27212 19808 27445 19836
rect 27212 19796 27218 19808
rect 27433 19805 27445 19808
rect 27479 19805 27491 19839
rect 27433 19799 27491 19805
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 24912 19740 25452 19768
rect 24912 19728 24918 19740
rect 26142 19728 26148 19780
rect 26200 19768 26206 19780
rect 26881 19771 26939 19777
rect 26881 19768 26893 19771
rect 26200 19740 26893 19768
rect 26200 19728 26206 19740
rect 26881 19737 26893 19740
rect 26927 19737 26939 19771
rect 27890 19768 27896 19780
rect 26881 19731 26939 19737
rect 27172 19740 27476 19768
rect 27851 19740 27896 19768
rect 27172 19712 27200 19740
rect 18233 19703 18291 19709
rect 18233 19700 18245 19703
rect 18156 19672 18245 19700
rect 18233 19669 18245 19672
rect 18279 19669 18291 19703
rect 18233 19663 18291 19669
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 19426 19700 19432 19712
rect 18840 19672 18885 19700
rect 19387 19672 19432 19700
rect 18840 19660 18846 19672
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 19843 19672 20545 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20533 19669 20545 19672
rect 20579 19700 20591 19703
rect 21358 19700 21364 19712
rect 20579 19672 21364 19700
rect 20579 19669 20591 19672
rect 20533 19663 20591 19669
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 22839 19703 22897 19709
rect 22839 19669 22851 19703
rect 22885 19700 22897 19703
rect 23382 19700 23388 19712
rect 22885 19672 23388 19700
rect 22885 19669 22897 19672
rect 22839 19663 22897 19669
rect 23382 19660 23388 19672
rect 23440 19660 23446 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 24673 19703 24731 19709
rect 24673 19700 24685 19703
rect 23624 19672 24685 19700
rect 23624 19660 23630 19672
rect 24673 19669 24685 19672
rect 24719 19669 24731 19703
rect 27154 19700 27160 19712
rect 27115 19672 27160 19700
rect 24673 19663 24731 19669
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 27246 19660 27252 19712
rect 27304 19700 27310 19712
rect 27448 19700 27476 19740
rect 27890 19728 27896 19740
rect 27948 19728 27954 19780
rect 28077 19703 28135 19709
rect 28077 19700 28089 19703
rect 27304 19672 27349 19700
rect 27448 19672 28089 19700
rect 27304 19660 27310 19672
rect 28077 19669 28089 19672
rect 28123 19669 28135 19703
rect 28077 19663 28135 19669
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 3421 19499 3479 19505
rect 3421 19496 3433 19499
rect 3292 19468 3433 19496
rect 3292 19456 3298 19468
rect 3421 19465 3433 19468
rect 3467 19465 3479 19499
rect 3421 19459 3479 19465
rect 4249 19499 4307 19505
rect 4249 19465 4261 19499
rect 4295 19496 4307 19499
rect 5994 19496 6000 19508
rect 4295 19468 6000 19496
rect 4295 19465 4307 19468
rect 4249 19459 4307 19465
rect 5994 19456 6000 19468
rect 6052 19456 6058 19508
rect 8021 19499 8079 19505
rect 8021 19465 8033 19499
rect 8067 19496 8079 19499
rect 8294 19496 8300 19508
rect 8067 19468 8300 19496
rect 8067 19465 8079 19468
rect 8021 19459 8079 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 12710 19496 12716 19508
rect 9640 19456 9674 19496
rect 12671 19468 12716 19496
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 13170 19456 13176 19508
rect 13228 19496 13234 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13228 19468 13461 19496
rect 13228 19456 13234 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 15470 19496 15476 19508
rect 13449 19459 13507 19465
rect 13740 19468 15476 19496
rect 2308 19431 2366 19437
rect 2308 19397 2320 19431
rect 2354 19428 2366 19431
rect 2866 19428 2872 19440
rect 2354 19400 2872 19428
rect 2354 19397 2366 19400
rect 2308 19391 2366 19397
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 5350 19428 5356 19440
rect 5311 19400 5356 19428
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 5442 19388 5448 19440
rect 5500 19428 5506 19440
rect 6908 19431 6966 19437
rect 5500 19400 5545 19428
rect 5500 19388 5506 19400
rect 6908 19397 6920 19431
rect 6954 19428 6966 19431
rect 7006 19428 7012 19440
rect 6954 19400 7012 19428
rect 6954 19397 6966 19400
rect 6908 19391 6966 19397
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 7650 19388 7656 19440
rect 7708 19428 7714 19440
rect 9493 19431 9551 19437
rect 9493 19428 9505 19431
rect 7708 19400 9505 19428
rect 7708 19388 7714 19400
rect 9493 19397 9505 19400
rect 9539 19397 9551 19431
rect 9493 19391 9551 19397
rect 2038 19360 2044 19372
rect 1999 19332 2044 19360
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19360 4215 19363
rect 4430 19360 4436 19372
rect 4203 19332 4292 19360
rect 4391 19332 4436 19360
rect 4203 19329 4215 19332
rect 4157 19323 4215 19329
rect 4264 19292 4292 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5261 19363 5319 19369
rect 5261 19360 5273 19363
rect 4948 19332 5273 19360
rect 4948 19320 4954 19332
rect 5261 19329 5273 19332
rect 5307 19329 5319 19363
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5261 19323 5319 19329
rect 5368 19332 5641 19360
rect 5074 19292 5080 19304
rect 4264 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5166 19184 5172 19236
rect 5224 19224 5230 19236
rect 5368 19224 5396 19332
rect 5629 19329 5641 19332
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 6730 19360 6736 19372
rect 6687 19332 6736 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 8665 19363 8723 19369
rect 8665 19360 8677 19363
rect 7524 19332 8677 19360
rect 7524 19320 7530 19332
rect 8665 19329 8677 19332
rect 8711 19329 8723 19363
rect 8665 19323 8723 19329
rect 8754 19320 8760 19372
rect 8812 19360 8818 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 8812 19332 9137 19360
rect 8812 19320 8818 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 9214 19320 9220 19372
rect 9272 19360 9278 19372
rect 9646 19369 9674 19456
rect 10321 19431 10379 19437
rect 10321 19397 10333 19431
rect 10367 19428 10379 19431
rect 10410 19428 10416 19440
rect 10367 19400 10416 19428
rect 10367 19397 10379 19400
rect 10321 19391 10379 19397
rect 10410 19388 10416 19400
rect 10468 19428 10474 19440
rect 13740 19428 13768 19468
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 18417 19499 18475 19505
rect 18417 19465 18429 19499
rect 18463 19496 18475 19499
rect 19058 19496 19064 19508
rect 18463 19468 19064 19496
rect 18463 19465 18475 19468
rect 18417 19459 18475 19465
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19705 19499 19763 19505
rect 19705 19496 19717 19499
rect 19199 19468 19717 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19705 19465 19717 19468
rect 19751 19465 19763 19499
rect 19705 19459 19763 19465
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 24578 19496 24584 19508
rect 21232 19468 24584 19496
rect 21232 19456 21238 19468
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 26050 19496 26056 19508
rect 24780 19468 26056 19496
rect 10468 19400 13768 19428
rect 10468 19388 10474 19400
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 17304 19431 17362 19437
rect 15436 19400 17264 19428
rect 15436 19388 15442 19400
rect 9401 19363 9459 19369
rect 9272 19332 9317 19360
rect 9272 19320 9278 19332
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9631 19363 9689 19369
rect 9447 19332 9536 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 5224 19196 5396 19224
rect 9508 19224 9536 19332
rect 9631 19329 9643 19363
rect 9677 19329 9689 19363
rect 11698 19360 11704 19372
rect 11659 19332 11704 19360
rect 9631 19323 9689 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19360 12403 19363
rect 13446 19360 13452 19372
rect 12391 19332 13452 19360
rect 12391 19329 12403 19332
rect 12345 19323 12403 19329
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13817 19363 13875 19369
rect 13817 19329 13829 19363
rect 13863 19360 13875 19363
rect 13998 19360 14004 19372
rect 13863 19332 14004 19360
rect 13863 19329 13875 19332
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 13556 19301 13676 19326
rect 13817 19323 13875 19329
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 15988 19332 17049 19360
rect 15988 19320 15994 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17236 19360 17264 19400
rect 17304 19397 17316 19431
rect 17350 19428 17362 19431
rect 19426 19428 19432 19440
rect 17350 19400 19432 19428
rect 17350 19397 17362 19400
rect 17304 19391 17362 19397
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 21266 19388 21272 19440
rect 21324 19428 21330 19440
rect 21324 19400 22416 19428
rect 21324 19388 21330 19400
rect 18414 19360 18420 19372
rect 17236 19332 18420 19360
rect 17037 19323 17095 19329
rect 18414 19320 18420 19332
rect 18472 19360 18478 19372
rect 18690 19360 18696 19372
rect 18472 19332 18696 19360
rect 18472 19320 18478 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19015 19332 19196 19360
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 13556 19298 13691 19301
rect 13556 19292 13584 19298
rect 13372 19264 13584 19292
rect 13633 19295 13691 19298
rect 9674 19224 9680 19236
rect 9508 19196 9680 19224
rect 5224 19184 5230 19196
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 13372 19224 13400 19264
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 13902 19295 13960 19301
rect 13902 19261 13914 19295
rect 13948 19261 13960 19295
rect 19168 19292 19196 19332
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19300 19332 19345 19360
rect 19300 19320 19306 19332
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19668 19332 19717 19360
rect 19668 19320 19674 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 21174 19360 21180 19372
rect 21135 19332 21180 19360
rect 19889 19323 19947 19329
rect 19168 19264 19288 19292
rect 13902 19255 13960 19261
rect 13446 19224 13452 19236
rect 13372 19196 13452 19224
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 4617 19159 4675 19165
rect 4617 19125 4629 19159
rect 4663 19156 4675 19159
rect 4890 19156 4896 19168
rect 4663 19128 4896 19156
rect 4663 19125 4675 19128
rect 4617 19119 4675 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 9766 19156 9772 19168
rect 9727 19128 9772 19156
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10413 19159 10471 19165
rect 10413 19156 10425 19159
rect 10100 19128 10425 19156
rect 10100 19116 10106 19128
rect 10413 19125 10425 19128
rect 10459 19156 10471 19159
rect 10502 19156 10508 19168
rect 10459 19128 10508 19156
rect 10459 19125 10471 19128
rect 10413 19119 10471 19125
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 11882 19156 11888 19168
rect 11843 19128 11888 19156
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12492 19128 12537 19156
rect 12492 19116 12498 19128
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 13740 19156 13768 19255
rect 13924 19224 13952 19255
rect 19260 19224 19288 19264
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19904 19292 19932 19323
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22388 19369 22416 19400
rect 22554 19388 22560 19440
rect 22612 19428 22618 19440
rect 24780 19428 24808 19468
rect 26050 19456 26056 19468
rect 26108 19496 26114 19508
rect 27522 19496 27528 19508
rect 26108 19468 27200 19496
rect 27483 19468 27528 19496
rect 26108 19456 26114 19468
rect 22612 19400 24808 19428
rect 22612 19388 22618 19400
rect 24854 19388 24860 19440
rect 24912 19428 24918 19440
rect 27172 19437 27200 19468
rect 27522 19456 27528 19468
rect 27580 19456 27586 19508
rect 25133 19431 25191 19437
rect 25133 19428 25145 19431
rect 24912 19400 25145 19428
rect 24912 19388 24918 19400
rect 25133 19397 25145 19400
rect 25179 19397 25191 19431
rect 25133 19391 25191 19397
rect 25317 19431 25375 19437
rect 25317 19397 25329 19431
rect 25363 19428 25375 19431
rect 27157 19431 27215 19437
rect 25363 19400 26096 19428
rect 25363 19397 25375 19400
rect 25317 19391 25375 19397
rect 26068 19372 26096 19400
rect 27157 19397 27169 19431
rect 27203 19397 27215 19431
rect 27157 19391 27215 19397
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19360 22431 19363
rect 23569 19363 23627 19369
rect 23569 19360 23581 19363
rect 22419 19332 23581 19360
rect 22419 19329 22431 19332
rect 22373 19323 22431 19329
rect 23569 19329 23581 19332
rect 23615 19329 23627 19363
rect 23569 19323 23627 19329
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 25038 19360 25044 19372
rect 24995 19332 25044 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25866 19360 25872 19372
rect 25827 19332 25872 19360
rect 25866 19320 25872 19332
rect 25924 19320 25930 19372
rect 25961 19363 26019 19369
rect 25961 19329 25973 19363
rect 26007 19329 26019 19363
rect 25961 19323 26019 19329
rect 19392 19264 19932 19292
rect 19392 19252 19398 19264
rect 20806 19252 20812 19304
rect 20864 19292 20870 19304
rect 23014 19292 23020 19304
rect 20864 19264 23020 19292
rect 20864 19252 20870 19264
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23474 19292 23480 19304
rect 23435 19264 23480 19292
rect 23474 19252 23480 19264
rect 23532 19252 23538 19304
rect 24397 19295 24455 19301
rect 24397 19261 24409 19295
rect 24443 19261 24455 19295
rect 24397 19255 24455 19261
rect 21082 19224 21088 19236
rect 13924 19196 14044 19224
rect 19260 19196 21088 19224
rect 14016 19168 14044 19196
rect 21082 19184 21088 19196
rect 21140 19184 21146 19236
rect 22373 19227 22431 19233
rect 22373 19193 22385 19227
rect 22419 19224 22431 19227
rect 24302 19224 24308 19236
rect 22419 19196 24308 19224
rect 22419 19193 22431 19196
rect 22373 19187 22431 19193
rect 24302 19184 24308 19196
rect 24360 19184 24366 19236
rect 24412 19224 24440 19255
rect 24486 19252 24492 19304
rect 24544 19292 24550 19304
rect 25976 19292 26004 19323
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 27172 19360 27200 19391
rect 27338 19388 27344 19440
rect 27396 19437 27402 19440
rect 27396 19431 27415 19437
rect 27403 19397 27415 19431
rect 27396 19391 27415 19397
rect 27396 19388 27402 19391
rect 27890 19360 27896 19372
rect 26108 19332 26201 19360
rect 27172 19332 27896 19360
rect 26108 19320 26114 19332
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 26142 19292 26148 19304
rect 24544 19264 26148 19292
rect 24544 19252 24550 19264
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 25958 19224 25964 19236
rect 24412 19196 25964 19224
rect 25958 19184 25964 19196
rect 26016 19184 26022 19236
rect 13596 19128 13768 19156
rect 13596 19116 13602 19128
rect 13998 19116 14004 19168
rect 14056 19116 14062 19168
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 14332 19128 15761 19156
rect 14332 19116 14338 19128
rect 15749 19125 15761 19128
rect 15795 19125 15807 19159
rect 18966 19156 18972 19168
rect 18927 19128 18972 19156
rect 15749 19119 15807 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 20438 19156 20444 19168
rect 20399 19128 20444 19156
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 20993 19159 21051 19165
rect 20993 19156 21005 19159
rect 20588 19128 21005 19156
rect 20588 19116 20594 19128
rect 20993 19125 21005 19128
rect 21039 19156 21051 19159
rect 23566 19156 23572 19168
rect 21039 19128 23572 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 26234 19156 26240 19168
rect 26195 19128 26240 19156
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 27154 19116 27160 19168
rect 27212 19156 27218 19168
rect 27341 19159 27399 19165
rect 27341 19156 27353 19159
rect 27212 19128 27353 19156
rect 27212 19116 27218 19128
rect 27341 19125 27353 19128
rect 27387 19125 27399 19159
rect 27341 19119 27399 19125
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 5350 18912 5356 18964
rect 5408 18952 5414 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5408 18924 6101 18952
rect 5408 18912 5414 18924
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 6089 18915 6147 18921
rect 7742 18912 7748 18964
rect 7800 18952 7806 18964
rect 13354 18952 13360 18964
rect 7800 18924 13360 18952
rect 7800 18912 7806 18924
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 13504 18924 13645 18952
rect 13504 18912 13510 18924
rect 13633 18921 13645 18924
rect 13679 18952 13691 18955
rect 14642 18952 14648 18964
rect 13679 18924 14648 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 15562 18952 15568 18964
rect 15523 18924 15568 18952
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 18012 18924 18061 18952
rect 18012 18912 18018 18924
rect 18049 18921 18061 18924
rect 18095 18921 18107 18955
rect 18049 18915 18107 18921
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 19886 18952 19892 18964
rect 18748 18924 19892 18952
rect 18748 18912 18754 18924
rect 19886 18912 19892 18924
rect 19944 18952 19950 18964
rect 21637 18955 21695 18961
rect 21637 18952 21649 18955
rect 19944 18924 21649 18952
rect 19944 18912 19950 18924
rect 21637 18921 21649 18924
rect 21683 18921 21695 18955
rect 23937 18955 23995 18961
rect 23937 18952 23949 18955
rect 21637 18915 21695 18921
rect 21744 18924 23949 18952
rect 14550 18844 14556 18896
rect 14608 18884 14614 18896
rect 16577 18887 16635 18893
rect 16577 18884 16589 18887
rect 14608 18856 16589 18884
rect 14608 18844 14614 18856
rect 16577 18853 16589 18856
rect 16623 18853 16635 18887
rect 21744 18884 21772 18924
rect 23937 18921 23949 18924
rect 23983 18921 23995 18955
rect 23937 18915 23995 18921
rect 26697 18955 26755 18961
rect 26697 18921 26709 18955
rect 26743 18952 26755 18955
rect 27338 18952 27344 18964
rect 26743 18924 27344 18952
rect 26743 18921 26755 18924
rect 26697 18915 26755 18921
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 16577 18847 16635 18853
rect 18248 18856 21772 18884
rect 23477 18887 23535 18893
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 15896 18788 17632 18816
rect 15896 18776 15902 18788
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1636 18720 1685 18748
rect 1636 18708 1642 18720
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 4249 18751 4307 18757
rect 4249 18748 4261 18751
rect 4212 18720 4261 18748
rect 4212 18708 4218 18720
rect 4249 18717 4261 18720
rect 4295 18717 4307 18751
rect 4249 18711 4307 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 4982 18757 4988 18760
rect 4976 18711 4988 18757
rect 5040 18748 5046 18760
rect 8297 18751 8355 18757
rect 5040 18720 5076 18748
rect 4982 18708 4988 18711
rect 5040 18708 5046 18720
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 8478 18748 8484 18760
rect 8343 18720 8484 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9548 18720 9597 18748
rect 9548 18708 9554 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 11701 18751 11759 18757
rect 11701 18717 11713 18751
rect 11747 18748 11759 18751
rect 12710 18748 12716 18760
rect 11747 18720 12716 18748
rect 11747 18717 11759 18720
rect 11701 18711 11759 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13688 18720 13737 18748
rect 13688 18708 13694 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 13725 18711 13783 18717
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16632 18720 16681 18748
rect 16632 18708 16638 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17218 18748 17224 18760
rect 16908 18720 17224 18748
rect 16908 18708 16914 18720
rect 17218 18708 17224 18720
rect 17276 18748 17282 18760
rect 17604 18757 17632 18788
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17276 18720 17325 18748
rect 17276 18708 17282 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18248 18757 18276 18856
rect 23477 18853 23489 18887
rect 23523 18884 23535 18887
rect 25038 18884 25044 18896
rect 23523 18856 25044 18884
rect 23523 18853 23535 18856
rect 23477 18847 23535 18853
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 26326 18844 26332 18896
rect 26384 18844 26390 18896
rect 26510 18844 26516 18896
rect 26568 18884 26574 18896
rect 26568 18856 27660 18884
rect 26568 18844 26574 18856
rect 19794 18816 19800 18828
rect 18432 18788 19800 18816
rect 18432 18757 18460 18788
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 20714 18816 20720 18828
rect 20675 18788 20720 18816
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 20898 18776 20904 18828
rect 20956 18816 20962 18828
rect 22833 18819 22891 18825
rect 22833 18816 22845 18819
rect 20956 18788 22845 18816
rect 20956 18776 20962 18788
rect 22833 18785 22845 18788
rect 22879 18816 22891 18819
rect 22879 18788 23520 18816
rect 22879 18785 22891 18788
rect 22833 18779 22891 18785
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 18012 18720 18245 18748
rect 18012 18708 18018 18720
rect 18233 18717 18245 18720
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 18690 18748 18696 18760
rect 18555 18720 18696 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 18932 18720 19625 18748
rect 18932 18708 18938 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19886 18748 19892 18760
rect 19847 18720 19892 18748
rect 19705 18711 19763 18717
rect 9858 18689 9864 18692
rect 9852 18643 9864 18689
rect 9916 18680 9922 18692
rect 11974 18689 11980 18692
rect 9916 18652 9952 18680
rect 9858 18640 9864 18643
rect 9916 18640 9922 18652
rect 11968 18643 11980 18689
rect 12032 18680 12038 18692
rect 12032 18652 12068 18680
rect 11974 18640 11980 18643
rect 12032 18640 12038 18652
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 14274 18680 14280 18692
rect 13044 18652 14280 18680
rect 13044 18640 13050 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 17494 18680 17500 18692
rect 17407 18652 17500 18680
rect 17494 18640 17500 18652
rect 17552 18680 17558 18692
rect 19720 18680 19748 18711
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20806 18748 20812 18760
rect 20036 18720 20081 18748
rect 20767 18720 20812 18748
rect 20036 18708 20042 18720
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 22388 18680 22416 18711
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23014 18748 23020 18760
rect 22796 18720 23020 18748
rect 22796 18708 22802 18720
rect 23014 18708 23020 18720
rect 23072 18748 23078 18760
rect 23492 18757 23520 18788
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 24854 18816 24860 18828
rect 23624 18788 24860 18816
rect 23624 18776 23630 18788
rect 24854 18776 24860 18788
rect 24912 18816 24918 18828
rect 24949 18819 25007 18825
rect 24949 18816 24961 18819
rect 24912 18788 24961 18816
rect 24912 18776 24918 18788
rect 24949 18785 24961 18788
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 26237 18819 26295 18825
rect 25740 18788 26188 18816
rect 25740 18776 25746 18788
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 23072 18720 23305 18748
rect 23072 18708 23078 18720
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18717 23535 18751
rect 23477 18711 23535 18717
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25133 18751 25191 18757
rect 25133 18748 25145 18751
rect 25096 18720 25145 18748
rect 25096 18708 25102 18720
rect 25133 18717 25145 18720
rect 25179 18717 25191 18751
rect 25133 18711 25191 18717
rect 25317 18751 25375 18757
rect 25317 18717 25329 18751
rect 25363 18748 25375 18751
rect 25866 18748 25872 18760
rect 25363 18720 25872 18748
rect 25363 18717 25375 18720
rect 25317 18711 25375 18717
rect 25866 18708 25872 18720
rect 25924 18708 25930 18760
rect 25958 18708 25964 18760
rect 26016 18748 26022 18760
rect 26160 18748 26188 18788
rect 26237 18785 26249 18819
rect 26283 18816 26295 18819
rect 26344 18816 26372 18844
rect 26283 18788 26372 18816
rect 26283 18785 26295 18788
rect 26237 18779 26295 18785
rect 26418 18776 26424 18828
rect 26476 18816 26482 18828
rect 27525 18819 27583 18825
rect 27525 18816 27537 18819
rect 26476 18788 27537 18816
rect 26476 18776 26482 18788
rect 27525 18785 27537 18788
rect 27571 18785 27583 18819
rect 27525 18779 27583 18785
rect 26329 18751 26387 18757
rect 26329 18748 26341 18751
rect 26016 18720 26061 18748
rect 26160 18720 26341 18748
rect 26016 18708 26022 18720
rect 26329 18717 26341 18720
rect 26375 18748 26387 18751
rect 26510 18748 26516 18760
rect 26375 18720 26516 18748
rect 26375 18717 26387 18720
rect 26329 18711 26387 18717
rect 26510 18708 26516 18720
rect 26568 18708 26574 18760
rect 27632 18757 27660 18856
rect 26789 18751 26847 18757
rect 26789 18717 26801 18751
rect 26835 18717 26847 18751
rect 26789 18711 26847 18717
rect 27617 18751 27675 18757
rect 27617 18717 27629 18751
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 23750 18680 23756 18692
rect 17552 18652 19656 18680
rect 19720 18652 20944 18680
rect 17552 18640 17558 18652
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 4062 18612 4068 18624
rect 4023 18584 4068 18612
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 5166 18612 5172 18624
rect 4764 18584 5172 18612
rect 4764 18572 4770 18584
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 7006 18612 7012 18624
rect 6967 18584 7012 18612
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 10226 18612 10232 18624
rect 8536 18584 10232 18612
rect 8536 18572 8542 18584
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10376 18584 10977 18612
rect 10376 18572 10382 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 13081 18615 13139 18621
rect 13081 18581 13093 18615
rect 13127 18612 13139 18615
rect 13446 18612 13452 18624
rect 13127 18584 13452 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 17129 18615 17187 18621
rect 17129 18612 17141 18615
rect 16632 18584 17141 18612
rect 16632 18572 16638 18584
rect 17129 18581 17141 18584
rect 17175 18581 17187 18615
rect 17129 18575 17187 18581
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 19429 18615 19487 18621
rect 19429 18612 19441 18615
rect 19116 18584 19441 18612
rect 19116 18572 19122 18584
rect 19429 18581 19441 18584
rect 19475 18581 19487 18615
rect 19628 18612 19656 18652
rect 20806 18612 20812 18624
rect 19628 18584 20812 18612
rect 19429 18575 19487 18581
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 20916 18612 20944 18652
rect 21109 18652 23756 18680
rect 21109 18612 21137 18652
rect 23750 18640 23756 18652
rect 23808 18680 23814 18692
rect 24486 18680 24492 18692
rect 23808 18652 24492 18680
rect 23808 18640 23814 18652
rect 24486 18640 24492 18652
rect 24544 18640 24550 18692
rect 25774 18640 25780 18692
rect 25832 18680 25838 18692
rect 26050 18680 26056 18692
rect 25832 18652 26056 18680
rect 25832 18640 25838 18652
rect 26050 18640 26056 18652
rect 26108 18680 26114 18692
rect 26804 18680 26832 18711
rect 26108 18652 26832 18680
rect 26108 18640 26114 18652
rect 20916 18584 21137 18612
rect 21177 18615 21235 18621
rect 21177 18581 21189 18615
rect 21223 18612 21235 18615
rect 21542 18612 21548 18624
rect 21223 18584 21548 18612
rect 21223 18581 21235 18584
rect 21177 18575 21235 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 22465 18615 22523 18621
rect 22465 18612 22477 18615
rect 21692 18584 22477 18612
rect 21692 18572 21698 18584
rect 22465 18581 22477 18584
rect 22511 18581 22523 18615
rect 22465 18575 22523 18581
rect 22557 18615 22615 18621
rect 22557 18581 22569 18615
rect 22603 18612 22615 18615
rect 23198 18612 23204 18624
rect 22603 18584 23204 18612
rect 22603 18581 22615 18584
rect 22557 18575 22615 18581
rect 23198 18572 23204 18584
rect 23256 18572 23262 18624
rect 27154 18572 27160 18624
rect 27212 18612 27218 18624
rect 27249 18615 27307 18621
rect 27249 18612 27261 18615
rect 27212 18584 27261 18612
rect 27212 18572 27218 18584
rect 27249 18581 27261 18584
rect 27295 18581 27307 18615
rect 27249 18575 27307 18581
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 5074 18368 5080 18420
rect 5132 18368 5138 18420
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18408 5503 18411
rect 5491 18380 7604 18408
rect 5491 18377 5503 18380
rect 5445 18371 5503 18377
rect 4338 18340 4344 18352
rect 4299 18312 4344 18340
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 5092 18340 5120 18368
rect 4816 18312 5120 18340
rect 7000 18343 7058 18349
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 1949 18275 2007 18281
rect 1949 18241 1961 18275
rect 1995 18272 2007 18275
rect 2222 18272 2228 18284
rect 1995 18244 2228 18272
rect 1995 18241 2007 18244
rect 1949 18235 2007 18241
rect 1780 18204 1808 18235
rect 2222 18232 2228 18244
rect 2280 18272 2286 18284
rect 3878 18272 3884 18284
rect 2280 18244 3884 18272
rect 2280 18232 2286 18244
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 4816 18281 4844 18312
rect 7000 18309 7012 18343
rect 7046 18340 7058 18343
rect 7098 18340 7104 18352
rect 7046 18312 7104 18340
rect 7046 18309 7058 18312
rect 7000 18303 7058 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 7576 18340 7604 18380
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7708 18380 8125 18408
rect 7708 18368 7714 18380
rect 8113 18377 8125 18380
rect 8159 18377 8171 18411
rect 8113 18371 8171 18377
rect 8665 18411 8723 18417
rect 8665 18377 8677 18411
rect 8711 18408 8723 18411
rect 9214 18408 9220 18420
rect 8711 18380 9220 18408
rect 8711 18377 8723 18380
rect 8665 18371 8723 18377
rect 9214 18368 9220 18380
rect 9272 18408 9278 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 9272 18380 10885 18408
rect 9272 18368 9278 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 11974 18408 11980 18420
rect 11931 18380 11980 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 13412 18380 19809 18408
rect 13412 18368 13418 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 20809 18411 20867 18417
rect 20809 18408 20821 18411
rect 19944 18380 20821 18408
rect 19944 18368 19950 18380
rect 20809 18377 20821 18380
rect 20855 18377 20867 18411
rect 20809 18371 20867 18377
rect 21542 18368 21548 18420
rect 21600 18408 21606 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 21600 18380 22201 18408
rect 21600 18368 21606 18380
rect 22189 18377 22201 18380
rect 22235 18377 22247 18411
rect 23566 18408 23572 18420
rect 23527 18380 23572 18408
rect 22189 18371 22247 18377
rect 23566 18368 23572 18380
rect 23624 18368 23630 18420
rect 9033 18343 9091 18349
rect 7576 18312 8984 18340
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18241 4859 18275
rect 4801 18235 4859 18241
rect 4894 18275 4952 18281
rect 4894 18241 4906 18275
rect 4940 18241 4952 18275
rect 5074 18272 5080 18284
rect 5035 18244 5080 18272
rect 4894 18235 4952 18241
rect 3234 18204 3240 18216
rect 1780 18176 3240 18204
rect 3234 18164 3240 18176
rect 3292 18204 3298 18216
rect 4908 18204 4936 18235
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 5350 18281 5356 18284
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18241 5227 18275
rect 5169 18235 5227 18241
rect 5307 18275 5356 18281
rect 5307 18241 5319 18275
rect 5353 18241 5356 18275
rect 5307 18235 5356 18241
rect 5184 18204 5212 18235
rect 5350 18232 5356 18235
rect 5408 18272 5414 18284
rect 7742 18272 7748 18284
rect 5408 18244 7748 18272
rect 5408 18232 5414 18244
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8536 18244 8585 18272
rect 8536 18232 8542 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18241 8907 18275
rect 8956 18272 8984 18312
rect 9033 18309 9045 18343
rect 9079 18340 9091 18343
rect 9738 18343 9796 18349
rect 9738 18340 9750 18343
rect 9079 18312 9750 18340
rect 9079 18309 9091 18312
rect 9033 18303 9091 18309
rect 9738 18309 9750 18312
rect 9784 18309 9796 18343
rect 9738 18303 9796 18309
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 12253 18343 12311 18349
rect 10284 18312 12204 18340
rect 10284 18300 10290 18312
rect 11054 18272 11060 18284
rect 8956 18244 11060 18272
rect 8849 18235 8907 18241
rect 6730 18204 6736 18216
rect 3292 18176 4936 18204
rect 5092 18176 5212 18204
rect 6691 18176 6736 18204
rect 3292 18164 3298 18176
rect 2498 18096 2504 18148
rect 2556 18136 2562 18148
rect 2556 18108 2774 18136
rect 2556 18096 2562 18108
rect 2133 18071 2191 18077
rect 2133 18037 2145 18071
rect 2179 18068 2191 18071
rect 2222 18068 2228 18080
rect 2179 18040 2228 18068
rect 2179 18037 2191 18040
rect 2133 18031 2191 18037
rect 2222 18028 2228 18040
rect 2280 18028 2286 18080
rect 2746 18068 2774 18108
rect 3326 18096 3332 18148
rect 3384 18136 3390 18148
rect 5092 18136 5120 18176
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 8864 18204 8892 18235
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11238 18232 11244 18284
rect 11296 18272 11302 18284
rect 11974 18272 11980 18284
rect 11296 18244 11980 18272
rect 11296 18232 11302 18244
rect 11974 18232 11980 18244
rect 12032 18272 12038 18284
rect 12069 18275 12127 18281
rect 12069 18272 12081 18275
rect 12032 18244 12081 18272
rect 12032 18232 12038 18244
rect 12069 18241 12081 18244
rect 12115 18241 12127 18275
rect 12176 18272 12204 18312
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 13446 18340 13452 18352
rect 12299 18312 13452 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 13446 18300 13452 18312
rect 13504 18300 13510 18352
rect 14734 18340 14740 18352
rect 14695 18312 14740 18340
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15749 18343 15807 18349
rect 15749 18309 15761 18343
rect 15795 18340 15807 18343
rect 16117 18343 16175 18349
rect 15795 18312 16073 18340
rect 15795 18309 15807 18312
rect 15749 18303 15807 18309
rect 12342 18272 12348 18284
rect 12176 18244 12348 18272
rect 12069 18235 12127 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18272 13047 18275
rect 15194 18272 15200 18284
rect 13035 18244 15200 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15396 18244 15669 18272
rect 8938 18204 8944 18216
rect 8864 18176 8944 18204
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9490 18204 9496 18216
rect 9272 18176 9496 18204
rect 9272 18164 9278 18176
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 10870 18204 10876 18216
rect 10560 18176 10876 18204
rect 10560 18164 10566 18176
rect 10870 18164 10876 18176
rect 10928 18204 10934 18216
rect 10928 18176 14044 18204
rect 10928 18164 10934 18176
rect 3384 18108 5120 18136
rect 3384 18096 3390 18108
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 9030 18136 9036 18148
rect 7984 18108 9036 18136
rect 7984 18096 7990 18108
rect 9030 18096 9036 18108
rect 9088 18096 9094 18148
rect 14016 18136 14044 18176
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 15396 18204 15424 18244
rect 15657 18241 15669 18244
rect 15703 18272 15715 18275
rect 15838 18272 15844 18284
rect 15703 18244 15844 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 16045 18272 16073 18312
rect 16117 18309 16129 18343
rect 16163 18340 16175 18343
rect 17098 18343 17156 18349
rect 17098 18340 17110 18343
rect 16163 18312 17110 18340
rect 16163 18309 16175 18312
rect 16117 18303 16175 18309
rect 17098 18309 17110 18312
rect 17144 18309 17156 18343
rect 19518 18340 19524 18352
rect 17098 18303 17156 18309
rect 19168 18312 19524 18340
rect 17862 18272 17868 18284
rect 16045 18244 17868 18272
rect 15933 18235 15991 18241
rect 14148 18176 15424 18204
rect 14148 18164 14154 18176
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 15948 18204 15976 18235
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18874 18272 18880 18284
rect 18196 18244 18880 18272
rect 18196 18232 18202 18244
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19168 18281 19196 18312
rect 19518 18300 19524 18312
rect 19576 18300 19582 18352
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18272 19303 18275
rect 19889 18275 19947 18281
rect 19291 18244 19472 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 15804 18176 15976 18204
rect 15804 18164 15810 18176
rect 14550 18136 14556 18148
rect 14016 18108 14556 18136
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 15948 18136 15976 18176
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 16080 18176 16865 18204
rect 16080 18164 16086 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 18690 18204 18696 18216
rect 16853 18167 16911 18173
rect 18064 18176 18276 18204
rect 18651 18176 18696 18204
rect 16758 18136 16764 18148
rect 15948 18108 16764 18136
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 18064 18136 18092 18176
rect 17788 18108 18092 18136
rect 18248 18136 18276 18176
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 18984 18204 19012 18235
rect 19334 18204 19340 18216
rect 18984 18176 19340 18204
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19444 18136 19472 18244
rect 19889 18241 19901 18275
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 20073 18275 20131 18281
rect 20073 18241 20085 18275
rect 20119 18272 20131 18275
rect 20162 18272 20168 18284
rect 20119 18244 20168 18272
rect 20119 18241 20131 18244
rect 20073 18235 20131 18241
rect 19904 18204 19932 18235
rect 20162 18232 20168 18244
rect 20220 18272 20226 18284
rect 20993 18275 21051 18281
rect 20220 18244 20944 18272
rect 20220 18232 20226 18244
rect 20714 18204 20720 18216
rect 19904 18176 20720 18204
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 18248 18108 19472 18136
rect 20916 18136 20944 18244
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21082 18272 21088 18284
rect 21039 18244 21088 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 21266 18272 21272 18284
rect 21227 18244 21272 18272
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18272 21511 18275
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21499 18244 22017 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18241 22339 18275
rect 22281 18235 22339 18241
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 22296 18204 22324 18235
rect 22370 18232 22376 18284
rect 22428 18272 22434 18284
rect 23198 18272 23204 18284
rect 22428 18244 22473 18272
rect 23159 18244 23204 18272
rect 22428 18232 22434 18244
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 23569 18275 23627 18281
rect 23569 18241 23581 18275
rect 23615 18272 23627 18275
rect 25038 18272 25044 18284
rect 23615 18244 25044 18272
rect 23615 18241 23627 18244
rect 23569 18235 23627 18241
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25958 18232 25964 18284
rect 26016 18272 26022 18284
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 26016 18244 26157 18272
rect 26016 18232 26022 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 26145 18235 26203 18241
rect 26326 18232 26332 18284
rect 26384 18272 26390 18284
rect 27341 18275 27399 18281
rect 27341 18272 27353 18275
rect 26384 18244 27353 18272
rect 26384 18232 26390 18244
rect 27341 18241 27353 18244
rect 27387 18241 27399 18275
rect 27341 18235 27399 18241
rect 23750 18204 23756 18216
rect 21692 18176 22324 18204
rect 23711 18176 23756 18204
rect 21692 18164 21698 18176
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 25590 18204 25596 18216
rect 25551 18176 25596 18204
rect 25590 18164 25596 18176
rect 25648 18164 25654 18216
rect 26234 18204 26240 18216
rect 26195 18176 26240 18204
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 27246 18204 27252 18216
rect 27207 18176 27252 18204
rect 27246 18164 27252 18176
rect 27304 18164 27310 18216
rect 20916 18108 22094 18136
rect 5905 18071 5963 18077
rect 5905 18068 5917 18071
rect 2746 18040 5917 18068
rect 5905 18037 5917 18040
rect 5951 18068 5963 18071
rect 9398 18068 9404 18080
rect 5951 18040 9404 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 17788 18068 17816 18108
rect 9824 18040 17816 18068
rect 9824 18028 9830 18040
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 17920 18040 18245 18068
rect 17920 18028 17926 18040
rect 18233 18037 18245 18040
rect 18279 18068 18291 18071
rect 21174 18068 21180 18080
rect 18279 18040 21180 18068
rect 18279 18037 18291 18040
rect 18233 18031 18291 18037
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 22066 18068 22094 18108
rect 22278 18096 22284 18148
rect 22336 18136 22342 18148
rect 22557 18139 22615 18145
rect 22557 18136 22569 18139
rect 22336 18108 22569 18136
rect 22336 18096 22342 18108
rect 22557 18105 22569 18108
rect 22603 18105 22615 18139
rect 24765 18139 24823 18145
rect 24765 18136 24777 18139
rect 22557 18099 22615 18105
rect 23400 18108 24777 18136
rect 23400 18068 23428 18108
rect 24765 18105 24777 18108
rect 24811 18105 24823 18139
rect 24765 18099 24823 18105
rect 27709 18139 27767 18145
rect 27709 18105 27721 18139
rect 27755 18136 27767 18139
rect 27890 18136 27896 18148
rect 27755 18108 27896 18136
rect 27755 18105 27767 18108
rect 27709 18099 27767 18105
rect 27890 18096 27896 18108
rect 27948 18096 27954 18148
rect 24302 18068 24308 18080
rect 22066 18040 23428 18068
rect 24263 18040 24308 18068
rect 24302 18028 24308 18040
rect 24360 18028 24366 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 6730 17864 6736 17876
rect 6691 17836 6736 17864
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 8386 17864 8392 17876
rect 6840 17836 8392 17864
rect 3436 17728 3464 17824
rect 5902 17756 5908 17808
rect 5960 17796 5966 17808
rect 6840 17796 6868 17836
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 10962 17864 10968 17876
rect 9180 17836 10968 17864
rect 9180 17824 9186 17836
rect 10962 17824 10968 17836
rect 11020 17864 11026 17876
rect 13078 17864 13084 17876
rect 11020 17836 13084 17864
rect 11020 17824 11026 17836
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 13722 17864 13728 17876
rect 13683 17836 13728 17864
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 18230 17864 18236 17876
rect 15252 17836 18236 17864
rect 15252 17824 15258 17836
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21545 17867 21603 17873
rect 21545 17864 21557 17867
rect 21324 17836 21557 17864
rect 21324 17824 21330 17836
rect 21545 17833 21557 17836
rect 21591 17833 21603 17867
rect 25682 17864 25688 17876
rect 21545 17827 21603 17833
rect 22664 17836 25688 17864
rect 8570 17796 8576 17808
rect 5960 17768 6868 17796
rect 7852 17768 8576 17796
rect 5960 17756 5966 17768
rect 3436 17700 4292 17728
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2130 17660 2136 17672
rect 2087 17632 2136 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2314 17669 2320 17672
rect 2308 17660 2320 17669
rect 2275 17632 2320 17660
rect 2308 17623 2320 17632
rect 2314 17620 2320 17623
rect 2372 17620 2378 17672
rect 3970 17660 3976 17672
rect 3931 17632 3976 17660
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 4264 17669 4292 17700
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17629 4307 17663
rect 4249 17623 4307 17629
rect 4338 17620 4344 17672
rect 4396 17660 4402 17672
rect 5350 17660 5356 17672
rect 4396 17632 5356 17660
rect 4396 17620 4402 17632
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17660 7711 17663
rect 7852 17660 7880 17768
rect 8570 17756 8576 17768
rect 8628 17756 8634 17808
rect 9769 17799 9827 17805
rect 9769 17765 9781 17799
rect 9815 17796 9827 17799
rect 9858 17796 9864 17808
rect 9815 17768 9864 17796
rect 9815 17765 9827 17768
rect 9769 17759 9827 17765
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 16577 17799 16635 17805
rect 16577 17796 16589 17799
rect 13228 17768 16589 17796
rect 13228 17756 13234 17768
rect 16577 17765 16589 17768
rect 16623 17765 16635 17799
rect 16577 17759 16635 17765
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 16724 17768 19472 17796
rect 16724 17756 16730 17768
rect 9217 17731 9275 17737
rect 9217 17697 9229 17731
rect 9263 17728 9275 17731
rect 9263 17700 11192 17728
rect 9263 17697 9275 17700
rect 9217 17691 9275 17697
rect 9784 17672 9812 17700
rect 7699 17632 7880 17660
rect 7699 17629 7711 17632
rect 7653 17623 7711 17629
rect 7926 17620 7932 17672
rect 7984 17660 7990 17672
rect 8386 17660 8392 17672
rect 7984 17632 8029 17660
rect 8347 17632 8392 17660
rect 7984 17620 7990 17632
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 4157 17595 4215 17601
rect 4157 17561 4169 17595
rect 4203 17592 4215 17595
rect 5074 17592 5080 17604
rect 4203 17564 5080 17592
rect 4203 17561 4215 17564
rect 4157 17555 4215 17561
rect 4356 17536 4384 17564
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5261 17595 5319 17601
rect 5261 17561 5273 17595
rect 5307 17592 5319 17595
rect 7006 17592 7012 17604
rect 5307 17564 7012 17592
rect 5307 17561 5319 17564
rect 5261 17555 5319 17561
rect 7006 17552 7012 17564
rect 7064 17552 7070 17604
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 7837 17595 7895 17601
rect 7837 17592 7849 17595
rect 7800 17564 7849 17592
rect 7800 17552 7806 17564
rect 7837 17561 7849 17564
rect 7883 17561 7895 17595
rect 8588 17592 8616 17623
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8904 17632 9137 17660
rect 8904 17620 8910 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9306 17660 9312 17672
rect 9267 17632 9312 17660
rect 9125 17623 9183 17629
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9916 17632 9965 17660
rect 9916 17620 9922 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 10226 17660 10232 17672
rect 10187 17632 10232 17660
rect 9953 17623 10011 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 10137 17595 10195 17601
rect 8588 17564 9352 17592
rect 7837 17555 7895 17561
rect 4338 17484 4344 17536
rect 4396 17484 4402 17536
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 6454 17524 6460 17536
rect 4571 17496 6460 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 7248 17496 7481 17524
rect 7248 17484 7254 17496
rect 7469 17493 7481 17496
rect 7515 17493 7527 17527
rect 7469 17487 7527 17493
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8352 17496 8493 17524
rect 8352 17484 8358 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 9324 17524 9352 17564
rect 10137 17561 10149 17595
rect 10183 17592 10195 17595
rect 10318 17592 10324 17604
rect 10183 17564 10324 17592
rect 10183 17561 10195 17564
rect 10137 17555 10195 17561
rect 10318 17552 10324 17564
rect 10376 17552 10382 17604
rect 11164 17592 11192 17700
rect 16758 17688 16764 17740
rect 16816 17728 16822 17740
rect 17497 17731 17555 17737
rect 17497 17728 17509 17731
rect 16816 17700 17509 17728
rect 16816 17688 16822 17700
rect 17497 17697 17509 17700
rect 17543 17728 17555 17731
rect 17586 17728 17592 17740
rect 17543 17700 17592 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 17586 17688 17592 17700
rect 17644 17728 17650 17740
rect 17954 17728 17960 17740
rect 17644 17700 17960 17728
rect 17644 17688 17650 17700
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 18966 17728 18972 17740
rect 18248 17700 18972 17728
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12437 17663 12495 17669
rect 12437 17660 12449 17663
rect 11940 17632 12449 17660
rect 11940 17620 11946 17632
rect 12437 17629 12449 17632
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13136 17632 13185 17660
rect 13136 17620 13142 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13538 17660 13544 17672
rect 13499 17632 13544 17660
rect 13173 17623 13231 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13648 17632 14289 17660
rect 12158 17592 12164 17604
rect 11164 17564 12164 17592
rect 12158 17552 12164 17564
rect 12216 17592 12222 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 12216 17564 13369 17592
rect 12216 17552 12222 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 13504 17564 13549 17592
rect 13504 17552 13510 17564
rect 10226 17524 10232 17536
rect 9324 17496 10232 17524
rect 8481 17487 8539 17493
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 11146 17524 11152 17536
rect 11107 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 13262 17524 13268 17536
rect 12400 17496 13268 17524
rect 12400 17484 12406 17496
rect 13262 17484 13268 17496
rect 13320 17524 13326 17536
rect 13648 17524 13676 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 18248 17669 18276 17700
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 19444 17737 19472 17768
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 20438 17796 20444 17808
rect 19576 17768 20444 17796
rect 19576 17756 19582 17768
rect 20438 17756 20444 17768
rect 20496 17756 20502 17808
rect 21358 17756 21364 17808
rect 21416 17796 21422 17808
rect 21416 17768 22324 17796
rect 21416 17756 21422 17768
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 20530 17728 20536 17740
rect 19475 17700 20536 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 21266 17688 21272 17740
rect 21324 17728 21330 17740
rect 21450 17728 21456 17740
rect 21324 17700 21456 17728
rect 21324 17688 21330 17700
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 22296 17728 22324 17768
rect 22664 17728 22692 17836
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 25958 17864 25964 17876
rect 25919 17836 25964 17864
rect 25958 17824 25964 17836
rect 26016 17824 26022 17876
rect 26053 17867 26111 17873
rect 26053 17833 26065 17867
rect 26099 17864 26111 17867
rect 26418 17864 26424 17876
rect 26099 17836 26424 17864
rect 26099 17833 26111 17836
rect 26053 17827 26111 17833
rect 26418 17824 26424 17836
rect 26476 17824 26482 17876
rect 27065 17867 27123 17873
rect 27065 17833 27077 17867
rect 27111 17864 27123 17867
rect 27246 17864 27252 17876
rect 27111 17836 27252 17864
rect 27111 17833 27123 17836
rect 27065 17827 27123 17833
rect 27246 17824 27252 17836
rect 27304 17824 27310 17876
rect 23477 17799 23535 17805
rect 23477 17765 23489 17799
rect 23523 17765 23535 17799
rect 23477 17759 23535 17765
rect 23492 17728 23520 17759
rect 22296 17700 22692 17728
rect 18233 17663 18291 17669
rect 14608 17632 17632 17660
rect 14608 17620 14614 17632
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 15286 17592 15292 17604
rect 13872 17564 14872 17592
rect 15247 17564 15292 17592
rect 13872 17552 13878 17564
rect 13320 17496 13676 17524
rect 13320 17484 13326 17496
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 14056 17496 14381 17524
rect 14056 17484 14062 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14734 17524 14740 17536
rect 14695 17496 14740 17524
rect 14369 17487 14427 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 14844 17524 14872 17564
rect 15286 17552 15292 17564
rect 15344 17552 15350 17604
rect 17402 17524 17408 17536
rect 14844 17496 17408 17524
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 17604 17524 17632 17632
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18322 17620 18328 17672
rect 18380 17660 18386 17672
rect 18601 17663 18659 17669
rect 18380 17632 18425 17660
rect 18380 17620 18386 17632
rect 18601 17629 18613 17663
rect 18647 17660 18659 17663
rect 18690 17660 18696 17672
rect 18647 17632 18696 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19610 17660 19616 17672
rect 19571 17632 19616 17660
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20625 17663 20683 17669
rect 20625 17660 20637 17663
rect 20128 17632 20637 17660
rect 20128 17620 20134 17632
rect 20625 17629 20637 17632
rect 20671 17629 20683 17663
rect 21542 17660 21548 17672
rect 21503 17632 21548 17660
rect 20625 17623 20683 17629
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 21949 17663 22007 17669
rect 21949 17629 21961 17663
rect 21995 17660 22007 17663
rect 22186 17660 22192 17672
rect 21995 17632 22192 17660
rect 21995 17629 22007 17632
rect 21949 17623 22007 17629
rect 22186 17620 22192 17632
rect 22244 17660 22250 17672
rect 22370 17660 22376 17672
rect 22244 17632 22376 17660
rect 22244 17620 22250 17632
rect 22370 17620 22376 17632
rect 22428 17660 22434 17672
rect 22664 17669 22692 17700
rect 22940 17700 23520 17728
rect 23753 17731 23811 17737
rect 22940 17669 22968 17700
rect 23753 17697 23765 17731
rect 23799 17728 23811 17731
rect 23842 17728 23848 17740
rect 23799 17700 23848 17728
rect 23799 17697 23811 17700
rect 23753 17691 23811 17697
rect 23842 17688 23848 17700
rect 23900 17728 23906 17740
rect 24673 17731 24731 17737
rect 24673 17728 24685 17731
rect 23900 17700 24685 17728
rect 23900 17688 23906 17700
rect 24673 17697 24685 17700
rect 24719 17697 24731 17731
rect 24673 17691 24731 17697
rect 25774 17688 25780 17740
rect 25832 17728 25838 17740
rect 26145 17731 26203 17737
rect 26145 17728 26157 17731
rect 25832 17700 26157 17728
rect 25832 17688 25838 17700
rect 26145 17697 26157 17700
rect 26191 17697 26203 17731
rect 26145 17691 26203 17697
rect 22649 17663 22707 17669
rect 22428 17632 22600 17660
rect 22428 17620 22434 17632
rect 18782 17592 18788 17604
rect 18743 17564 18788 17592
rect 18782 17552 18788 17564
rect 18840 17552 18846 17604
rect 18874 17552 18880 17604
rect 18932 17592 18938 17604
rect 19150 17592 19156 17604
rect 18932 17564 19156 17592
rect 18932 17552 18938 17564
rect 19150 17552 19156 17564
rect 19208 17552 19214 17604
rect 19628 17592 19656 17620
rect 20257 17595 20315 17601
rect 20257 17592 20269 17595
rect 19628 17564 20269 17592
rect 20257 17561 20269 17564
rect 20303 17561 20315 17595
rect 20257 17555 20315 17561
rect 20441 17595 20499 17601
rect 20441 17561 20453 17595
rect 20487 17592 20499 17595
rect 20530 17592 20536 17604
rect 20487 17564 20536 17592
rect 20487 17561 20499 17564
rect 20441 17555 20499 17561
rect 20530 17552 20536 17564
rect 20588 17552 20594 17604
rect 21729 17595 21787 17601
rect 21729 17592 21741 17595
rect 21560 17564 21741 17592
rect 21560 17536 21588 17564
rect 21729 17561 21741 17564
rect 21775 17561 21787 17595
rect 21729 17555 21787 17561
rect 21821 17595 21879 17601
rect 21821 17561 21833 17595
rect 21867 17592 21879 17595
rect 22278 17592 22284 17604
rect 21867 17564 22284 17592
rect 21867 17561 21879 17564
rect 21821 17555 21879 17561
rect 22278 17552 22284 17564
rect 22336 17552 22342 17604
rect 22572 17592 22600 17632
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17629 22983 17663
rect 23382 17660 23388 17672
rect 23343 17632 23388 17660
rect 22925 17623 22983 17629
rect 22940 17592 22968 17623
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24581 17623 24639 17629
rect 22572 17564 22968 17592
rect 23477 17595 23535 17601
rect 23477 17561 23489 17595
rect 23523 17592 23535 17595
rect 23750 17592 23756 17604
rect 23523 17564 23756 17592
rect 23523 17561 23535 17564
rect 23477 17555 23535 17561
rect 23750 17552 23756 17564
rect 23808 17552 23814 17604
rect 24596 17592 24624 17623
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25866 17660 25872 17672
rect 25827 17632 25872 17660
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 26234 17620 26240 17672
rect 26292 17660 26298 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26292 17632 26985 17660
rect 26292 17620 26298 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 27154 17660 27160 17672
rect 27115 17632 27160 17660
rect 26973 17623 27031 17629
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 24854 17592 24860 17604
rect 24596 17564 24860 17592
rect 24854 17552 24860 17564
rect 24912 17552 24918 17604
rect 19518 17524 19524 17536
rect 17604 17496 19524 17524
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20346 17524 20352 17536
rect 19843 17496 20352 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 21542 17484 21548 17536
rect 21600 17484 21606 17536
rect 22462 17524 22468 17536
rect 22423 17496 22468 17524
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 22830 17524 22836 17536
rect 22791 17496 22836 17524
rect 22830 17484 22836 17496
rect 22888 17484 22894 17536
rect 23566 17524 23572 17536
rect 23527 17496 23572 17524
rect 23566 17484 23572 17496
rect 23624 17524 23630 17536
rect 23934 17524 23940 17536
rect 23624 17496 23940 17524
rect 23624 17484 23630 17496
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 8386 17320 8392 17332
rect 1719 17292 8392 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 8386 17280 8392 17292
rect 8444 17320 8450 17332
rect 11057 17323 11115 17329
rect 8444 17292 10732 17320
rect 8444 17280 8450 17292
rect 2400 17255 2458 17261
rect 2400 17221 2412 17255
rect 2446 17252 2458 17255
rect 2774 17252 2780 17264
rect 2446 17224 2780 17252
rect 2446 17221 2458 17224
rect 2400 17215 2458 17221
rect 2774 17212 2780 17224
rect 2832 17212 2838 17264
rect 5626 17252 5632 17264
rect 3988 17224 5632 17252
rect 3988 17193 4016 17224
rect 5626 17212 5632 17224
rect 5684 17212 5690 17264
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 10704 17261 10732 17292
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11698 17320 11704 17332
rect 11103 17292 11704 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 12529 17323 12587 17329
rect 11808 17292 12434 17320
rect 10689 17255 10747 17261
rect 6512 17224 10364 17252
rect 6512 17212 6518 17224
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17153 4031 17187
rect 3973 17147 4031 17153
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17184 4675 17187
rect 4706 17184 4712 17196
rect 4663 17156 4712 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 4890 17193 4896 17196
rect 4884 17184 4896 17193
rect 4851 17156 4896 17184
rect 4884 17147 4896 17156
rect 4890 17144 4896 17147
rect 4948 17144 4954 17196
rect 6546 17184 6552 17196
rect 6507 17156 6552 17184
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6642 17187 6700 17193
rect 6642 17153 6654 17187
rect 6688 17153 6700 17187
rect 6822 17184 6828 17196
rect 6783 17156 6828 17184
rect 6642 17147 6700 17153
rect 2130 17116 2136 17128
rect 2091 17088 2136 17116
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 6656 17116 6684 17147
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7055 17187 7113 17193
rect 6972 17156 7017 17184
rect 6972 17144 6978 17156
rect 7055 17153 7067 17187
rect 7101 17184 7113 17187
rect 7650 17184 7656 17196
rect 7101 17156 7656 17184
rect 7101 17153 7113 17156
rect 7055 17147 7113 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7800 17156 7849 17184
rect 7800 17144 7806 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9950 17184 9956 17196
rect 9364 17156 9956 17184
rect 9364 17144 9370 17156
rect 9950 17144 9956 17156
rect 10008 17184 10014 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 10008 17156 10057 17184
rect 10008 17144 10014 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 10045 17147 10103 17153
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 10336 17184 10364 17224
rect 10689 17221 10701 17255
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 10778 17212 10784 17264
rect 10836 17252 10842 17264
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 10836 17224 10885 17252
rect 10836 17212 10842 17224
rect 10873 17221 10885 17224
rect 10919 17252 10931 17255
rect 11808 17252 11836 17292
rect 12158 17252 12164 17264
rect 10919 17224 11836 17252
rect 12119 17224 12164 17252
rect 10919 17221 10931 17224
rect 10873 17215 10931 17221
rect 12158 17212 12164 17224
rect 12216 17212 12222 17264
rect 11885 17187 11943 17193
rect 11885 17184 11897 17187
rect 10336 17156 11897 17184
rect 11885 17153 11897 17156
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 11978 17187 12036 17193
rect 11978 17153 11990 17187
rect 12024 17153 12036 17187
rect 11978 17147 12036 17153
rect 6012 17088 6684 17116
rect 6012 17060 6040 17088
rect 3510 17048 3516 17060
rect 3471 17020 3516 17048
rect 3510 17008 3516 17020
rect 3568 17008 3574 17060
rect 5994 17048 6000 17060
rect 5955 17020 6000 17048
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 7193 17051 7251 17057
rect 7193 17017 7205 17051
rect 7239 17048 7251 17051
rect 7282 17048 7288 17060
rect 7239 17020 7288 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 9122 17048 9128 17060
rect 9083 17020 9128 17048
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 9732 17020 10057 17048
rect 9732 17008 9738 17020
rect 10045 17017 10057 17020
rect 10091 17048 10103 17051
rect 10410 17048 10416 17060
rect 10091 17020 10416 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10410 17008 10416 17020
rect 10468 17048 10474 17060
rect 10778 17048 10784 17060
rect 10468 17020 10784 17048
rect 10468 17008 10474 17020
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 5350 16980 5356 16992
rect 4203 16952 5356 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 10594 16980 10600 16992
rect 9456 16952 10600 16980
rect 9456 16940 9462 16952
rect 10594 16940 10600 16952
rect 10652 16980 10658 16992
rect 10873 16983 10931 16989
rect 10873 16980 10885 16983
rect 10652 16952 10885 16980
rect 10652 16940 10658 16952
rect 10873 16949 10885 16952
rect 10919 16949 10931 16983
rect 11992 16980 12020 17147
rect 12250 17144 12256 17196
rect 12308 17193 12314 17196
rect 12406 17193 12434 17292
rect 12529 17289 12541 17323
rect 12575 17320 12587 17323
rect 13906 17320 13912 17332
rect 12575 17292 13912 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 15289 17323 15347 17329
rect 15289 17289 15301 17323
rect 15335 17320 15347 17323
rect 15335 17292 19196 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13170 17252 13176 17264
rect 13035 17224 13176 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15764 17224 15945 17252
rect 12308 17184 12319 17193
rect 12391 17187 12449 17193
rect 12308 17156 12353 17184
rect 12308 17147 12319 17156
rect 12391 17153 12403 17187
rect 12437 17184 12449 17187
rect 13538 17184 13544 17196
rect 12437 17156 13544 17184
rect 12437 17153 12449 17156
rect 12391 17147 12449 17153
rect 12308 17144 12314 17147
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 15194 17184 15200 17196
rect 15155 17156 15200 17184
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15764 17184 15792 17224
rect 15933 17221 15945 17224
rect 15979 17252 15991 17255
rect 18690 17252 18696 17264
rect 15979 17224 18696 17252
rect 15979 17221 15991 17224
rect 15933 17215 15991 17221
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 19168 17252 19196 17292
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 19300 17292 19349 17320
rect 19300 17280 19306 17292
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20404 17292 22140 17320
rect 20404 17280 20410 17292
rect 19610 17252 19616 17264
rect 19168 17224 19616 17252
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 21131 17221 21189 17227
rect 15427 17156 15792 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16117 17187 16175 17193
rect 15896 17156 15941 17184
rect 15896 17144 15902 17156
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16206 17184 16212 17196
rect 16163 17156 16212 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 17109 17187 17167 17193
rect 17109 17184 17121 17187
rect 16816 17156 17121 17184
rect 16816 17144 16822 17156
rect 17109 17153 17121 17156
rect 17155 17153 17167 17187
rect 17109 17147 17167 17153
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19886 17184 19892 17196
rect 19107 17156 19892 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 20070 17184 20076 17196
rect 20031 17156 20076 17184
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20346 17184 20352 17196
rect 20307 17156 20352 17184
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 21131 17187 21143 17221
rect 21177 17218 21189 17221
rect 21177 17187 21199 17218
rect 21266 17212 21272 17264
rect 21324 17252 21330 17264
rect 21361 17255 21419 17261
rect 21361 17252 21373 17255
rect 21324 17224 21373 17252
rect 21324 17212 21330 17224
rect 21361 17221 21373 17224
rect 21407 17221 21419 17255
rect 21361 17215 21419 17221
rect 21450 17212 21456 17264
rect 21508 17252 21514 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21508 17224 22017 17252
rect 21508 17212 21514 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22112 17252 22140 17292
rect 22186 17280 22192 17332
rect 22244 17329 22250 17332
rect 22244 17323 22263 17329
rect 22251 17289 22263 17323
rect 22244 17283 22263 17289
rect 22244 17280 22250 17283
rect 22830 17280 22836 17332
rect 22888 17320 22894 17332
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 22888 17292 23489 17320
rect 22888 17280 22894 17292
rect 23477 17289 23489 17292
rect 23523 17289 23535 17323
rect 23477 17283 23535 17289
rect 22646 17252 22652 17264
rect 22112 17224 22652 17252
rect 22005 17215 22063 17221
rect 22646 17212 22652 17224
rect 22704 17212 22710 17264
rect 22925 17255 22983 17261
rect 22925 17221 22937 17255
rect 22971 17252 22983 17255
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 22971 17224 24501 17252
rect 22971 17221 22983 17224
rect 22925 17215 22983 17221
rect 24489 17221 24501 17224
rect 24535 17252 24547 17255
rect 24762 17252 24768 17264
rect 24535 17224 24768 17252
rect 24535 17221 24547 17224
rect 24489 17215 24547 17221
rect 24762 17212 24768 17224
rect 24820 17252 24826 17264
rect 24820 17224 25544 17252
rect 24820 17212 24826 17224
rect 21131 17184 21199 17187
rect 21634 17184 21640 17196
rect 21131 17181 21640 17184
rect 21171 17156 21640 17181
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 21726 17144 21732 17196
rect 21784 17184 21790 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 21784 17156 22845 17184
rect 21784 17144 21790 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 23014 17184 23020 17196
rect 22975 17156 23020 17184
rect 22833 17147 22891 17153
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 23842 17184 23848 17196
rect 23803 17156 23848 17184
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24673 17187 24731 17193
rect 23992 17156 24037 17184
rect 23992 17144 23998 17156
rect 24673 17153 24685 17187
rect 24719 17184 24731 17187
rect 24854 17184 24860 17196
rect 24719 17156 24860 17184
rect 24719 17153 24731 17156
rect 24673 17147 24731 17153
rect 24854 17144 24860 17156
rect 24912 17184 24918 17196
rect 25516 17193 25544 17224
rect 25317 17187 25375 17193
rect 25317 17184 25329 17187
rect 24912 17156 25329 17184
rect 24912 17144 24918 17156
rect 25317 17153 25329 17156
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17184 27307 17187
rect 27338 17184 27344 17196
rect 27295 17156 27344 17184
rect 27295 17153 27307 17156
rect 27249 17147 27307 17153
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17184 27491 17187
rect 27890 17184 27896 17196
rect 27479 17156 27896 17184
rect 27479 17153 27491 17156
rect 27433 17147 27491 17153
rect 27890 17144 27896 17156
rect 27948 17144 27954 17196
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 16022 17116 16028 17128
rect 14783 17088 16028 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15212 17060 15240 17088
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16724 17088 16865 17116
rect 16724 17076 16730 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 19334 17116 19340 17128
rect 19199 17088 19340 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 19334 17076 19340 17088
rect 19392 17116 19398 17128
rect 19794 17116 19800 17128
rect 19392 17088 19800 17116
rect 19392 17076 19398 17088
rect 19794 17076 19800 17088
rect 19852 17076 19858 17128
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17116 20223 17119
rect 21358 17116 21364 17128
rect 20211 17088 21364 17116
rect 20211 17085 20223 17088
rect 20165 17079 20223 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 21652 17116 21680 17144
rect 23382 17116 23388 17128
rect 21652 17088 23388 17116
rect 23382 17076 23388 17088
rect 23440 17116 23446 17128
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23440 17088 23673 17116
rect 23440 17076 23446 17088
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23661 17079 23719 17085
rect 15194 17008 15200 17060
rect 15252 17008 15258 17060
rect 20257 17051 20315 17057
rect 20257 17017 20269 17051
rect 20303 17048 20315 17051
rect 20993 17051 21051 17057
rect 20993 17048 21005 17051
rect 20303 17020 21005 17048
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 20993 17017 21005 17020
rect 21039 17048 21051 17051
rect 21450 17048 21456 17060
rect 21039 17020 21456 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 22278 17048 22284 17060
rect 22191 17020 22284 17048
rect 12158 16980 12164 16992
rect 11992 16952 12164 16980
rect 10873 16943 10931 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 17218 16980 17224 16992
rect 16347 16952 17224 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 18230 16980 18236 16992
rect 18191 16952 18236 16980
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 20533 16983 20591 16989
rect 20533 16949 20545 16983
rect 20579 16980 20591 16983
rect 20806 16980 20812 16992
rect 20579 16952 20812 16980
rect 20579 16949 20591 16952
rect 20533 16943 20591 16949
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 21174 16980 21180 16992
rect 21135 16952 21180 16980
rect 21174 16940 21180 16952
rect 21232 16980 21238 16992
rect 21726 16980 21732 16992
rect 21232 16952 21732 16980
rect 21232 16940 21238 16952
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 22204 16989 22232 17020
rect 22278 17008 22284 17020
rect 22336 17048 22342 17060
rect 22738 17048 22744 17060
rect 22336 17020 22744 17048
rect 22336 17008 22342 17020
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16949 22247 16983
rect 22370 16980 22376 16992
rect 22331 16952 22376 16980
rect 22189 16943 22247 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23676 16980 23704 17079
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 23808 17088 23853 17116
rect 23808 17076 23814 17088
rect 23768 17048 23796 17076
rect 24857 17051 24915 17057
rect 24857 17048 24869 17051
rect 23768 17020 24869 17048
rect 24857 17017 24869 17020
rect 24903 17048 24915 17051
rect 24946 17048 24952 17060
rect 24903 17020 24952 17048
rect 24903 17017 24915 17020
rect 24857 17011 24915 17017
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 24762 16980 24768 16992
rect 23676 16952 24768 16980
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 25682 16980 25688 16992
rect 25643 16952 25688 16980
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 27120 16952 27353 16980
rect 27120 16940 27126 16952
rect 27341 16949 27353 16952
rect 27387 16949 27399 16983
rect 27341 16943 27399 16949
rect 27614 16940 27620 16992
rect 27672 16980 27678 16992
rect 27985 16983 28043 16989
rect 27985 16980 27997 16983
rect 27672 16952 27997 16980
rect 27672 16940 27678 16952
rect 27985 16949 27997 16952
rect 28031 16949 28043 16983
rect 27985 16943 28043 16949
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 5534 16776 5540 16788
rect 5495 16748 5540 16776
rect 5534 16736 5540 16748
rect 5592 16776 5598 16788
rect 5718 16776 5724 16788
rect 5592 16748 5724 16776
rect 5592 16736 5598 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 8754 16776 8760 16788
rect 8435 16748 8760 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 11333 16779 11391 16785
rect 10284 16748 10364 16776
rect 10284 16736 10290 16748
rect 5258 16668 5264 16720
rect 5316 16708 5322 16720
rect 5316 16680 8156 16708
rect 5316 16668 5322 16680
rect 3510 16600 3516 16652
rect 3568 16640 3574 16652
rect 3568 16612 4200 16640
rect 3568 16600 3574 16612
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16572 4031 16575
rect 4172 16572 4200 16612
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 7524 16612 7972 16640
rect 7524 16600 7530 16612
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 4019 16544 4108 16572
rect 4172 16544 4261 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 2308 16507 2366 16513
rect 2308 16473 2320 16507
rect 2354 16504 2366 16507
rect 2682 16504 2688 16516
rect 2354 16476 2688 16504
rect 2354 16473 2366 16476
rect 2308 16467 2366 16473
rect 2682 16464 2688 16476
rect 2740 16464 2746 16516
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 4080 16436 4108 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 6730 16572 6736 16584
rect 4396 16544 4441 16572
rect 5000 16544 6736 16572
rect 4396 16532 4402 16544
rect 4157 16507 4215 16513
rect 4157 16473 4169 16507
rect 4203 16504 4215 16507
rect 4430 16504 4436 16516
rect 4203 16476 4436 16504
rect 4203 16473 4215 16476
rect 4157 16467 4215 16473
rect 4430 16464 4436 16476
rect 4488 16504 4494 16516
rect 5000 16504 5028 16544
rect 6730 16532 6736 16544
rect 6788 16532 6794 16584
rect 7944 16581 7972 16612
rect 8128 16581 8156 16680
rect 9306 16640 9312 16652
rect 9267 16612 9312 16640
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16572 8263 16575
rect 8570 16572 8576 16584
rect 8251 16544 8576 16572
rect 8251 16541 8263 16544
rect 8205 16535 8263 16541
rect 4488 16476 5028 16504
rect 7009 16507 7067 16513
rect 4488 16464 4494 16476
rect 7009 16473 7021 16507
rect 7055 16504 7067 16507
rect 7742 16504 7748 16516
rect 7055 16476 7748 16504
rect 7055 16473 7067 16476
rect 7009 16467 7067 16473
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 7852 16504 7880 16535
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10336 16572 10364 16748
rect 11333 16745 11345 16779
rect 11379 16776 11391 16779
rect 12342 16776 12348 16788
rect 11379 16748 12348 16776
rect 11379 16745 11391 16748
rect 11333 16739 11391 16745
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 13998 16776 14004 16788
rect 12400 16748 14004 16776
rect 12400 16736 12406 16748
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16942 16776 16948 16788
rect 16264 16748 16948 16776
rect 16264 16736 16270 16748
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 18230 16776 18236 16788
rect 17144 16748 18236 16776
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 13725 16711 13783 16717
rect 13725 16708 13737 16711
rect 13688 16680 13737 16708
rect 13688 16668 13694 16680
rect 13725 16677 13737 16680
rect 13771 16677 13783 16711
rect 13725 16671 13783 16677
rect 16390 16668 16396 16720
rect 16448 16708 16454 16720
rect 17144 16708 17172 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 18509 16779 18567 16785
rect 18509 16745 18521 16779
rect 18555 16776 18567 16779
rect 18690 16776 18696 16788
rect 18555 16748 18696 16776
rect 18555 16745 18567 16748
rect 18509 16739 18567 16745
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 21358 16776 21364 16788
rect 21319 16748 21364 16776
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 24581 16779 24639 16785
rect 24581 16776 24593 16779
rect 24360 16748 24593 16776
rect 24360 16736 24366 16748
rect 24581 16745 24593 16748
rect 24627 16745 24639 16779
rect 27798 16776 27804 16788
rect 27759 16748 27804 16776
rect 24581 16739 24639 16745
rect 27798 16736 27804 16748
rect 27856 16736 27862 16788
rect 21082 16708 21088 16720
rect 16448 16680 17172 16708
rect 19628 16680 21088 16708
rect 16448 16668 16454 16680
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15252 16612 15301 16640
rect 15252 16600 15258 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 19628 16649 19656 16680
rect 21082 16668 21088 16680
rect 21140 16708 21146 16720
rect 21266 16708 21272 16720
rect 21140 16680 21272 16708
rect 21140 16668 21146 16680
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 25682 16708 25688 16720
rect 25424 16680 25688 16708
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16724 16612 17141 16640
rect 16724 16600 16730 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20254 16640 20260 16652
rect 19751 16612 20260 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 10192 16544 10364 16572
rect 10192 16532 10198 16544
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 12676 16544 14381 16572
rect 12676 16532 12682 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14550 16572 14556 16584
rect 14511 16544 14556 16572
rect 14369 16535 14427 16541
rect 14550 16532 14556 16544
rect 14608 16572 14614 16584
rect 15556 16575 15614 16581
rect 14608 16544 15516 16572
rect 14608 16532 14614 16544
rect 8478 16504 8484 16516
rect 7852 16476 8484 16504
rect 8478 16464 8484 16476
rect 8536 16464 8542 16516
rect 9576 16507 9634 16513
rect 9576 16473 9588 16507
rect 9622 16504 9634 16507
rect 10042 16504 10048 16516
rect 9622 16476 10048 16504
rect 9622 16473 9634 16476
rect 9576 16467 9634 16473
rect 10042 16464 10048 16476
rect 10100 16464 10106 16516
rect 12468 16507 12526 16513
rect 12468 16473 12480 16507
rect 12514 16504 12526 16507
rect 12514 16476 13308 16504
rect 12514 16473 12526 16476
rect 12468 16467 12526 16473
rect 4338 16436 4344 16448
rect 3467 16408 4344 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 6546 16436 6552 16448
rect 4571 16408 6552 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8938 16436 8944 16448
rect 8352 16408 8944 16436
rect 8352 16396 8358 16408
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 10686 16436 10692 16448
rect 10647 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 13280 16436 13308 16476
rect 13354 16464 13360 16516
rect 13412 16504 13418 16516
rect 13538 16504 13544 16516
rect 13412 16476 13457 16504
rect 13499 16476 13544 16504
rect 13412 16464 13418 16476
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 14734 16504 14740 16516
rect 13648 16476 14740 16504
rect 13648 16436 13676 16476
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 15488 16504 15516 16544
rect 15556 16541 15568 16575
rect 15602 16572 15614 16575
rect 16574 16572 16580 16584
rect 15602 16544 16580 16572
rect 15602 16541 15614 16544
rect 15556 16535 15614 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17385 16575 17443 16581
rect 17385 16572 17397 16575
rect 17276 16544 17397 16572
rect 17276 16532 17282 16544
rect 17385 16541 17397 16544
rect 17431 16541 17443 16575
rect 19628 16572 19656 16603
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 21542 16640 21548 16652
rect 20456 16612 21548 16640
rect 17385 16535 17443 16541
rect 18156 16544 19656 16572
rect 18156 16504 18184 16544
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 20073 16575 20131 16581
rect 20073 16572 20085 16575
rect 19852 16544 20085 16572
rect 19852 16532 19858 16544
rect 20073 16541 20085 16544
rect 20119 16572 20131 16575
rect 20456 16572 20484 16612
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 22462 16640 22468 16652
rect 22112 16612 22468 16640
rect 20119 16544 20484 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 20714 16572 20720 16584
rect 20588 16544 20633 16572
rect 20675 16544 20720 16572
rect 20588 16532 20594 16544
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21634 16572 21640 16584
rect 20864 16544 21496 16572
rect 21595 16544 21640 16572
rect 20864 16532 20870 16544
rect 15488 16476 18184 16504
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 21174 16504 21180 16516
rect 18288 16476 21180 16504
rect 18288 16464 18294 16476
rect 21174 16464 21180 16476
rect 21232 16504 21238 16516
rect 21361 16507 21419 16513
rect 21361 16504 21373 16507
rect 21232 16476 21373 16504
rect 21232 16464 21238 16476
rect 21361 16473 21373 16476
rect 21407 16473 21419 16507
rect 21468 16504 21496 16544
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 22112 16581 22140 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 25424 16649 25452 16680
rect 25682 16668 25688 16680
rect 25740 16668 25746 16720
rect 27893 16711 27951 16717
rect 27893 16677 27905 16711
rect 27939 16677 27951 16711
rect 27893 16671 27951 16677
rect 25409 16643 25467 16649
rect 25409 16609 25421 16643
rect 25455 16609 25467 16643
rect 25590 16640 25596 16652
rect 25551 16612 25596 16640
rect 25409 16603 25467 16609
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 26053 16643 26111 16649
rect 26053 16609 26065 16643
rect 26099 16640 26111 16643
rect 27908 16640 27936 16671
rect 26099 16612 26924 16640
rect 26099 16609 26111 16612
rect 26053 16603 26111 16609
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16541 22155 16575
rect 22370 16572 22376 16584
rect 22331 16544 22376 16572
rect 22097 16535 22155 16541
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 23293 16575 23351 16581
rect 23293 16572 23305 16575
rect 22612 16544 23305 16572
rect 22612 16532 22618 16544
rect 23293 16541 23305 16544
rect 23339 16572 23351 16575
rect 23382 16572 23388 16584
rect 23339 16544 23388 16572
rect 23339 16541 23351 16544
rect 23293 16535 23351 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23474 16532 23480 16584
rect 23532 16572 23538 16584
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 23532 16544 23581 16572
rect 23532 16532 23538 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 23934 16532 23940 16584
rect 23992 16572 23998 16584
rect 24762 16572 24768 16584
rect 23992 16544 24768 16572
rect 23992 16532 23998 16544
rect 24762 16532 24768 16544
rect 24820 16572 24826 16584
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 24820 16544 25329 16572
rect 24820 16532 24826 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16572 25743 16575
rect 25774 16572 25780 16584
rect 25731 16544 25780 16572
rect 25731 16541 25743 16544
rect 25685 16535 25743 16541
rect 25774 16532 25780 16544
rect 25832 16532 25838 16584
rect 26896 16581 26924 16612
rect 27264 16612 27936 16640
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26881 16575 26939 16581
rect 26881 16541 26893 16575
rect 26927 16572 26939 16575
rect 27154 16572 27160 16584
rect 26927 16544 27160 16572
rect 26927 16541 26939 16544
rect 26881 16535 26939 16541
rect 22189 16507 22247 16513
rect 22189 16504 22201 16507
rect 21468 16476 22201 16504
rect 21361 16467 21419 16473
rect 22189 16473 22201 16476
rect 22235 16473 22247 16507
rect 23400 16504 23428 16532
rect 23400 16476 24900 16504
rect 22189 16467 22247 16473
rect 13280 16408 13676 16436
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16436 14611 16439
rect 15286 16436 15292 16448
rect 14599 16408 15292 16436
rect 14599 16405 14611 16408
rect 14553 16399 14611 16405
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 16669 16439 16727 16445
rect 16669 16405 16681 16439
rect 16715 16436 16727 16439
rect 17494 16436 17500 16448
rect 16715 16408 17500 16436
rect 16715 16405 16727 16408
rect 16669 16399 16727 16405
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 19426 16436 19432 16448
rect 19387 16408 19432 16436
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19886 16436 19892 16448
rect 19847 16408 19892 16436
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 19981 16439 20039 16445
rect 19981 16405 19993 16439
rect 20027 16436 20039 16439
rect 20070 16436 20076 16448
rect 20027 16408 20076 16436
rect 20027 16405 20039 16408
rect 19981 16399 20039 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20622 16436 20628 16448
rect 20583 16408 20628 16436
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21545 16439 21603 16445
rect 21545 16436 21557 16439
rect 21048 16408 21557 16436
rect 21048 16396 21054 16408
rect 21545 16405 21557 16408
rect 21591 16405 21603 16439
rect 21545 16399 21603 16405
rect 22274 16439 22332 16445
rect 22274 16405 22286 16439
rect 22320 16436 22332 16439
rect 22738 16436 22744 16448
rect 22320 16408 22744 16436
rect 22320 16405 22332 16408
rect 22274 16399 22332 16405
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 23106 16436 23112 16448
rect 23067 16408 23112 16436
rect 23106 16396 23112 16408
rect 23164 16396 23170 16448
rect 23477 16439 23535 16445
rect 23477 16405 23489 16439
rect 23523 16436 23535 16439
rect 23566 16436 23572 16448
rect 23523 16408 23572 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 24872 16436 24900 16476
rect 24946 16464 24952 16516
rect 25004 16504 25010 16516
rect 26160 16504 26188 16535
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27264 16581 27292 16612
rect 27982 16600 27988 16652
rect 28040 16640 28046 16652
rect 28040 16612 28085 16640
rect 28040 16600 28046 16612
rect 27249 16575 27307 16581
rect 27249 16541 27261 16575
rect 27295 16541 27307 16575
rect 27249 16535 27307 16541
rect 27430 16532 27436 16584
rect 27488 16572 27494 16584
rect 27709 16575 27767 16581
rect 27709 16572 27721 16575
rect 27488 16544 27721 16572
rect 27488 16532 27494 16544
rect 27709 16541 27721 16544
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 26694 16504 26700 16516
rect 25004 16476 26188 16504
rect 26655 16476 26700 16504
rect 25004 16464 25010 16476
rect 26694 16464 26700 16476
rect 26752 16464 26758 16516
rect 26050 16436 26056 16448
rect 24872 16408 26056 16436
rect 26050 16396 26056 16408
rect 26108 16396 26114 16448
rect 26970 16436 26976 16448
rect 26931 16408 26976 16436
rect 26970 16396 26976 16408
rect 27028 16396 27034 16448
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 27120 16408 27165 16436
rect 27120 16396 27126 16408
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2869 16235 2927 16241
rect 2869 16232 2881 16235
rect 2188 16204 2881 16232
rect 2188 16192 2194 16204
rect 2869 16201 2881 16204
rect 2915 16201 2927 16235
rect 2869 16195 2927 16201
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 6880 16204 7512 16232
rect 6880 16192 6886 16204
rect 1581 16167 1639 16173
rect 1581 16133 1593 16167
rect 1627 16164 1639 16167
rect 2958 16164 2964 16176
rect 1627 16136 2964 16164
rect 1627 16133 1639 16136
rect 1581 16127 1639 16133
rect 2958 16124 2964 16136
rect 3016 16124 3022 16176
rect 5997 16167 6055 16173
rect 5997 16133 6009 16167
rect 6043 16164 6055 16167
rect 7374 16164 7380 16176
rect 6043 16136 7380 16164
rect 6043 16133 6055 16136
rect 5997 16127 6055 16133
rect 7374 16124 7380 16136
rect 7432 16124 7438 16176
rect 7484 16164 7512 16204
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 7800 16204 9137 16232
rect 7800 16192 7806 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 12434 16232 12440 16244
rect 10827 16204 12440 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 12768 16204 14289 16232
rect 12768 16192 12774 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 14277 16195 14335 16201
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16758 16232 16764 16244
rect 16163 16204 16764 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 16942 16232 16948 16244
rect 16903 16204 16948 16232
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 21634 16232 21640 16244
rect 18555 16204 21640 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 22649 16235 22707 16241
rect 22649 16201 22661 16235
rect 22695 16232 22707 16235
rect 23106 16232 23112 16244
rect 22695 16204 23112 16232
rect 22695 16201 22707 16204
rect 22649 16195 22707 16201
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 27430 16232 27436 16244
rect 23400 16204 27436 16232
rect 9490 16164 9496 16176
rect 7484 16136 9496 16164
rect 9490 16124 9496 16136
rect 9548 16124 9554 16176
rect 10410 16164 10416 16176
rect 10371 16136 10416 16164
rect 10410 16124 10416 16136
rect 10468 16124 10474 16176
rect 11146 16124 11152 16176
rect 11204 16164 11210 16176
rect 12989 16167 13047 16173
rect 12989 16164 13001 16167
rect 11204 16136 13001 16164
rect 11204 16124 11210 16136
rect 12989 16133 13001 16136
rect 13035 16133 13047 16167
rect 12989 16127 13047 16133
rect 13354 16124 13360 16176
rect 13412 16164 13418 16176
rect 13906 16164 13912 16176
rect 13412 16136 13912 16164
rect 13412 16124 13418 16136
rect 13906 16124 13912 16136
rect 13964 16124 13970 16176
rect 15749 16167 15807 16173
rect 15749 16133 15761 16167
rect 15795 16164 15807 16167
rect 16390 16164 16396 16176
rect 15795 16136 16396 16164
rect 15795 16133 15807 16136
rect 15749 16127 15807 16133
rect 16390 16124 16396 16136
rect 16448 16124 16454 16176
rect 17402 16124 17408 16176
rect 17460 16164 17466 16176
rect 20993 16167 21051 16173
rect 20993 16164 21005 16167
rect 17460 16136 21005 16164
rect 17460 16124 17466 16136
rect 20993 16133 21005 16136
rect 21039 16133 21051 16167
rect 20993 16127 21051 16133
rect 21542 16124 21548 16176
rect 21600 16164 21606 16176
rect 22554 16164 22560 16176
rect 21600 16136 22560 16164
rect 21600 16124 21606 16136
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 22738 16164 22744 16176
rect 22699 16136 22744 16164
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 3786 16056 3792 16108
rect 3844 16096 3850 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 3844 16068 6561 16096
rect 3844 16056 3850 16068
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 6730 16096 6736 16108
rect 6691 16068 6736 16096
rect 6549 16059 6607 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16065 6975 16099
rect 7834 16096 7840 16108
rect 7795 16068 7840 16096
rect 6917 16059 6975 16065
rect 6840 16028 6868 16059
rect 6564 16000 6868 16028
rect 6564 15972 6592 16000
rect 6546 15920 6552 15972
rect 6604 15920 6610 15972
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 6923 15960 6951 16059
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 10134 16096 10140 16108
rect 10095 16068 10140 16096
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10318 16105 10324 16108
rect 10285 16099 10324 16105
rect 10285 16065 10297 16099
rect 10285 16059 10324 16065
rect 10318 16056 10324 16059
rect 10376 16056 10382 16108
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 10643 16099 10701 16105
rect 10560 16068 10605 16096
rect 10560 16056 10566 16068
rect 10643 16065 10655 16099
rect 10689 16096 10701 16099
rect 10778 16096 10784 16108
rect 10689 16068 10784 16096
rect 10689 16065 10701 16068
rect 10643 16059 10701 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11112 16068 11713 16096
rect 11112 16056 11118 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11848 16068 12173 16096
rect 11848 16056 11854 16068
rect 12161 16065 12173 16068
rect 12207 16096 12219 16099
rect 15010 16096 15016 16108
rect 12207 16068 15016 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15838 16096 15844 16108
rect 15703 16068 15844 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16114 16096 16120 16108
rect 15979 16068 16120 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16942 16096 16948 16108
rect 16855 16068 16948 16096
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 13998 16028 14004 16040
rect 10008 16000 14004 16028
rect 10008 15988 10014 16000
rect 13998 15988 14004 16000
rect 14056 16028 14062 16040
rect 14826 16028 14832 16040
rect 14056 16000 14832 16028
rect 14056 15988 14062 16000
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15562 15988 15568 16040
rect 15620 16028 15626 16040
rect 16960 16028 16988 16056
rect 15620 16000 16988 16028
rect 15620 15988 15626 16000
rect 6788 15932 6951 15960
rect 6788 15920 6794 15932
rect 10134 15920 10140 15972
rect 10192 15960 10198 15972
rect 10594 15960 10600 15972
rect 10192 15932 10600 15960
rect 10192 15920 10198 15932
rect 10594 15920 10600 15932
rect 10652 15920 10658 15972
rect 17034 15960 17040 15972
rect 12406 15932 17040 15960
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 4890 15892 4896 15904
rect 4755 15864 4896 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11296 15864 11805 15892
rect 11296 15852 11302 15864
rect 11793 15861 11805 15864
rect 11839 15892 11851 15895
rect 12406 15892 12434 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 17144 15960 17172 16059
rect 17218 16056 17224 16108
rect 17276 16096 17282 16108
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17276 16068 17969 16096
rect 17276 16056 17282 16068
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16065 18475 16099
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 18417 16059 18475 16065
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18138 16028 18144 16040
rect 17920 16000 18144 16028
rect 17920 15988 17926 16000
rect 18138 15988 18144 16000
rect 18196 16028 18202 16040
rect 18432 16028 18460 16059
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19886 16096 19892 16108
rect 19847 16068 19892 16096
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20254 16096 20260 16108
rect 20027 16068 20260 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 21174 16096 21180 16108
rect 21135 16068 21180 16096
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 22462 16096 22468 16108
rect 22423 16068 22468 16096
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 23400 16105 23428 16204
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 27525 16235 27583 16241
rect 27525 16201 27537 16235
rect 27571 16232 27583 16235
rect 27614 16232 27620 16244
rect 27571 16204 27620 16232
rect 27571 16201 27583 16204
rect 27525 16195 27583 16201
rect 27614 16192 27620 16204
rect 27672 16192 27678 16244
rect 24762 16124 24768 16176
rect 24820 16164 24826 16176
rect 24820 16136 25176 16164
rect 24820 16124 24826 16136
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22756 16068 23397 16096
rect 19794 16028 19800 16040
rect 18196 16000 18460 16028
rect 19755 16000 19800 16028
rect 18196 15988 18202 16000
rect 19794 15988 19800 16000
rect 19852 15988 19858 16040
rect 20070 15988 20076 16040
rect 20128 16028 20134 16040
rect 20714 16028 20720 16040
rect 20128 16000 20720 16028
rect 20128 15988 20134 16000
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 21453 16031 21511 16037
rect 21453 15997 21465 16031
rect 21499 16028 21511 16031
rect 21542 16028 21548 16040
rect 21499 16000 21548 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 22756 16028 22784 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23658 16096 23664 16108
rect 23523 16068 23664 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 24946 16096 24952 16108
rect 24907 16068 24952 16096
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 25148 16105 25176 16136
rect 25590 16124 25596 16176
rect 25648 16164 25654 16176
rect 25648 16136 25912 16164
rect 25648 16124 25654 16136
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 25682 16096 25688 16108
rect 25271 16068 25688 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 25884 16105 25912 16136
rect 25958 16124 25964 16176
rect 26016 16164 26022 16176
rect 26053 16167 26111 16173
rect 26053 16164 26065 16167
rect 26016 16136 26065 16164
rect 26016 16124 26022 16136
rect 26053 16133 26065 16136
rect 26099 16164 26111 16167
rect 26602 16164 26608 16176
rect 26099 16136 26608 16164
rect 26099 16133 26111 16136
rect 26053 16127 26111 16133
rect 26602 16124 26608 16136
rect 26660 16124 26666 16176
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16065 25927 16099
rect 25869 16059 25927 16065
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16096 26203 16099
rect 26694 16096 26700 16108
rect 26191 16068 26700 16096
rect 26191 16065 26203 16068
rect 26145 16059 26203 16065
rect 22428 16000 22784 16028
rect 22428 15988 22434 16000
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 22888 16000 23305 16028
rect 22888 15988 22894 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 23569 16031 23627 16037
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 23842 16028 23848 16040
rect 23615 16000 23848 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 23842 15988 23848 16000
rect 23900 16028 23906 16040
rect 23900 16000 24808 16028
rect 23900 15988 23906 16000
rect 20898 15960 20904 15972
rect 17144 15932 20904 15960
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15960 21419 15963
rect 21634 15960 21640 15972
rect 21407 15932 21640 15960
rect 21407 15929 21419 15932
rect 21361 15923 21419 15929
rect 21634 15920 21640 15932
rect 21692 15960 21698 15972
rect 23753 15963 23811 15969
rect 23753 15960 23765 15963
rect 21692 15932 23765 15960
rect 21692 15920 21698 15932
rect 23753 15929 23765 15932
rect 23799 15929 23811 15963
rect 24780 15960 24808 16000
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25958 16028 25964 16040
rect 24912 16000 25964 16028
rect 24912 15988 24918 16000
rect 25958 15988 25964 16000
rect 26016 16028 26022 16040
rect 26160 16028 26188 16059
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 26016 16000 26188 16028
rect 27617 16031 27675 16037
rect 26016 15988 26022 16000
rect 27617 15997 27629 16031
rect 27663 15997 27675 16031
rect 27617 15991 27675 15997
rect 27157 15963 27215 15969
rect 27157 15960 27169 15963
rect 24780 15932 27169 15960
rect 23753 15923 23811 15929
rect 27157 15929 27169 15932
rect 27203 15929 27215 15963
rect 27632 15960 27660 15991
rect 27706 15988 27712 16040
rect 27764 16028 27770 16040
rect 27764 16000 27809 16028
rect 27764 15988 27770 16000
rect 28074 15960 28080 15972
rect 27632 15932 28080 15960
rect 27157 15923 27215 15929
rect 28074 15920 28080 15932
rect 28132 15920 28138 15972
rect 11839 15864 12434 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 14090 15892 14096 15904
rect 13596 15864 14096 15892
rect 13596 15852 13602 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 15896 15864 17785 15892
rect 15896 15852 15902 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 17773 15855 17831 15861
rect 18877 15895 18935 15901
rect 18877 15861 18889 15895
rect 18923 15892 18935 15895
rect 19334 15892 19340 15904
rect 18923 15864 19340 15892
rect 18923 15861 18935 15864
rect 18877 15855 18935 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19702 15892 19708 15904
rect 19659 15864 19708 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 22281 15895 22339 15901
rect 22281 15861 22293 15895
rect 22327 15892 22339 15895
rect 22554 15892 22560 15904
rect 22327 15864 22560 15892
rect 22327 15861 22339 15864
rect 22281 15855 22339 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 22922 15852 22928 15904
rect 22980 15892 22986 15904
rect 24213 15895 24271 15901
rect 24213 15892 24225 15895
rect 22980 15864 24225 15892
rect 22980 15852 22986 15864
rect 24213 15861 24225 15864
rect 24259 15861 24271 15895
rect 24213 15855 24271 15861
rect 24857 15895 24915 15901
rect 24857 15861 24869 15895
rect 24903 15892 24915 15895
rect 24946 15892 24952 15904
rect 24903 15864 24952 15892
rect 24903 15861 24915 15864
rect 24857 15855 24915 15861
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 25685 15895 25743 15901
rect 25685 15861 25697 15895
rect 25731 15892 25743 15895
rect 25774 15892 25780 15904
rect 25731 15864 25780 15892
rect 25731 15861 25743 15864
rect 25685 15855 25743 15861
rect 25774 15852 25780 15864
rect 25832 15852 25838 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 2038 15688 2044 15700
rect 1999 15660 2044 15688
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 8478 15688 8484 15700
rect 8439 15660 8484 15688
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 12618 15688 12624 15700
rect 10919 15660 12624 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14884 15660 15025 15688
rect 14884 15648 14890 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15930 15688 15936 15700
rect 15891 15660 15936 15688
rect 15013 15651 15071 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 20622 15688 20628 15700
rect 16500 15660 20628 15688
rect 7742 15580 7748 15632
rect 7800 15620 7806 15632
rect 7800 15592 8340 15620
rect 7800 15580 7806 15592
rect 4356 15524 4752 15552
rect 4356 15493 4384 15524
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15453 4399 15487
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4341 15447 4399 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4724 15484 4752 15524
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 4856 15524 5273 15552
rect 4856 15512 4862 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 6638 15512 6644 15564
rect 6696 15552 6702 15564
rect 8312 15552 8340 15592
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 16500 15620 16528 15660
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 21361 15691 21419 15697
rect 21361 15688 21373 15691
rect 21232 15660 21373 15688
rect 21232 15648 21238 15660
rect 21361 15657 21373 15660
rect 21407 15657 21419 15691
rect 25130 15688 25136 15700
rect 21361 15651 21419 15657
rect 22066 15660 25136 15688
rect 19702 15620 19708 15632
rect 9548 15592 16528 15620
rect 18156 15592 19564 15620
rect 19663 15592 19708 15620
rect 9548 15580 9554 15592
rect 10686 15552 10692 15564
rect 6696 15524 8248 15552
rect 8312 15524 8345 15552
rect 6696 15512 6702 15524
rect 4982 15484 4988 15496
rect 4724 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 7006 15484 7012 15496
rect 6967 15456 7012 15484
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 8018 15493 8024 15496
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7156 15456 7849 15484
rect 7156 15444 7162 15456
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7985 15487 8024 15493
rect 7985 15453 7997 15487
rect 7985 15447 8024 15453
rect 8018 15444 8024 15447
rect 8076 15444 8082 15496
rect 8220 15493 8248 15524
rect 8317 15493 8345 15524
rect 9233 15524 10692 15552
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8302 15487 8360 15493
rect 8302 15453 8314 15487
rect 8348 15453 8360 15487
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 8302 15447 8360 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9233 15493 9261 15524
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 12912 15524 15240 15552
rect 9218 15487 9276 15493
rect 9218 15453 9230 15487
rect 9264 15453 9276 15487
rect 9590 15487 9648 15493
rect 9590 15484 9602 15487
rect 9218 15447 9276 15453
rect 9324 15456 9602 15484
rect 3326 15416 3332 15428
rect 3287 15388 3332 15416
rect 3326 15376 3332 15388
rect 3384 15376 3390 15428
rect 4433 15419 4491 15425
rect 4433 15385 4445 15419
rect 4479 15416 4491 15419
rect 5442 15416 5448 15428
rect 4479 15388 5448 15416
rect 4479 15385 4491 15388
rect 4433 15379 4491 15385
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 8113 15419 8171 15425
rect 8113 15385 8125 15419
rect 8159 15385 8171 15419
rect 8113 15379 8171 15385
rect 4801 15351 4859 15357
rect 4801 15317 4813 15351
rect 4847 15348 4859 15351
rect 5258 15348 5264 15360
rect 4847 15320 5264 15348
rect 4847 15317 4859 15320
rect 4801 15311 4859 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 8128 15348 8156 15379
rect 8938 15376 8944 15428
rect 8996 15416 9002 15428
rect 9324 15416 9352 15456
rect 9590 15453 9602 15456
rect 9636 15453 9648 15487
rect 9590 15447 9648 15453
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12802 15484 12808 15496
rect 12207 15456 12808 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 8996 15388 9352 15416
rect 9401 15419 9459 15425
rect 8996 15376 9002 15388
rect 9401 15385 9413 15419
rect 9447 15385 9459 15419
rect 9401 15379 9459 15385
rect 9416 15348 9444 15379
rect 9490 15376 9496 15428
rect 9548 15416 9554 15428
rect 9548 15388 9593 15416
rect 9548 15376 9554 15388
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 12912 15416 12940 15524
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15453 13139 15487
rect 13446 15484 13452 15496
rect 13407 15456 13452 15484
rect 13081 15447 13139 15453
rect 13096 15416 13124 15447
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 15212 15493 15240 15524
rect 15104 15487 15162 15493
rect 15104 15484 15116 15487
rect 15068 15456 15116 15484
rect 15068 15444 15074 15456
rect 15104 15453 15116 15456
rect 15150 15453 15162 15487
rect 15104 15447 15162 15453
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15484 15255 15487
rect 16298 15484 16304 15496
rect 15243 15456 16304 15484
rect 15243 15453 15255 15456
rect 15197 15447 15255 15453
rect 11112 15388 12940 15416
rect 13004 15388 13124 15416
rect 13265 15419 13323 15425
rect 11112 15376 11118 15388
rect 13004 15360 13032 15388
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13354 15416 13360 15428
rect 13311 15388 13360 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 15120 15416 15148 15447
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15484 17463 15487
rect 18046 15484 18052 15496
rect 17451 15456 18052 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18156 15493 18184 15592
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 18506 15552 18512 15564
rect 18279 15524 18512 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 19426 15552 19432 15564
rect 19387 15524 19432 15552
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19536 15552 19564 15592
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 22066 15620 22094 15660
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 25682 15648 25688 15700
rect 25740 15688 25746 15700
rect 26513 15691 26571 15697
rect 25740 15660 26096 15688
rect 25740 15648 25746 15660
rect 20272 15592 22094 15620
rect 22281 15623 22339 15629
rect 20070 15552 20076 15564
rect 19536 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 20272 15484 20300 15592
rect 22281 15589 22293 15623
rect 22327 15620 22339 15623
rect 22462 15620 22468 15632
rect 22327 15592 22468 15620
rect 22327 15589 22339 15592
rect 22281 15583 22339 15589
rect 22462 15580 22468 15592
rect 22520 15620 22526 15632
rect 23293 15623 23351 15629
rect 23293 15620 23305 15623
rect 22520 15592 23305 15620
rect 22520 15580 22526 15592
rect 23293 15589 23305 15592
rect 23339 15589 23351 15623
rect 23293 15583 23351 15589
rect 23382 15580 23388 15632
rect 23440 15620 23446 15632
rect 23440 15592 23704 15620
rect 23440 15580 23446 15592
rect 21542 15512 21548 15564
rect 21600 15552 21606 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21600 15524 22109 15552
rect 21600 15512 21606 15524
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 22738 15552 22744 15564
rect 22603 15524 22744 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 22738 15512 22744 15524
rect 22796 15512 22802 15564
rect 23474 15552 23480 15564
rect 23435 15524 23480 15552
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 18463 15456 20300 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 17678 15416 17684 15428
rect 15120 15388 17684 15416
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 18230 15376 18236 15428
rect 18288 15416 18294 15428
rect 18340 15416 18368 15447
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20533 15487 20591 15493
rect 20404 15456 20449 15484
rect 20404 15444 20410 15456
rect 20533 15453 20545 15487
rect 20579 15484 20591 15487
rect 20622 15484 20628 15496
rect 20579 15456 20628 15484
rect 20579 15453 20591 15456
rect 20533 15447 20591 15453
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 21324 15456 21373 15484
rect 21324 15444 21330 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21634 15484 21640 15496
rect 21595 15456 21640 15484
rect 21361 15447 21419 15453
rect 21634 15444 21640 15456
rect 21692 15444 21698 15496
rect 23566 15484 23572 15496
rect 23479 15456 23572 15484
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 23676 15493 23704 15592
rect 25590 15580 25596 15632
rect 25648 15620 25654 15632
rect 25648 15592 26004 15620
rect 25648 15580 25654 15592
rect 24964 15524 25728 15552
rect 24964 15496 24992 15524
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15484 23811 15487
rect 23842 15484 23848 15496
rect 23799 15456 23848 15484
rect 23799 15453 23811 15456
rect 23753 15447 23811 15453
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24946 15484 24952 15496
rect 24907 15456 24952 15484
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 25225 15487 25283 15493
rect 25225 15453 25237 15487
rect 25271 15484 25283 15487
rect 25590 15484 25596 15496
rect 25271 15456 25596 15484
rect 25271 15453 25283 15456
rect 25225 15447 25283 15453
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 25700 15493 25728 15524
rect 25685 15487 25743 15493
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 25685 15447 25743 15453
rect 25774 15444 25780 15496
rect 25832 15484 25838 15496
rect 25976 15493 26004 15592
rect 25961 15487 26019 15493
rect 25832 15456 25877 15484
rect 25832 15444 25838 15456
rect 25961 15453 25973 15487
rect 26007 15453 26019 15487
rect 26068 15484 26096 15660
rect 26513 15657 26525 15691
rect 26559 15688 26571 15691
rect 26970 15688 26976 15700
rect 26559 15660 26976 15688
rect 26559 15657 26571 15660
rect 26513 15651 26571 15657
rect 26970 15648 26976 15660
rect 27028 15648 27034 15700
rect 27525 15691 27583 15697
rect 27525 15657 27537 15691
rect 27571 15688 27583 15691
rect 27706 15688 27712 15700
rect 27571 15660 27712 15688
rect 27571 15657 27583 15660
rect 27525 15651 27583 15657
rect 27706 15648 27712 15660
rect 27764 15648 27770 15700
rect 28074 15688 28080 15700
rect 28035 15660 28080 15688
rect 28074 15648 28080 15660
rect 28132 15648 28138 15700
rect 27338 15552 27344 15564
rect 27299 15524 27344 15552
rect 27338 15512 27344 15524
rect 27396 15512 27402 15564
rect 27614 15512 27620 15564
rect 27672 15552 27678 15564
rect 27672 15524 28304 15552
rect 27672 15512 27678 15524
rect 26421 15487 26479 15493
rect 26421 15484 26433 15487
rect 26068 15456 26433 15484
rect 25961 15447 26019 15453
rect 26421 15453 26433 15456
rect 26467 15453 26479 15487
rect 26602 15484 26608 15496
rect 26563 15456 26608 15484
rect 26421 15447 26479 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 27249 15487 27307 15493
rect 27249 15484 27261 15487
rect 26712 15456 27261 15484
rect 18288 15388 18368 15416
rect 18288 15376 18294 15388
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 20441 15419 20499 15425
rect 20441 15416 20453 15419
rect 18840 15388 20453 15416
rect 18840 15376 18846 15388
rect 20441 15385 20453 15388
rect 20487 15385 20499 15419
rect 21542 15416 21548 15428
rect 21503 15388 21548 15416
rect 20441 15379 20499 15385
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 23584 15416 23612 15444
rect 24762 15416 24768 15428
rect 23584 15388 23980 15416
rect 24723 15388 24768 15416
rect 23952 15360 23980 15388
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 25133 15419 25191 15425
rect 25133 15385 25145 15419
rect 25179 15416 25191 15419
rect 25792 15416 25820 15444
rect 25179 15388 25820 15416
rect 25179 15385 25191 15388
rect 25133 15379 25191 15385
rect 9674 15348 9680 15360
rect 8128 15320 9680 15348
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 12526 15348 12532 15360
rect 9815 15320 12532 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 12986 15308 12992 15360
rect 13044 15308 13050 15360
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13780 15320 14289 15348
rect 13780 15308 13786 15320
rect 14277 15317 14289 15320
rect 14323 15348 14335 15351
rect 15562 15348 15568 15360
rect 14323 15320 15568 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18874 15348 18880 15360
rect 18647 15320 18880 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 19889 15351 19947 15357
rect 19889 15348 19901 15351
rect 19576 15320 19901 15348
rect 19576 15308 19582 15320
rect 19889 15317 19901 15320
rect 19935 15317 19947 15351
rect 19889 15311 19947 15317
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 23566 15348 23572 15360
rect 20864 15320 23572 15348
rect 20864 15308 20870 15320
rect 23566 15308 23572 15320
rect 23624 15308 23630 15360
rect 23934 15308 23940 15360
rect 23992 15348 23998 15360
rect 25685 15351 25743 15357
rect 25685 15348 25697 15351
rect 23992 15320 25697 15348
rect 23992 15308 23998 15320
rect 25685 15317 25697 15320
rect 25731 15317 25743 15351
rect 25685 15311 25743 15317
rect 26050 15308 26056 15360
rect 26108 15348 26114 15360
rect 26712 15348 26740 15456
rect 27249 15453 27261 15456
rect 27295 15453 27307 15487
rect 27249 15447 27307 15453
rect 27982 15444 27988 15496
rect 28040 15484 28046 15496
rect 28276 15493 28304 15524
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 28040 15456 28089 15484
rect 28040 15444 28046 15456
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 26108 15320 26740 15348
rect 26108 15308 26114 15320
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5500 15116 6009 15144
rect 5500 15104 5506 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 5997 15107 6055 15113
rect 4062 15076 4068 15088
rect 4023 15048 4068 15076
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 5074 15076 5080 15088
rect 4540 15048 5080 15076
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 4540 15008 4568 15048
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 6012 15076 6040 15107
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 8297 15147 8355 15153
rect 6788 15116 6960 15144
rect 6788 15104 6794 15116
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 6012 15048 6837 15076
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 6825 15039 6883 15045
rect 1903 14980 4568 15008
rect 4617 15011 4675 15017
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 4617 14977 4629 15011
rect 4663 15008 4675 15011
rect 4706 15008 4712 15020
rect 4663 14980 4712 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 4873 15011 4931 15017
rect 4873 14977 4885 15011
rect 4919 15008 4931 15011
rect 5258 15008 5264 15020
rect 4919 14980 5264 15008
rect 4919 14977 4931 14980
rect 4873 14971 4931 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 6932 15017 6960 15116
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 9030 15144 9036 15156
rect 8343 15116 9036 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 9824 15116 10793 15144
rect 9824 15104 9830 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 11974 15104 11980 15156
rect 12032 15104 12038 15156
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12618 15144 12624 15156
rect 12216 15116 12624 15144
rect 12216 15104 12222 15116
rect 12618 15104 12624 15116
rect 12676 15144 12682 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12676 15116 13093 15144
rect 12676 15104 12682 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 15657 15147 15715 15153
rect 13081 15107 13139 15113
rect 13556 15116 14872 15144
rect 10962 15076 10968 15088
rect 10923 15048 10968 15076
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11992 15076 12020 15104
rect 12342 15076 12348 15088
rect 11992 15048 12348 15076
rect 12342 15036 12348 15048
rect 12400 15076 12406 15088
rect 13556 15076 13584 15116
rect 12400 15048 13584 15076
rect 12400 15036 12406 15048
rect 14090 15036 14096 15088
rect 14148 15076 14154 15088
rect 14737 15079 14795 15085
rect 14737 15076 14749 15079
rect 14148 15048 14749 15076
rect 14148 15036 14154 15048
rect 14737 15045 14749 15048
rect 14783 15045 14795 15079
rect 14844 15076 14872 15116
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 16114 15144 16120 15156
rect 15703 15116 16120 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 16114 15104 16120 15116
rect 16172 15144 16178 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 16172 15116 16221 15144
rect 16172 15104 16178 15116
rect 16209 15113 16221 15116
rect 16255 15113 16267 15147
rect 20070 15144 20076 15156
rect 16209 15107 16267 15113
rect 17236 15116 19380 15144
rect 20031 15116 20076 15144
rect 17236 15076 17264 15116
rect 18230 15076 18236 15088
rect 14844 15048 17264 15076
rect 17328 15048 18236 15076
rect 14737 15039 14795 15045
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5868 14980 6561 15008
rect 5868 14968 5874 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7098 15008 7104 15020
rect 6963 14980 7104 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 6748 14940 6776 14971
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 9585 15011 9643 15017
rect 8536 14980 8708 15008
rect 8536 14968 8542 14980
rect 8570 14940 8576 14952
rect 6748 14912 8576 14940
rect 1762 14832 1768 14884
rect 1820 14872 1826 14884
rect 1820 14844 4660 14872
rect 1820 14832 1826 14844
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 3326 14804 3332 14816
rect 2823 14776 3332 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 4632 14804 4660 14844
rect 6748 14804 6776 14912
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 8680 14940 8708 14980
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 11146 15008 11152 15020
rect 9631 14980 11152 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 11968 15011 12026 15017
rect 11968 14977 11980 15011
rect 12014 15008 12026 15011
rect 12526 15008 12532 15020
rect 12014 14980 12532 15008
rect 12014 14977 12026 14980
rect 11968 14971 12026 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13538 15008 13544 15020
rect 13044 14980 13544 15008
rect 13044 14968 13050 14980
rect 13538 14968 13544 14980
rect 13596 15008 13602 15020
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13596 14980 14013 15008
rect 13596 14968 13602 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 14918 15008 14924 15020
rect 14599 14980 14924 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 15381 14971 15439 14977
rect 11698 14940 11704 14952
rect 8680 14912 11560 14940
rect 11659 14912 11704 14940
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 9122 14872 9128 14884
rect 7147 14844 9128 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10192 14844 10824 14872
rect 10192 14832 10198 14844
rect 10594 14804 10600 14816
rect 4632 14776 6776 14804
rect 10555 14776 10600 14804
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 10796 14813 10824 14844
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14773 10839 14807
rect 11532 14804 11560 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13504 14912 13737 14940
rect 13504 14900 13510 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 13740 14872 13768 14903
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 15396 14940 15424 14971
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 17000 14980 17049 15008
rect 17000 14968 17006 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 16850 14940 16856 14952
rect 13872 14912 15424 14940
rect 16811 14912 16856 14940
rect 13872 14900 13878 14912
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 17052 14940 17080 14971
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 17328 15017 17356 15048
rect 18230 15036 18236 15048
rect 18288 15076 18294 15088
rect 19245 15079 19303 15085
rect 19245 15076 19257 15079
rect 18288 15048 18460 15076
rect 18288 15036 18294 15048
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 17184 14980 17325 15008
rect 17184 14968 17190 14980
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 18322 15008 18328 15020
rect 18283 14980 18328 15008
rect 17313 14971 17371 14977
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 18432 15017 18460 15048
rect 18616 15048 19257 15076
rect 18616 15017 18644 15048
rect 19245 15045 19257 15048
rect 19291 15045 19303 15079
rect 19352 15076 19380 15116
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 20438 15104 20444 15156
rect 20496 15144 20502 15156
rect 20622 15144 20628 15156
rect 20496 15116 20628 15144
rect 20496 15104 20502 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 21361 15147 21419 15153
rect 21361 15144 21373 15147
rect 20772 15116 21373 15144
rect 20772 15104 20778 15116
rect 21361 15113 21373 15116
rect 21407 15113 21419 15147
rect 21361 15107 21419 15113
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22428 15116 22661 15144
rect 22428 15104 22434 15116
rect 22649 15113 22661 15116
rect 22695 15113 22707 15147
rect 23658 15144 23664 15156
rect 22649 15107 22707 15113
rect 22848 15116 23664 15144
rect 22002 15076 22008 15088
rect 19352 15048 22008 15076
rect 19245 15039 19303 15045
rect 22002 15036 22008 15048
rect 22060 15036 22066 15088
rect 22848 15085 22876 15116
rect 23658 15104 23664 15116
rect 23716 15144 23722 15156
rect 23937 15147 23995 15153
rect 23937 15144 23949 15147
rect 23716 15116 23949 15144
rect 23716 15104 23722 15116
rect 23937 15113 23949 15116
rect 23983 15113 23995 15147
rect 25590 15144 25596 15156
rect 25551 15116 25596 15144
rect 23937 15107 23995 15113
rect 25590 15104 25596 15116
rect 25648 15104 25654 15156
rect 27338 15144 27344 15156
rect 27299 15116 27344 15144
rect 27338 15104 27344 15116
rect 27396 15104 27402 15156
rect 22833 15079 22891 15085
rect 22833 15045 22845 15079
rect 22879 15045 22891 15079
rect 22833 15039 22891 15045
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 24762 15076 24768 15088
rect 23532 15048 24768 15076
rect 23532 15036 23538 15048
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18601 14971 18659 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19518 15008 19524 15020
rect 19479 14980 19524 15008
rect 19518 14968 19524 14980
rect 19576 14968 19582 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 20128 14980 20177 15008
rect 20128 14968 20134 14980
rect 20165 14977 20177 14980
rect 20211 15008 20223 15011
rect 20346 15008 20352 15020
rect 20211 14980 20352 15008
rect 20211 14977 20223 14980
rect 20165 14971 20223 14977
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 20806 15008 20812 15020
rect 20767 14980 20812 15008
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 21266 15008 21272 15020
rect 21227 14980 21272 15008
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 21450 15008 21456 15020
rect 21411 14980 21456 15008
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22554 15008 22560 15020
rect 22515 14980 22560 15008
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 22738 14968 22744 15020
rect 22796 15008 22802 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 22796 14980 23305 15008
rect 22796 14968 22802 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23934 15008 23940 15020
rect 23895 14980 23940 15008
rect 23293 14971 23351 14977
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 24136 15017 24164 15048
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 25682 15076 25688 15088
rect 25643 15048 25688 15076
rect 25682 15036 25688 15048
rect 25740 15036 25746 15088
rect 25869 15079 25927 15085
rect 25869 15045 25881 15079
rect 25915 15076 25927 15079
rect 25958 15076 25964 15088
rect 25915 15048 25964 15076
rect 25915 15045 25927 15048
rect 25869 15039 25927 15045
rect 25958 15036 25964 15048
rect 26016 15036 26022 15088
rect 26970 15036 26976 15088
rect 27028 15076 27034 15088
rect 27028 15048 27384 15076
rect 27028 15036 27034 15048
rect 24121 15011 24179 15017
rect 24121 14977 24133 15011
rect 24167 14977 24179 15011
rect 24121 14971 24179 14977
rect 25593 15011 25651 15017
rect 25593 14977 25605 15011
rect 25639 15008 25651 15011
rect 26602 15008 26608 15020
rect 25639 14980 26608 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 26602 14968 26608 14980
rect 26660 14968 26666 15020
rect 27154 15008 27160 15020
rect 27115 14980 27160 15008
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 27356 15017 27384 15048
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 19242 14940 19248 14952
rect 17052 14912 18920 14940
rect 19203 14912 19248 14940
rect 14274 14872 14280 14884
rect 13740 14844 14280 14872
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 14366 14832 14372 14884
rect 14424 14872 14430 14884
rect 14642 14872 14648 14884
rect 14424 14844 14648 14872
rect 14424 14832 14430 14844
rect 14642 14832 14648 14844
rect 14700 14872 14706 14884
rect 17862 14872 17868 14884
rect 14700 14844 17868 14872
rect 14700 14832 14706 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 18506 14832 18512 14884
rect 18564 14872 18570 14884
rect 18782 14872 18788 14884
rect 18564 14844 18788 14872
rect 18564 14832 18570 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 18892 14872 18920 14912
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19392 14912 19441 14940
rect 19392 14900 19398 14912
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 19996 14912 20208 14940
rect 19996 14872 20024 14912
rect 18892 14844 20024 14872
rect 20180 14872 20208 14912
rect 20254 14900 20260 14952
rect 20312 14940 20318 14952
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 20312 14912 23397 14940
rect 20312 14900 20318 14912
rect 23385 14909 23397 14912
rect 23431 14909 23443 14943
rect 28350 14940 28356 14952
rect 28311 14912 28356 14940
rect 23385 14903 23443 14909
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 21082 14872 21088 14884
rect 20180 14844 21088 14872
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 22830 14872 22836 14884
rect 22791 14844 22836 14872
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 13722 14804 13728 14816
rect 11532 14776 13728 14804
rect 10781 14767 10839 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14608 14776 14841 14804
rect 14608 14764 14614 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15470 14804 15476 14816
rect 14976 14776 15476 14804
rect 14976 14764 14982 14776
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16758 14804 16764 14816
rect 15804 14776 16764 14804
rect 15804 14764 15810 14776
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 18138 14804 18144 14816
rect 18099 14776 18144 14804
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 20070 14804 20076 14816
rect 18288 14776 20076 14804
rect 18288 14764 18294 14776
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 20898 14804 20904 14816
rect 20763 14776 20904 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22186 14804 22192 14816
rect 22143 14776 22192 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22186 14764 22192 14776
rect 22244 14804 22250 14816
rect 22922 14804 22928 14816
rect 22244 14776 22928 14804
rect 22244 14764 22250 14776
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 24578 14804 24584 14816
rect 23440 14776 24584 14804
rect 23440 14764 23446 14776
rect 24578 14764 24584 14776
rect 24636 14764 24642 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 1912 14572 3188 14600
rect 1912 14560 1918 14572
rect 3160 14532 3188 14572
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3292 14572 3433 14600
rect 3292 14560 3298 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 11238 14600 11244 14612
rect 3421 14563 3479 14569
rect 4264 14572 11244 14600
rect 4264 14532 4292 14572
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 16942 14600 16948 14612
rect 12032 14572 16948 14600
rect 12032 14560 12038 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 18598 14600 18604 14612
rect 17828 14572 18604 14600
rect 17828 14560 17834 14572
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 21177 14603 21235 14609
rect 21177 14600 21189 14603
rect 18840 14572 21189 14600
rect 18840 14560 18846 14572
rect 21177 14569 21189 14572
rect 21223 14569 21235 14603
rect 23566 14600 23572 14612
rect 23479 14572 23572 14600
rect 21177 14563 21235 14569
rect 23566 14560 23572 14572
rect 23624 14600 23630 14612
rect 24302 14600 24308 14612
rect 23624 14572 24308 14600
rect 23624 14560 23630 14572
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 24578 14560 24584 14612
rect 24636 14600 24642 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 24636 14572 25237 14600
rect 24636 14560 24642 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 25225 14563 25283 14569
rect 3160 14504 4292 14532
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 5629 14535 5687 14541
rect 5629 14532 5641 14535
rect 5316 14504 5641 14532
rect 5316 14492 5322 14504
rect 5629 14501 5641 14504
rect 5675 14532 5687 14535
rect 5675 14504 9720 14532
rect 5675 14501 5687 14504
rect 5629 14495 5687 14501
rect 2038 14464 2044 14476
rect 1999 14436 2044 14464
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 7098 14464 7104 14476
rect 5500 14436 7104 14464
rect 5500 14424 5506 14436
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 9398 14464 9404 14476
rect 7156 14436 9404 14464
rect 7156 14424 7162 14436
rect 9398 14424 9404 14436
rect 9456 14464 9462 14476
rect 9456 14436 9536 14464
rect 9456 14424 9462 14436
rect 2314 14405 2320 14408
rect 2308 14359 2320 14405
rect 2372 14396 2378 14408
rect 4246 14396 4252 14408
rect 2372 14368 2408 14396
rect 4207 14368 4252 14396
rect 2314 14356 2320 14359
rect 2372 14356 2378 14368
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5408 14368 6101 14396
rect 5408 14356 5414 14368
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 8294 14396 8300 14408
rect 6420 14368 8300 14396
rect 6420 14356 6426 14368
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8536 14368 8585 14396
rect 8536 14356 8542 14368
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9508 14405 9536 14436
rect 9692 14405 9720 14504
rect 10870 14492 10876 14544
rect 10928 14532 10934 14544
rect 12894 14532 12900 14544
rect 10928 14504 12900 14532
rect 10928 14492 10934 14504
rect 12894 14492 12900 14504
rect 12952 14492 12958 14544
rect 15381 14535 15439 14541
rect 15381 14501 15393 14535
rect 15427 14532 15439 14535
rect 15746 14532 15752 14544
rect 15427 14504 15752 14532
rect 15427 14501 15439 14504
rect 15381 14495 15439 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 19058 14532 19064 14544
rect 18472 14504 19064 14532
rect 18472 14492 18478 14504
rect 19058 14492 19064 14504
rect 19116 14492 19122 14544
rect 20070 14492 20076 14544
rect 20128 14532 20134 14544
rect 21821 14535 21879 14541
rect 21821 14532 21833 14535
rect 20128 14504 21833 14532
rect 20128 14492 20134 14504
rect 21821 14501 21833 14504
rect 21867 14501 21879 14535
rect 21821 14495 21879 14501
rect 23109 14535 23167 14541
rect 23109 14501 23121 14535
rect 23155 14532 23167 14535
rect 23658 14532 23664 14544
rect 23155 14504 23664 14532
rect 23155 14501 23167 14504
rect 23109 14495 23167 14501
rect 23658 14492 23664 14504
rect 23716 14492 23722 14544
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 13596 14436 14504 14464
rect 13596 14424 13602 14436
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8996 14368 9321 14396
rect 8996 14356 9002 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12400 14368 13001 14396
rect 12400 14356 12406 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13136 14368 13185 14396
rect 13136 14356 13142 14368
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 14274 14396 14280 14408
rect 13320 14368 13365 14396
rect 14235 14368 14280 14396
rect 13320 14356 13326 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14476 14405 14504 14436
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 16908 14436 17448 14464
rect 16908 14424 16914 14436
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14792 14368 15117 14396
rect 14792 14356 14798 14368
rect 15105 14365 15117 14368
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15562 14396 15568 14408
rect 15427 14368 15568 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15804 14368 15945 14396
rect 15804 14356 15810 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 17420 14396 17448 14436
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 22462 14464 22468 14476
rect 18196 14436 22468 14464
rect 18196 14424 18202 14436
rect 22462 14424 22468 14436
rect 22520 14464 22526 14476
rect 25777 14467 25835 14473
rect 25777 14464 25789 14467
rect 22520 14436 22876 14464
rect 22520 14424 22526 14436
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17420 14368 18245 14396
rect 15933 14359 15991 14365
rect 4516 14331 4574 14337
rect 4516 14297 4528 14331
rect 4562 14328 4574 14331
rect 4890 14328 4896 14340
rect 4562 14300 4896 14328
rect 4562 14297 4574 14300
rect 4516 14291 4574 14297
rect 4890 14288 4896 14300
rect 4948 14288 4954 14340
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 8496 14328 8524 14356
rect 18156 14340 18184 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18414 14396 18420 14408
rect 18375 14368 18420 14396
rect 18233 14359 18291 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18598 14396 18604 14408
rect 18559 14368 18604 14396
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 18874 14356 18880 14408
rect 18932 14396 18938 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18932 14368 19625 14396
rect 18932 14356 18938 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19886 14396 19892 14408
rect 19847 14368 19892 14396
rect 19613 14359 19671 14365
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14396 20407 14399
rect 20714 14396 20720 14408
rect 20395 14368 20720 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 20714 14356 20720 14368
rect 20772 14396 20778 14408
rect 21082 14396 21088 14408
rect 20772 14368 20944 14396
rect 21043 14368 21088 14396
rect 20772 14356 20778 14368
rect 5132 14300 8524 14328
rect 9401 14331 9459 14337
rect 5132 14288 5138 14300
rect 9401 14297 9413 14331
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8389 14263 8447 14269
rect 8389 14229 8401 14263
rect 8435 14260 8447 14263
rect 8662 14260 8668 14272
rect 8435 14232 8668 14260
rect 8435 14229 8447 14232
rect 8389 14223 8447 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9122 14260 9128 14272
rect 9083 14232 9128 14260
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9416 14260 9444 14291
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 10597 14331 10655 14337
rect 10597 14328 10609 14331
rect 9640 14300 10609 14328
rect 9640 14288 9646 14300
rect 10597 14297 10609 14300
rect 10643 14297 10655 14331
rect 10597 14291 10655 14297
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 13722 14328 13728 14340
rect 12952 14300 13728 14328
rect 12952 14288 12958 14300
rect 13722 14288 13728 14300
rect 13780 14328 13786 14340
rect 14645 14331 14703 14337
rect 14645 14328 14657 14331
rect 13780 14300 14657 14328
rect 13780 14288 13786 14300
rect 14645 14297 14657 14300
rect 14691 14328 14703 14331
rect 16209 14331 16267 14337
rect 14691 14300 15332 14328
rect 14691 14297 14703 14300
rect 14645 14291 14703 14297
rect 10318 14260 10324 14272
rect 9416 14232 10324 14260
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10410 14220 10416 14272
rect 10468 14260 10474 14272
rect 11885 14263 11943 14269
rect 11885 14260 11897 14263
rect 10468 14232 11897 14260
rect 10468 14220 10474 14232
rect 11885 14229 11897 14232
rect 11931 14229 11943 14263
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 11885 14223 11943 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 15304 14260 15332 14300
rect 16209 14297 16221 14331
rect 16255 14328 16267 14331
rect 16482 14328 16488 14340
rect 16255 14300 16488 14328
rect 16255 14297 16267 14300
rect 16209 14291 16267 14297
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 18046 14328 18052 14340
rect 17434 14300 18052 14328
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 18138 14288 18144 14340
rect 18196 14288 18202 14340
rect 18322 14288 18328 14340
rect 18380 14328 18386 14340
rect 18509 14331 18567 14337
rect 18509 14328 18521 14331
rect 18380 14300 18521 14328
rect 18380 14288 18386 14300
rect 18509 14297 18521 14300
rect 18555 14297 18567 14331
rect 18509 14291 18567 14297
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 18748 14300 19809 14328
rect 18748 14288 18754 14300
rect 19797 14297 19809 14300
rect 19843 14297 19855 14331
rect 20438 14328 20444 14340
rect 19797 14291 19855 14297
rect 19904 14300 20444 14328
rect 17218 14260 17224 14272
rect 15304 14232 17224 14260
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 17681 14263 17739 14269
rect 17681 14229 17693 14263
rect 17727 14260 17739 14263
rect 18230 14260 18236 14272
rect 17727 14232 18236 14260
rect 17727 14229 17739 14232
rect 17681 14223 17739 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18782 14260 18788 14272
rect 18743 14232 18788 14260
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19904 14269 19932 14300
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 20625 14331 20683 14337
rect 20625 14297 20637 14331
rect 20671 14297 20683 14331
rect 20916 14328 20944 14368
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21542 14356 21548 14408
rect 21600 14396 21606 14408
rect 22848 14405 22876 14436
rect 23032 14436 25789 14464
rect 21729 14399 21787 14405
rect 21729 14396 21741 14399
rect 21600 14368 21741 14396
rect 21600 14356 21606 14368
rect 21729 14365 21741 14368
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 21560 14328 21588 14356
rect 20916 14300 21588 14328
rect 20625 14291 20683 14297
rect 19889 14263 19947 14269
rect 19889 14229 19901 14263
rect 19935 14229 19947 14263
rect 20346 14260 20352 14272
rect 20307 14232 20352 14260
rect 19889 14223 19947 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 20640 14260 20668 14291
rect 21634 14260 21640 14272
rect 20640 14232 21640 14260
rect 21634 14220 21640 14232
rect 21692 14260 21698 14272
rect 21928 14260 21956 14359
rect 22002 14288 22008 14340
rect 22060 14328 22066 14340
rect 23032 14328 23060 14436
rect 25777 14433 25789 14436
rect 25823 14433 25835 14467
rect 25777 14427 25835 14433
rect 24578 14396 24584 14408
rect 24539 14368 24584 14396
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 24946 14396 24952 14408
rect 24811 14368 24952 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 24946 14356 24952 14368
rect 25004 14356 25010 14408
rect 22060 14300 23060 14328
rect 23109 14331 23167 14337
rect 22060 14288 22066 14300
rect 23109 14297 23121 14331
rect 23155 14328 23167 14331
rect 24394 14328 24400 14340
rect 23155 14300 24400 14328
rect 23155 14297 23167 14300
rect 23109 14291 23167 14297
rect 24394 14288 24400 14300
rect 24452 14288 24458 14340
rect 22922 14260 22928 14272
rect 21692 14232 21956 14260
rect 22883 14232 22928 14260
rect 21692 14220 21698 14232
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24544 14232 24593 14260
rect 24544 14220 24550 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1820 14028 1869 14056
rect 1820 14016 1826 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 7282 14056 7288 14068
rect 5868 14028 7098 14056
rect 7243 14028 7288 14056
rect 5868 14016 5874 14028
rect 5534 13988 5540 14000
rect 4448 13960 5540 13988
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2222 13880 2228 13932
rect 2280 13920 2286 13932
rect 4448 13929 4476 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 2665 13923 2723 13929
rect 2665 13920 2677 13923
rect 2280 13892 2677 13920
rect 2280 13880 2286 13892
rect 2665 13889 2677 13892
rect 2711 13889 2723 13923
rect 2665 13883 2723 13889
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13889 4491 13923
rect 4689 13923 4747 13929
rect 4689 13920 4701 13923
rect 4433 13883 4491 13889
rect 4540 13892 4701 13920
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 2424 13784 2452 13815
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 4540 13852 4568 13892
rect 4689 13889 4701 13892
rect 4735 13889 4747 13923
rect 4689 13883 4747 13889
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7070 13929 7098 14028
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10686 14056 10692 14068
rect 10459 14028 10692 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 12434 14056 12440 14068
rect 11103 14028 12440 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 13078 14056 13084 14068
rect 13039 14028 13084 14056
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14642 14056 14648 14068
rect 13412 14028 14228 14056
rect 14603 14028 14648 14056
rect 13412 14016 13418 14028
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 11238 13988 11244 14000
rect 9631 13960 11244 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11968 13991 12026 13997
rect 11968 13957 11980 13991
rect 12014 13988 12026 13991
rect 12802 13988 12808 14000
rect 12014 13960 12808 13988
rect 12014 13957 12026 13960
rect 11968 13951 12026 13957
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 13909 13991 13967 13997
rect 13909 13957 13921 13991
rect 13955 13988 13967 13991
rect 13998 13988 14004 14000
rect 13955 13960 14004 13988
rect 13955 13957 13967 13960
rect 13909 13951 13967 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6512 13892 6653 13920
rect 6512 13880 6518 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6734 13923 6792 13929
rect 6734 13889 6746 13923
rect 6780 13889 6792 13923
rect 6734 13883 6792 13889
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 7017 13923 7098 13929
rect 7017 13889 7029 13923
rect 7063 13892 7098 13923
rect 7147 13923 7205 13929
rect 7063 13889 7075 13892
rect 7017 13883 7075 13889
rect 7147 13889 7159 13923
rect 7193 13920 7205 13923
rect 7282 13920 7288 13932
rect 7193 13892 7288 13920
rect 7193 13889 7205 13892
rect 7147 13883 7205 13889
rect 3476 13824 4568 13852
rect 3476 13812 3482 13824
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6749 13852 6777 13883
rect 6236 13824 6777 13852
rect 6236 13812 6242 13824
rect 3786 13784 3792 13796
rect 1912 13756 2452 13784
rect 3747 13756 3792 13784
rect 1912 13744 1918 13756
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 6932 13784 6960 13883
rect 7282 13880 7288 13892
rect 7340 13920 7346 13932
rect 7742 13920 7748 13932
rect 7340 13892 7748 13920
rect 7340 13880 7346 13892
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 10226 13920 10232 13932
rect 8352 13892 10232 13920
rect 8352 13880 8358 13892
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 10686 13920 10692 13932
rect 10551 13892 10692 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10928 13892 10977 13920
rect 10928 13880 10934 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 11146 13920 11152 13932
rect 11107 13892 11152 13920
rect 10965 13883 11023 13889
rect 11146 13880 11152 13892
rect 11204 13920 11210 13932
rect 11204 13892 13676 13920
rect 11204 13880 11210 13892
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8938 13852 8944 13864
rect 8536 13824 8944 13852
rect 8536 13812 8542 13824
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 10778 13852 10784 13864
rect 8996 13824 10784 13852
rect 8996 13812 9002 13824
rect 10778 13812 10784 13824
rect 10836 13852 10842 13864
rect 11698 13852 11704 13864
rect 10836 13824 11560 13852
rect 11659 13824 11704 13852
rect 10836 13812 10842 13824
rect 9030 13784 9036 13796
rect 6512 13756 9036 13784
rect 6512 13744 6518 13756
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 5810 13716 5816 13728
rect 3108 13688 5816 13716
rect 3108 13676 3114 13688
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 8297 13719 8355 13725
rect 8297 13685 8309 13719
rect 8343 13716 8355 13719
rect 8570 13716 8576 13728
rect 8343 13688 8576 13716
rect 8343 13685 8355 13688
rect 8297 13679 8355 13685
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 11532 13716 11560 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 13648 13852 13676 13892
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14200 13920 14228 14028
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 15930 14056 15936 14068
rect 15712 14028 15936 14056
rect 15712 14016 15718 14028
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16942 14056 16948 14068
rect 16903 14028 16948 14056
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 19981 14059 20039 14065
rect 17276 14028 19748 14056
rect 17276 14016 17282 14028
rect 16226 13991 16284 13997
rect 16226 13957 16238 13991
rect 16272 13988 16284 13991
rect 17126 13988 17132 14000
rect 16272 13960 17132 13988
rect 16272 13957 16284 13960
rect 16226 13951 16284 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 17678 13988 17684 14000
rect 17639 13960 17684 13988
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 19613 13991 19671 13997
rect 19613 13988 19625 13991
rect 18708 13960 19625 13988
rect 18708 13932 18736 13960
rect 19613 13957 19625 13960
rect 19659 13957 19671 13991
rect 19720 13988 19748 14028
rect 19981 14025 19993 14059
rect 20027 14056 20039 14059
rect 20714 14056 20720 14068
rect 20027 14028 20720 14056
rect 20027 14025 20039 14028
rect 19981 14019 20039 14025
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 22066 14028 23428 14056
rect 20530 13988 20536 14000
rect 19720 13960 20536 13988
rect 19613 13951 19671 13957
rect 20530 13948 20536 13960
rect 20588 13948 20594 14000
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 22066 13988 22094 14028
rect 23400 13988 23428 14028
rect 25685 13991 25743 13997
rect 25685 13988 25697 13991
rect 20680 13960 22094 13988
rect 22480 13960 23336 13988
rect 23400 13960 25697 13988
rect 20680 13948 20686 13960
rect 22480 13932 22508 13960
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 13780 13892 13825 13920
rect 14200 13892 14565 13920
rect 13780 13880 13786 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 14090 13852 14096 13864
rect 13648 13824 14096 13852
rect 14090 13812 14096 13824
rect 14148 13852 14154 13864
rect 14568 13852 14596 13883
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 14700 13892 14745 13920
rect 14700 13880 14706 13892
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15344 13892 15669 13920
rect 15344 13880 15350 13892
rect 15657 13889 15669 13892
rect 15703 13889 15715 13923
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15657 13883 15715 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 15948 13852 15976 13883
rect 16022 13880 16028 13932
rect 16080 13929 16086 13932
rect 16080 13920 16088 13929
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16080 13892 16125 13920
rect 16211 13892 16865 13920
rect 16080 13883 16088 13892
rect 16080 13880 16086 13883
rect 14148 13824 14504 13852
rect 14568 13824 14688 13852
rect 15948 13824 16068 13852
rect 14148 13812 14154 13824
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13906 13784 13912 13796
rect 12860 13756 13912 13784
rect 12860 13744 12866 13756
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 11974 13716 11980 13728
rect 11532 13688 11980 13716
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 13541 13719 13599 13725
rect 13541 13685 13553 13719
rect 13587 13716 13599 13719
rect 14182 13716 14188 13728
rect 13587 13688 14188 13716
rect 13587 13685 13599 13688
rect 13541 13679 13599 13685
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 14476 13716 14504 13824
rect 14660 13784 14688 13824
rect 15930 13784 15936 13796
rect 14660 13756 15936 13784
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 16040 13784 16068 13824
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 16211 13852 16239 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17310 13920 17316 13932
rect 17083 13892 17316 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13889 17923 13923
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 17865 13883 17923 13889
rect 16172 13824 16239 13852
rect 16172 13812 16178 13824
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 17880 13852 17908 13883
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18874 13880 18880 13892
rect 18932 13920 18938 13932
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 18932 13892 19533 13920
rect 18932 13880 18938 13892
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 19886 13920 19892 13932
rect 19843 13892 19892 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 19886 13880 19892 13892
rect 19944 13920 19950 13932
rect 22462 13920 22468 13932
rect 19944 13892 22094 13920
rect 22423 13892 22468 13920
rect 19944 13880 19950 13892
rect 16356 13824 17908 13852
rect 19061 13855 19119 13861
rect 16356 13812 16362 13824
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19702 13852 19708 13864
rect 19107 13824 19708 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 20533 13855 20591 13861
rect 20533 13821 20545 13855
rect 20579 13852 20591 13855
rect 20714 13852 20720 13864
rect 20579 13824 20720 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 22066 13852 22094 13892
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22922 13920 22928 13932
rect 22756 13892 22928 13920
rect 22756 13852 22784 13892
rect 22922 13880 22928 13892
rect 22980 13920 22986 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 22980 13892 23213 13920
rect 22980 13880 22986 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23308 13861 23336 13960
rect 25685 13957 25697 13960
rect 25731 13957 25743 13991
rect 25685 13951 25743 13957
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13920 24271 13923
rect 24578 13920 24584 13932
rect 24259 13892 24584 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 22066 13824 22784 13852
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 16942 13784 16948 13796
rect 16040 13756 16948 13784
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 18049 13787 18107 13793
rect 18049 13784 18061 13787
rect 17276 13756 18061 13784
rect 17276 13744 17282 13756
rect 18049 13753 18061 13756
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 20346 13744 20352 13796
rect 20404 13784 20410 13796
rect 20809 13787 20867 13793
rect 20809 13784 20821 13787
rect 20404 13756 20821 13784
rect 20404 13744 20410 13756
rect 20809 13753 20821 13756
rect 20855 13753 20867 13787
rect 20809 13747 20867 13753
rect 23569 13787 23627 13793
rect 23569 13753 23581 13787
rect 23615 13784 23627 13787
rect 24228 13784 24256 13883
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 25038 13920 25044 13932
rect 24999 13892 25044 13920
rect 25038 13880 25044 13892
rect 25096 13880 25102 13932
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13920 25283 13923
rect 25590 13920 25596 13932
rect 25271 13892 25596 13920
rect 25271 13889 25283 13892
rect 25225 13883 25283 13889
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13852 24363 13855
rect 25240 13852 25268 13883
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 24351 13824 24532 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 23615 13756 24256 13784
rect 23615 13753 23627 13756
rect 23569 13747 23627 13753
rect 14642 13716 14648 13728
rect 14476 13688 14648 13716
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 20162 13716 20168 13728
rect 15528 13688 20168 13716
rect 15528 13676 15534 13688
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 20993 13719 21051 13725
rect 20993 13685 21005 13719
rect 21039 13716 21051 13719
rect 21450 13716 21456 13728
rect 21039 13688 21456 13716
rect 21039 13685 21051 13688
rect 20993 13679 21051 13685
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 22373 13719 22431 13725
rect 22373 13685 22385 13719
rect 22419 13716 22431 13719
rect 23106 13716 23112 13728
rect 22419 13688 23112 13716
rect 22419 13685 22431 13688
rect 22373 13679 22431 13685
rect 23106 13676 23112 13688
rect 23164 13676 23170 13728
rect 24504 13716 24532 13824
rect 24596 13824 25268 13852
rect 24596 13793 24624 13824
rect 24581 13787 24639 13793
rect 24581 13753 24593 13787
rect 24627 13753 24639 13787
rect 24581 13747 24639 13753
rect 24946 13716 24952 13728
rect 24504 13688 24952 13716
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 25130 13716 25136 13728
rect 25091 13688 25136 13716
rect 25130 13676 25136 13688
rect 25188 13676 25194 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3421 13515 3479 13521
rect 3421 13512 3433 13515
rect 2832 13484 3433 13512
rect 2832 13472 2838 13484
rect 3421 13481 3433 13484
rect 3467 13512 3479 13515
rect 3970 13512 3976 13524
rect 3467 13484 3976 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 6546 13472 6552 13524
rect 6604 13512 6610 13524
rect 7929 13515 7987 13521
rect 7929 13512 7941 13515
rect 6604 13484 7941 13512
rect 6604 13472 6610 13484
rect 7929 13481 7941 13484
rect 7975 13481 7987 13515
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 7929 13475 7987 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12584 13484 12633 13512
rect 12584 13472 12590 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 13633 13515 13691 13521
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 13814 13512 13820 13524
rect 13679 13484 13820 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14516 13484 14565 13512
rect 14516 13472 14522 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 16196 13515 16254 13521
rect 16196 13481 16208 13515
rect 16242 13512 16254 13515
rect 16574 13512 16580 13524
rect 16242 13484 16580 13512
rect 16242 13481 16254 13484
rect 16196 13475 16254 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 20898 13512 20904 13524
rect 19843 13484 20904 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21039 13484 24348 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 14734 13444 14740 13456
rect 8527 13416 14740 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 14734 13404 14740 13416
rect 14792 13404 14798 13456
rect 18785 13447 18843 13453
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 19610 13444 19616 13456
rect 18831 13416 19616 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 19610 13404 19616 13416
rect 19668 13444 19674 13456
rect 19978 13444 19984 13456
rect 19668 13416 19984 13444
rect 19668 13404 19674 13416
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 20438 13404 20444 13456
rect 20496 13444 20502 13456
rect 21729 13447 21787 13453
rect 20496 13416 21496 13444
rect 20496 13404 20502 13416
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9088 13348 9352 13376
rect 9088 13336 9094 13348
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1912 13280 2053 13308
rect 1912 13268 1918 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4522 13308 4528 13320
rect 4019 13280 4528 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 4856 13280 6561 13308
rect 4856 13268 4862 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6816 13311 6874 13317
rect 6816 13277 6828 13311
rect 6862 13308 6874 13311
rect 7190 13308 7196 13320
rect 6862 13280 7196 13308
rect 6862 13277 6874 13280
rect 6816 13271 6874 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 9122 13308 9128 13320
rect 9083 13280 9128 13308
rect 8389 13271 8447 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9218 13311 9276 13317
rect 9218 13277 9230 13311
rect 9264 13277 9276 13311
rect 9218 13271 9276 13277
rect 2130 13200 2136 13252
rect 2188 13240 2194 13252
rect 2286 13243 2344 13249
rect 2286 13240 2298 13243
rect 2188 13212 2298 13240
rect 2188 13200 2194 13212
rect 2286 13209 2298 13212
rect 2332 13209 2344 13243
rect 2286 13203 2344 13209
rect 4976 13243 5034 13249
rect 4976 13209 4988 13243
rect 5022 13240 5034 13243
rect 5810 13240 5816 13252
rect 5022 13212 5816 13240
rect 5022 13209 5034 13212
rect 4976 13203 5034 13209
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 6270 13200 6276 13252
rect 6328 13240 6334 13252
rect 9232 13240 9260 13271
rect 6328 13212 9260 13240
rect 9324 13240 9352 13348
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 16574 13376 16580 13388
rect 13556 13348 16580 13376
rect 9416 13308 9444 13336
rect 9590 13311 9648 13317
rect 9590 13308 9602 13311
rect 9416 13280 9602 13308
rect 9590 13277 9602 13280
rect 9636 13277 9648 13311
rect 10410 13308 10416 13320
rect 10371 13280 10416 13308
rect 9590 13271 9648 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 11020 13280 12817 13308
rect 11020 13268 11026 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13262 13308 13268 13320
rect 13127 13280 13268 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13556 13317 13584 13348
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 19702 13376 19708 13388
rect 19663 13348 19708 13376
rect 19702 13336 19708 13348
rect 19760 13336 19766 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20772 13348 20852 13376
rect 20772 13336 20778 13348
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 13541 13271 13599 13277
rect 13648 13280 14381 13308
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9324 13212 9413 13240
rect 6328 13200 6334 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13209 9551 13243
rect 9493 13203 9551 13209
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4157 13175 4215 13181
rect 4157 13172 4169 13175
rect 3752 13144 4169 13172
rect 3752 13132 3758 13144
rect 4157 13141 4169 13144
rect 4203 13172 4215 13175
rect 5350 13172 5356 13184
rect 4203 13144 5356 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 6089 13175 6147 13181
rect 6089 13172 6101 13175
rect 5960 13144 6101 13172
rect 5960 13132 5966 13144
rect 6089 13141 6101 13144
rect 6135 13172 6147 13175
rect 9508 13172 9536 13203
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 10980 13240 11008 13268
rect 10284 13212 11008 13240
rect 10284 13200 10290 13212
rect 12158 13200 12164 13252
rect 12216 13240 12222 13252
rect 13648 13240 13676 13280
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 14645 13311 14703 13317
rect 14645 13308 14657 13311
rect 14516 13280 14657 13308
rect 14516 13268 14522 13280
rect 14645 13277 14657 13280
rect 14691 13308 14703 13311
rect 14691 13280 15700 13308
rect 14691 13277 14703 13280
rect 14645 13271 14703 13277
rect 12216 13212 13676 13240
rect 12216 13200 12222 13212
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 14274 13240 14280 13252
rect 13964 13212 14280 13240
rect 13964 13200 13970 13212
rect 14274 13200 14280 13212
rect 14332 13240 14338 13252
rect 15105 13243 15163 13249
rect 15105 13240 15117 13243
rect 14332 13212 15117 13240
rect 14332 13200 14338 13212
rect 15105 13209 15117 13212
rect 15151 13209 15163 13243
rect 15105 13203 15163 13209
rect 15289 13243 15347 13249
rect 15289 13209 15301 13243
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 6135 13144 9536 13172
rect 9769 13175 9827 13181
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 9769 13141 9781 13175
rect 9815 13172 9827 13175
rect 11882 13172 11888 13184
rect 9815 13144 11888 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12676 13144 13001 13172
rect 12676 13132 12682 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 12989 13135 13047 13141
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 15304 13172 15332 13203
rect 15470 13172 15476 13184
rect 13136 13144 15332 13172
rect 15431 13144 15476 13172
rect 13136 13132 13142 13144
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 15672 13172 15700 13280
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15804 13280 15945 13308
rect 15804 13268 15810 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 18230 13268 18236 13320
rect 18288 13308 18294 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 18288 13280 18613 13308
rect 18288 13268 18294 13280
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 20254 13308 20260 13320
rect 19475 13280 20260 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 17957 13243 18015 13249
rect 16356 13212 16698 13240
rect 16356 13200 16362 13212
rect 17957 13209 17969 13243
rect 18003 13240 18015 13243
rect 19444 13240 19472 13271
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20824 13317 20852 13348
rect 21468 13317 21496 13416
rect 21729 13413 21741 13447
rect 21775 13413 21787 13447
rect 24320 13444 24348 13484
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24452 13484 24593 13512
rect 24452 13472 24458 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 25038 13444 25044 13456
rect 24320 13416 25044 13444
rect 21729 13407 21787 13413
rect 21744 13376 21772 13407
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 24949 13379 25007 13385
rect 21744 13348 21956 13376
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13308 20591 13311
rect 20809 13311 20867 13317
rect 20579 13280 20760 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 18003 13212 19472 13240
rect 18003 13209 18015 13212
rect 17957 13203 18015 13209
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 20404 13212 20637 13240
rect 20404 13200 20410 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 19426 13172 19432 13184
rect 15672 13144 19432 13172
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 19978 13172 19984 13184
rect 19939 13144 19984 13172
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20732 13172 20760 13280
rect 20809 13277 20821 13311
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 20824 13240 20852 13271
rect 21542 13268 21548 13320
rect 21600 13308 21606 13320
rect 21600 13280 21645 13308
rect 21600 13268 21606 13280
rect 21726 13268 21732 13320
rect 21784 13308 21790 13320
rect 21784 13280 21829 13308
rect 21784 13268 21790 13280
rect 21928 13240 21956 13348
rect 24949 13345 24961 13379
rect 24995 13376 25007 13379
rect 25866 13376 25872 13388
rect 24995 13348 25872 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25866 13336 25872 13348
rect 25924 13336 25930 13388
rect 22554 13308 22560 13320
rect 22515 13280 22560 13308
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 23106 13268 23112 13320
rect 23164 13308 23170 13320
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 23164 13280 24777 13308
rect 23164 13268 23170 13280
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 25314 13308 25320 13320
rect 25087 13280 25320 13308
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 20824 13212 21956 13240
rect 22824 13243 22882 13249
rect 22824 13209 22836 13243
rect 22870 13240 22882 13243
rect 23198 13240 23204 13252
rect 22870 13212 23204 13240
rect 22870 13209 22882 13212
rect 22824 13203 22882 13209
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 24872 13240 24900 13271
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 25590 13308 25596 13320
rect 25551 13280 25596 13308
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 25958 13308 25964 13320
rect 25919 13280 25964 13308
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 23952 13212 24900 13240
rect 20806 13172 20812 13184
rect 20732 13144 20812 13172
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 23952 13181 23980 13212
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 21600 13144 23949 13172
rect 21600 13132 21606 13144
rect 23937 13141 23949 13144
rect 23983 13141 23995 13175
rect 24872 13172 24900 13212
rect 25130 13200 25136 13252
rect 25188 13240 25194 13252
rect 25777 13243 25835 13249
rect 25777 13240 25789 13243
rect 25188 13212 25789 13240
rect 25188 13200 25194 13212
rect 25777 13209 25789 13212
rect 25823 13209 25835 13243
rect 26421 13243 26479 13249
rect 26421 13240 26433 13243
rect 25777 13203 25835 13209
rect 25884 13212 26433 13240
rect 25682 13172 25688 13184
rect 24872 13144 25688 13172
rect 23937 13135 23995 13141
rect 25682 13132 25688 13144
rect 25740 13172 25746 13184
rect 25884 13172 25912 13212
rect 26421 13209 26433 13212
rect 26467 13209 26479 13243
rect 26421 13203 26479 13209
rect 25740 13144 25912 13172
rect 25740 13132 25746 13144
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12937 1915 12971
rect 1857 12931 1915 12937
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 4246 12968 4252 12980
rect 3099 12940 4252 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12869 1731 12903
rect 1872 12900 1900 12931
rect 4246 12928 4252 12940
rect 4304 12968 4310 12980
rect 4706 12968 4712 12980
rect 4304 12940 4712 12968
rect 4304 12928 4310 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 7374 12968 7380 12980
rect 5460 12940 7380 12968
rect 4341 12903 4399 12909
rect 1872 12872 4292 12900
rect 1673 12863 1731 12869
rect 1688 12696 1716 12863
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 4154 12832 4160 12844
rect 2179 12804 4160 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4264 12832 4292 12872
rect 4341 12869 4353 12903
rect 4387 12900 4399 12903
rect 5460 12900 5488 12940
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8297 12971 8355 12977
rect 8297 12937 8309 12971
rect 8343 12968 8355 12971
rect 9306 12968 9312 12980
rect 8343 12940 9312 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10410 12968 10416 12980
rect 9600 12940 10416 12968
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 4387 12872 5488 12900
rect 5644 12872 5825 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 4706 12832 4712 12844
rect 4264 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5074 12832 5080 12844
rect 4856 12804 5080 12832
rect 4856 12792 4862 12804
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 5644 12832 5672 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 5997 12903 6055 12909
rect 5997 12869 6009 12903
rect 6043 12869 6055 12903
rect 5997 12863 6055 12869
rect 5500 12804 5672 12832
rect 5500 12792 5506 12804
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6012 12832 6040 12863
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 9600 12909 9628 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 12250 12968 12256 12980
rect 12211 12940 12256 12968
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 19426 12968 19432 12980
rect 15948 12940 17080 12968
rect 19339 12940 19432 12968
rect 7101 12903 7159 12909
rect 7101 12900 7113 12903
rect 6512 12872 7113 12900
rect 6512 12860 6518 12872
rect 7101 12869 7113 12872
rect 7147 12869 7159 12903
rect 7101 12863 7159 12869
rect 9585 12903 9643 12909
rect 9585 12869 9597 12903
rect 9631 12869 9643 12903
rect 11698 12900 11704 12912
rect 9585 12863 9643 12869
rect 10152 12872 10548 12900
rect 6086 12832 6092 12844
rect 5776 12804 6092 12832
rect 5776 12792 5782 12804
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 6871 12835 6929 12841
rect 6871 12832 6883 12835
rect 6564 12804 6883 12832
rect 5626 12696 5632 12708
rect 1688 12668 5212 12696
rect 5587 12668 5632 12696
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 4430 12628 4436 12640
rect 1903 12600 4436 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5074 12628 5080 12640
rect 5031 12600 5080 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5184 12628 5212 12668
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 5718 12628 5724 12640
rect 5184 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 5994 12628 6000 12640
rect 5859 12600 6000 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6564 12628 6592 12804
rect 6871 12801 6883 12804
rect 6917 12801 6929 12835
rect 7006 12832 7012 12844
rect 6967 12804 7012 12832
rect 6871 12795 6929 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 7558 12832 7564 12844
rect 7423 12804 7564 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 10152 12832 10180 12872
rect 8720 12804 10180 12832
rect 8720 12792 8726 12804
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10410 12832 10416 12844
rect 10284 12804 10329 12832
rect 10371 12804 10416 12832
rect 10284 12792 10290 12804
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10520 12841 10548 12872
rect 10980 12872 11704 12900
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10686 12832 10692 12844
rect 10551 12804 10692 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10980 12841 11008 12872
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 12989 12903 13047 12909
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 13170 12900 13176 12912
rect 13035 12872 13176 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 15562 12900 15568 12912
rect 15212 12872 15568 12900
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 10965 12795 11023 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12529 12835 12587 12841
rect 12299 12804 12333 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 13998 12832 14004 12844
rect 12575 12804 14004 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 12268 12764 12296 12795
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 15212 12841 15240 12872
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 14148 12804 15209 12832
rect 14148 12792 14154 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15948 12841 15976 12940
rect 16298 12900 16304 12912
rect 16259 12872 16304 12900
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15344 12804 15945 12832
rect 15344 12792 15350 12804
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16163 12804 16957 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 17052 12832 17080 12940
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20714 12968 20720 12980
rect 20027 12940 20720 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 23198 12968 23204 12980
rect 23159 12940 23204 12968
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 25314 12968 25320 12980
rect 23308 12940 25320 12968
rect 18046 12900 18052 12912
rect 18007 12872 18052 12900
rect 18046 12860 18052 12872
rect 18104 12860 18110 12912
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 19444 12900 19472 12928
rect 22370 12900 22376 12912
rect 18196 12872 18644 12900
rect 19444 12872 22376 12900
rect 18196 12860 18202 12872
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 17052 12804 17141 12832
rect 16945 12795 17003 12801
rect 17129 12801 17141 12804
rect 17175 12832 17187 12835
rect 17678 12832 17684 12844
rect 17175 12804 17684 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 7708 12736 12434 12764
rect 7708 12724 7714 12736
rect 6733 12699 6791 12705
rect 6733 12665 6745 12699
rect 6779 12696 6791 12699
rect 7466 12696 7472 12708
rect 6779 12668 7472 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 6822 12628 6828 12640
rect 6564 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12628 6886 12640
rect 8478 12628 8484 12640
rect 6880 12600 8484 12628
rect 6880 12588 6886 12600
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9088 12600 10057 12628
rect 9088 12588 9094 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 12406 12628 12434 12736
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 15470 12764 15476 12776
rect 12676 12736 15476 12764
rect 12676 12724 12682 12736
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 14550 12656 14556 12708
rect 14608 12696 14614 12708
rect 16132 12696 16160 12795
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16816 12736 16865 12764
rect 16816 12724 16822 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16960 12764 16988 12795
rect 17678 12792 17684 12804
rect 17736 12792 17742 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 17880 12764 17908 12795
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 18288 12804 18521 12832
rect 18288 12792 18294 12804
rect 18509 12801 18521 12804
rect 18555 12801 18567 12835
rect 18616 12832 18644 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 19242 12841 19248 12844
rect 19233 12835 19248 12841
rect 19233 12832 19245 12835
rect 18616 12804 19245 12832
rect 18509 12795 18567 12801
rect 19233 12801 19245 12804
rect 19300 12832 19306 12844
rect 20530 12832 20536 12844
rect 19300 12804 20536 12832
rect 19233 12795 19248 12801
rect 19242 12792 19248 12795
rect 19300 12792 19306 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21094 12835 21152 12841
rect 21094 12832 21106 12835
rect 20772 12804 21106 12832
rect 20772 12792 20778 12804
rect 21094 12801 21106 12804
rect 21140 12801 21152 12835
rect 21094 12795 21152 12801
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 21450 12832 21456 12844
rect 21324 12804 21456 12832
rect 21324 12792 21330 12804
rect 21450 12792 21456 12804
rect 21508 12832 21514 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21508 12804 22017 12832
rect 21508 12792 21514 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22554 12832 22560 12844
rect 22005 12795 22063 12801
rect 22204 12804 22560 12832
rect 17954 12764 17960 12776
rect 16960 12736 17960 12764
rect 16853 12727 16911 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 22204 12764 22232 12804
rect 22554 12792 22560 12804
rect 22612 12832 22618 12844
rect 22738 12832 22744 12844
rect 22612 12804 22744 12832
rect 22612 12792 22618 12804
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 21407 12736 22232 12764
rect 22281 12767 22339 12773
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 22281 12733 22293 12767
rect 22327 12764 22339 12767
rect 23308 12764 23336 12940
rect 25314 12928 25320 12940
rect 25372 12968 25378 12980
rect 26050 12968 26056 12980
rect 25372 12940 26056 12968
rect 25372 12928 25378 12940
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 25958 12900 25964 12912
rect 23400 12872 25964 12900
rect 23400 12841 23428 12872
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 23385 12835 23443 12841
rect 23385 12801 23397 12835
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 23477 12835 23535 12841
rect 23477 12801 23489 12835
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12801 23627 12835
rect 23569 12795 23627 12801
rect 23492 12764 23520 12795
rect 22327 12736 23520 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 22572 12708 22600 12736
rect 16666 12696 16672 12708
rect 14608 12668 16160 12696
rect 16500 12668 16672 12696
rect 14608 12656 14614 12668
rect 12802 12628 12808 12640
rect 12406 12600 12808 12628
rect 10045 12591 10103 12597
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 14461 12631 14519 12637
rect 14461 12597 14473 12631
rect 14507 12628 14519 12631
rect 16500 12628 16528 12668
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 22189 12699 22247 12705
rect 22189 12696 22201 12699
rect 21508 12668 22201 12696
rect 21508 12656 21514 12668
rect 22189 12665 22201 12668
rect 22235 12665 22247 12699
rect 22189 12659 22247 12665
rect 22554 12656 22560 12708
rect 22612 12656 22618 12708
rect 23584 12696 23612 12795
rect 23658 12792 23664 12844
rect 23716 12841 23722 12844
rect 23716 12835 23745 12841
rect 23733 12801 23745 12835
rect 24486 12832 24492 12844
rect 24447 12804 24492 12832
rect 23716 12795 23745 12801
rect 23716 12792 23722 12795
rect 24486 12792 24492 12804
rect 24544 12832 24550 12844
rect 24762 12832 24768 12844
rect 24544 12804 24768 12832
rect 24544 12792 24550 12804
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12832 25559 12835
rect 25774 12832 25780 12844
rect 25547 12804 25780 12832
rect 25547 12801 25559 12804
rect 25501 12795 25559 12801
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 23842 12764 23848 12776
rect 23803 12736 23848 12764
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 24394 12764 24400 12776
rect 24355 12736 24400 12764
rect 24394 12724 24400 12736
rect 24452 12724 24458 12776
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24673 12767 24731 12773
rect 24673 12733 24685 12767
rect 24719 12764 24731 12767
rect 25590 12764 25596 12776
rect 24719 12736 25596 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 24596 12696 24624 12727
rect 25590 12724 25596 12736
rect 25648 12724 25654 12776
rect 25682 12724 25688 12776
rect 25740 12764 25746 12776
rect 26145 12767 26203 12773
rect 26145 12764 26157 12767
rect 25740 12736 26157 12764
rect 25740 12724 25746 12736
rect 26145 12733 26157 12736
rect 26191 12733 26203 12767
rect 26145 12727 26203 12733
rect 25222 12696 25228 12708
rect 23584 12668 25228 12696
rect 25222 12656 25228 12668
rect 25280 12696 25286 12708
rect 25958 12696 25964 12708
rect 25280 12668 25964 12696
rect 25280 12656 25286 12668
rect 25958 12656 25964 12668
rect 26016 12656 26022 12708
rect 14507 12600 16528 12628
rect 14507 12597 14519 12600
rect 14461 12591 14519 12597
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 18046 12628 18052 12640
rect 16632 12600 18052 12628
rect 16632 12588 16638 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18690 12628 18696 12640
rect 18651 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12628 18754 12640
rect 19334 12628 19340 12640
rect 18748 12600 19340 12628
rect 18748 12588 18754 12600
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 20990 12588 20996 12640
rect 21048 12628 21054 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21048 12600 22109 12628
rect 21048 12588 21054 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22097 12591 22155 12597
rect 24857 12631 24915 12637
rect 24857 12597 24869 12631
rect 24903 12628 24915 12631
rect 24946 12628 24952 12640
rect 24903 12600 24952 12628
rect 24903 12597 24915 12600
rect 24857 12591 24915 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25317 12631 25375 12637
rect 25317 12628 25329 12631
rect 25096 12600 25329 12628
rect 25096 12588 25102 12600
rect 25317 12597 25329 12600
rect 25363 12597 25375 12631
rect 25317 12591 25375 12597
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2406 12424 2412 12436
rect 2087 12396 2412 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2406 12384 2412 12396
rect 2464 12424 2470 12436
rect 6638 12424 6644 12436
rect 2464 12396 6644 12424
rect 2464 12384 2470 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 9122 12424 9128 12436
rect 6779 12396 9128 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 11296 12396 11621 12424
rect 11296 12384 11302 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 11609 12387 11667 12393
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12066 12424 12072 12436
rect 11940 12396 12072 12424
rect 11940 12384 11946 12396
rect 12066 12384 12072 12396
rect 12124 12424 12130 12436
rect 12710 12424 12716 12436
rect 12124 12396 12716 12424
rect 12124 12384 12130 12396
rect 12710 12384 12716 12396
rect 12768 12424 12774 12436
rect 14458 12424 14464 12436
rect 12768 12396 14464 12424
rect 12768 12384 12774 12396
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 17586 12424 17592 12436
rect 15488 12396 17592 12424
rect 7193 12359 7251 12365
rect 7193 12325 7205 12359
rect 7239 12325 7251 12359
rect 7193 12319 7251 12325
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 5534 12220 5540 12232
rect 3467 12192 5540 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6822 12220 6828 12232
rect 6595 12192 6828 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 3176 12155 3234 12161
rect 3176 12121 3188 12155
rect 3222 12152 3234 12155
rect 3694 12152 3700 12164
rect 3222 12124 3700 12152
rect 3222 12121 3234 12124
rect 3176 12115 3234 12121
rect 3694 12112 3700 12124
rect 3752 12112 3758 12164
rect 3970 12152 3976 12164
rect 3931 12124 3976 12152
rect 3970 12112 3976 12124
rect 4028 12112 4034 12164
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 6196 12152 6224 12183
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7208 12220 7236 12319
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 8720 12328 12633 12356
rect 8720 12316 8726 12328
rect 12621 12325 12633 12328
rect 12667 12325 12679 12359
rect 12621 12319 12679 12325
rect 13633 12359 13691 12365
rect 13633 12325 13645 12359
rect 13679 12356 13691 12359
rect 15488 12356 15516 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 20625 12427 20683 12433
rect 20625 12393 20637 12427
rect 20671 12424 20683 12427
rect 20714 12424 20720 12436
rect 20671 12396 20720 12424
rect 20671 12393 20683 12396
rect 20625 12387 20683 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 22370 12424 22376 12436
rect 22331 12396 22376 12424
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 23569 12427 23627 12433
rect 23569 12393 23581 12427
rect 23615 12424 23627 12427
rect 23842 12424 23848 12436
rect 23615 12396 23848 12424
rect 23615 12393 23627 12396
rect 23569 12387 23627 12393
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 13679 12328 15516 12356
rect 13679 12325 13691 12328
rect 13633 12319 13691 12325
rect 20438 12316 20444 12368
rect 20496 12316 20502 12368
rect 21361 12359 21419 12365
rect 21361 12325 21373 12359
rect 21407 12325 21419 12359
rect 25038 12356 25044 12368
rect 21361 12319 21419 12325
rect 24688 12328 25044 12356
rect 10410 12288 10416 12300
rect 8496 12260 10416 12288
rect 8496 12220 8524 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 15654 12288 15660 12300
rect 12636 12260 13492 12288
rect 15615 12260 15660 12288
rect 7208 12192 8524 12220
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8628 12192 8673 12220
rect 8628 12180 8634 12192
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8996 12192 9137 12220
rect 8996 12180 9002 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9401 12223 9459 12229
rect 9272 12192 9317 12220
rect 9272 12180 9278 12192
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9490 12220 9496 12232
rect 9447 12192 9496 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9490 12180 9496 12192
rect 9548 12220 9554 12232
rect 9674 12220 9680 12232
rect 9548 12192 9680 12220
rect 9548 12180 9554 12192
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 12636 12229 12664 12260
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 10744 12192 12633 12220
rect 10744 12180 10750 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12802 12220 12808 12232
rect 12763 12192 12808 12220
rect 12621 12183 12679 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 4120 12124 6224 12152
rect 6365 12155 6423 12161
rect 4120 12112 4126 12124
rect 6365 12121 6377 12155
rect 6411 12121 6423 12155
rect 6365 12115 6423 12121
rect 6457 12155 6515 12161
rect 6457 12121 6469 12155
rect 6503 12152 6515 12155
rect 7558 12152 7564 12164
rect 6503 12124 7564 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 5258 12084 5264 12096
rect 5219 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 6380 12084 6408 12115
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 8306 12155 8364 12161
rect 8306 12121 8318 12155
rect 8352 12121 8364 12155
rect 8306 12115 8364 12121
rect 6914 12084 6920 12096
rect 6380 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12084 6978 12096
rect 7190 12084 7196 12096
rect 6972 12056 7196 12084
rect 6972 12044 6978 12056
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8312 12084 8340 12115
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 8536 12124 10333 12152
rect 8536 12112 8542 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 10410 12112 10416 12164
rect 10468 12152 10474 12164
rect 13372 12152 13400 12183
rect 10468 12124 13400 12152
rect 10468 12112 10474 12124
rect 9030 12084 9036 12096
rect 8312 12056 9036 12084
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 9548 12056 9597 12084
rect 9548 12044 9554 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 13464 12084 13492 12260
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 16022 12248 16028 12300
rect 16080 12288 16086 12300
rect 19426 12288 19432 12300
rect 16080 12260 19432 12288
rect 16080 12248 16086 12260
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 20070 12288 20076 12300
rect 20031 12260 20076 12288
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 20456 12288 20484 12316
rect 21376 12288 21404 12319
rect 24118 12288 24124 12300
rect 20395 12260 20484 12288
rect 20916 12260 21404 12288
rect 22066 12260 24124 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12220 13691 12223
rect 14090 12220 14096 12232
rect 13679 12192 14096 12220
rect 13679 12189 13691 12192
rect 13633 12183 13691 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14550 12220 14556 12232
rect 14511 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15286 12220 15292 12232
rect 14783 12192 15292 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 14240 12124 14381 12152
rect 14240 12112 14246 12124
rect 14369 12121 14381 12124
rect 14415 12121 14427 12155
rect 15396 12152 15424 12183
rect 16758 12180 16764 12232
rect 16816 12180 16822 12232
rect 17678 12220 17684 12232
rect 17639 12192 17684 12220
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17954 12220 17960 12232
rect 17915 12192 17960 12220
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 19978 12220 19984 12232
rect 19939 12192 19984 12220
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20254 12220 20260 12232
rect 20180 12192 20260 12220
rect 15746 12152 15752 12164
rect 15396 12124 15752 12152
rect 14369 12115 14427 12121
rect 15746 12112 15752 12124
rect 15804 12112 15810 12164
rect 17218 12152 17224 12164
rect 16960 12124 17224 12152
rect 14458 12084 14464 12096
rect 13464 12056 14464 12084
rect 9585 12047 9643 12053
rect 14458 12044 14464 12056
rect 14516 12084 14522 12096
rect 16960 12084 16988 12124
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12152 18107 12155
rect 18138 12152 18144 12164
rect 18095 12124 18144 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18138 12112 18144 12124
rect 18196 12112 18202 12164
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 20180 12152 20208 12192
rect 20254 12180 20260 12192
rect 20312 12180 20318 12232
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 20916 12220 20944 12260
rect 21082 12220 21088 12232
rect 20487 12192 20944 12220
rect 21043 12192 21088 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21266 12220 21272 12232
rect 21223 12192 21272 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12220 21419 12223
rect 21450 12220 21456 12232
rect 21407 12192 21456 12220
rect 21407 12189 21419 12192
rect 21361 12183 21419 12189
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 22066 12152 22094 12260
rect 24118 12248 24124 12260
rect 24176 12248 24182 12300
rect 23106 12220 23112 12232
rect 23067 12192 23112 12220
rect 23106 12180 23112 12192
rect 23164 12180 23170 12232
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 24688 12220 24716 12328
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 25406 12316 25412 12368
rect 25464 12356 25470 12368
rect 25685 12359 25743 12365
rect 25685 12356 25697 12359
rect 25464 12328 25697 12356
rect 25464 12316 25470 12328
rect 25685 12325 25697 12328
rect 25731 12325 25743 12359
rect 25685 12319 25743 12325
rect 24762 12248 24768 12300
rect 24820 12288 24826 12300
rect 24820 12260 25544 12288
rect 24820 12248 24826 12260
rect 24946 12220 24952 12232
rect 23431 12192 24716 12220
rect 24907 12192 24952 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25038 12180 25044 12232
rect 25096 12220 25102 12232
rect 25406 12220 25412 12232
rect 25096 12192 25412 12220
rect 25096 12180 25102 12192
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 25516 12220 25544 12260
rect 25958 12220 25964 12232
rect 25516 12192 25820 12220
rect 25919 12192 25964 12220
rect 23290 12152 23296 12164
rect 18923 12124 20208 12152
rect 20272 12124 22094 12152
rect 22664 12124 23296 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 14516 12056 16988 12084
rect 17129 12087 17187 12093
rect 14516 12044 14522 12056
rect 17129 12053 17141 12087
rect 17175 12084 17187 12087
rect 17770 12084 17776 12096
rect 17175 12056 17776 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18288 12056 18521 12084
rect 18288 12044 18294 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 18677 12087 18735 12093
rect 18677 12053 18689 12087
rect 18723 12084 18735 12087
rect 18966 12084 18972 12096
rect 18723 12056 18972 12084
rect 18723 12053 18735 12056
rect 18677 12047 18735 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 20272 12093 20300 12124
rect 22664 12096 22692 12124
rect 23290 12112 23296 12124
rect 23348 12112 23354 12164
rect 24578 12152 24584 12164
rect 24539 12124 24584 12152
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 24728 12124 24773 12152
rect 24728 12112 24734 12124
rect 25130 12112 25136 12164
rect 25188 12152 25194 12164
rect 25590 12152 25596 12164
rect 25188 12124 25596 12152
rect 25188 12112 25194 12124
rect 25590 12112 25596 12124
rect 25648 12152 25654 12164
rect 25685 12155 25743 12161
rect 25685 12152 25697 12155
rect 25648 12124 25697 12152
rect 25648 12112 25654 12124
rect 25685 12121 25697 12124
rect 25731 12121 25743 12155
rect 25792 12152 25820 12192
rect 25958 12180 25964 12192
rect 26016 12180 26022 12232
rect 25869 12155 25927 12161
rect 25869 12152 25881 12155
rect 25792 12124 25881 12152
rect 25685 12115 25743 12121
rect 25869 12121 25881 12124
rect 25915 12121 25927 12155
rect 25869 12115 25927 12121
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12053 20315 12087
rect 20257 12047 20315 12053
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 21821 12087 21879 12093
rect 21821 12084 21833 12087
rect 20588 12056 21833 12084
rect 20588 12044 20594 12056
rect 21821 12053 21833 12056
rect 21867 12084 21879 12087
rect 22646 12084 22652 12096
rect 21867 12056 22652 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 23382 12084 23388 12096
rect 23247 12056 23388 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 25222 12084 25228 12096
rect 25183 12056 25228 12084
rect 25222 12044 25228 12056
rect 25280 12044 25286 12096
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 2222 11880 2228 11892
rect 2179 11852 2228 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3568 11852 3985 11880
rect 3568 11840 3574 11852
rect 3973 11849 3985 11852
rect 4019 11880 4031 11883
rect 6546 11880 6552 11892
rect 4019 11852 6552 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 8662 11880 8668 11892
rect 7064 11852 8668 11880
rect 7064 11840 7070 11852
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 9272 11852 10701 11880
rect 9272 11840 9278 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 11974 11880 11980 11892
rect 11935 11852 11980 11880
rect 10689 11843 10747 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 19153 11883 19211 11889
rect 19153 11880 19165 11883
rect 13464 11852 19165 11880
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 3786 11812 3792 11824
rect 1811 11784 3792 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 6641 11815 6699 11821
rect 5408 11784 6592 11812
rect 5408 11772 5414 11784
rect 6564 11756 6592 11784
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 6687 11784 9168 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2866 11753 2872 11756
rect 2860 11707 2872 11753
rect 2924 11744 2930 11756
rect 4884 11747 4942 11753
rect 2924 11716 2960 11744
rect 2866 11704 2872 11707
rect 2924 11704 2930 11716
rect 4884 11713 4896 11747
rect 4930 11744 4942 11747
rect 5626 11744 5632 11756
rect 4930 11716 5632 11744
rect 4930 11713 4942 11716
rect 4884 11707 4942 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 6546 11744 6552 11756
rect 6507 11716 6552 11744
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2096 11648 2605 11676
rect 2096 11636 2102 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4396 11648 4629 11676
rect 4396 11636 4402 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6840 11676 6868 11707
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 8582 11747 8640 11753
rect 8582 11744 8594 11747
rect 8352 11716 8594 11744
rect 8352 11704 8358 11716
rect 8582 11713 8594 11716
rect 8628 11713 8640 11747
rect 8582 11707 8640 11713
rect 6420 11648 6868 11676
rect 7009 11679 7067 11685
rect 6420 11636 6426 11648
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 8849 11679 8907 11685
rect 7055 11648 7880 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 5994 11540 6000 11552
rect 5955 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11540 6058 11552
rect 6270 11540 6276 11552
rect 6052 11512 6276 11540
rect 6052 11500 6058 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7558 11540 7564 11552
rect 7515 11512 7564 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7852 11540 7880 11648
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9030 11676 9036 11688
rect 8895 11648 9036 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 8662 11540 8668 11552
rect 7852 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9140 11540 9168 11784
rect 9490 11772 9496 11824
rect 9548 11812 9554 11824
rect 12158 11812 12164 11824
rect 9548 11784 9628 11812
rect 12119 11784 12164 11812
rect 9548 11772 9554 11784
rect 9306 11744 9312 11756
rect 9267 11716 9312 11744
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9600 11753 9628 11784
rect 12158 11772 12164 11784
rect 12216 11772 12222 11824
rect 13464 11821 13492 11852
rect 19153 11849 19165 11852
rect 19199 11849 19211 11883
rect 19153 11843 19211 11849
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 19484 11852 21373 11880
rect 19484 11840 19490 11852
rect 21361 11849 21373 11852
rect 21407 11880 21419 11883
rect 22186 11880 22192 11892
rect 21407 11852 22192 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 22186 11840 22192 11852
rect 22244 11880 22250 11892
rect 22830 11880 22836 11892
rect 22244 11852 22836 11880
rect 22244 11840 22250 11852
rect 22830 11840 22836 11852
rect 22888 11840 22894 11892
rect 24765 11883 24823 11889
rect 24765 11849 24777 11883
rect 24811 11880 24823 11883
rect 25958 11880 25964 11892
rect 24811 11852 25964 11880
rect 24811 11849 24823 11852
rect 24765 11843 24823 11849
rect 13449 11815 13507 11821
rect 13449 11781 13461 11815
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 14182 11772 14188 11824
rect 14240 11772 14246 11824
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 15841 11815 15899 11821
rect 15841 11812 15853 11815
rect 15620 11784 15853 11812
rect 15620 11772 15626 11784
rect 15841 11781 15853 11784
rect 15887 11812 15899 11815
rect 16022 11812 16028 11824
rect 15887 11784 16028 11812
rect 15887 11781 15899 11784
rect 15841 11775 15899 11781
rect 16022 11772 16028 11784
rect 16080 11772 16086 11824
rect 16209 11815 16267 11821
rect 16209 11781 16221 11815
rect 16255 11812 16267 11815
rect 17402 11812 17408 11824
rect 16255 11784 17408 11812
rect 16255 11781 16267 11784
rect 16209 11775 16267 11781
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 18138 11772 18144 11824
rect 18196 11772 18202 11824
rect 18782 11812 18788 11824
rect 18524 11784 18788 11812
rect 9576 11747 9634 11753
rect 9576 11713 9588 11747
rect 9622 11713 9634 11747
rect 9576 11707 9634 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 12618 11744 12624 11756
rect 10100 11716 12624 11744
rect 10100 11704 10106 11716
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12768 11648 13185 11676
rect 12768 11636 12774 11648
rect 13173 11645 13185 11648
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14700 11648 15209 11676
rect 14700 11636 14706 11648
rect 15197 11645 15209 11648
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 16850 11676 16856 11688
rect 15804 11648 16856 11676
rect 15804 11636 15810 11648
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 18524 11676 18552 11784
rect 18782 11772 18788 11784
rect 18840 11772 18846 11824
rect 19794 11812 19800 11824
rect 19306 11784 19800 11812
rect 19150 11704 19156 11756
rect 19208 11744 19214 11756
rect 19208 11716 19253 11744
rect 19208 11704 19214 11716
rect 17175 11648 18552 11676
rect 18601 11679 18659 11685
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 18601 11645 18613 11679
rect 18647 11676 18659 11679
rect 19306 11676 19334 11784
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 19978 11772 19984 11824
rect 20036 11812 20042 11824
rect 23652 11815 23710 11821
rect 20036 11784 22048 11812
rect 20036 11772 20042 11784
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 22020 11753 22048 11784
rect 23652 11781 23664 11815
rect 23698 11812 23710 11815
rect 25222 11812 25228 11824
rect 23698 11784 25228 11812
rect 23698 11781 23710 11784
rect 23652 11775 23710 11781
rect 25222 11772 25228 11784
rect 25280 11772 25286 11824
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 19944 11716 20729 11744
rect 19944 11704 19950 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 22005 11707 22063 11713
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 22520 11716 22753 11744
rect 22520 11704 22526 11716
rect 22741 11713 22753 11716
rect 22787 11744 22799 11747
rect 23474 11744 23480 11756
rect 22787 11716 23480 11744
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23474 11704 23480 11716
rect 23532 11744 23538 11756
rect 25608 11753 25636 11852
rect 25958 11840 25964 11852
rect 26016 11880 26022 11892
rect 26329 11883 26387 11889
rect 26329 11880 26341 11883
rect 26016 11852 26341 11880
rect 26016 11840 26022 11852
rect 26329 11849 26341 11852
rect 26375 11849 26387 11883
rect 26329 11843 26387 11849
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 23532 11716 25513 11744
rect 23532 11704 23538 11716
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11744 25835 11747
rect 26050 11744 26056 11756
rect 25823 11716 26056 11744
rect 25823 11713 25835 11716
rect 25777 11707 25835 11713
rect 26050 11704 26056 11716
rect 26108 11704 26114 11756
rect 18647 11648 19334 11676
rect 20257 11679 20315 11685
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 21358 11676 21364 11688
rect 20303 11648 21364 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 21358 11636 21364 11648
rect 21416 11676 21422 11688
rect 22094 11676 22100 11688
rect 21416 11648 22100 11676
rect 21416 11636 21422 11648
rect 22094 11636 22100 11648
rect 22152 11636 22158 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 22756 11648 23397 11676
rect 22756 11620 22784 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25685 11679 25743 11685
rect 25685 11676 25697 11679
rect 24912 11648 25697 11676
rect 24912 11636 24918 11648
rect 25685 11645 25697 11648
rect 25731 11676 25743 11679
rect 25866 11676 25872 11688
rect 25731 11648 25872 11676
rect 25731 11645 25743 11648
rect 25685 11639 25743 11645
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 19978 11608 19984 11620
rect 18616 11580 19984 11608
rect 10502 11540 10508 11552
rect 9140 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11540 10566 11552
rect 10778 11540 10784 11552
rect 10560 11512 10784 11540
rect 10560 11500 10566 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12066 11540 12072 11552
rect 12023 11512 12072 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18616 11540 18644 11580
rect 19978 11568 19984 11580
rect 20036 11608 20042 11620
rect 20165 11611 20223 11617
rect 20165 11608 20177 11611
rect 20036 11580 20177 11608
rect 20036 11568 20042 11580
rect 20165 11577 20177 11580
rect 20211 11577 20223 11611
rect 20806 11608 20812 11620
rect 20767 11580 20812 11608
rect 20165 11571 20223 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 22738 11568 22744 11620
rect 22796 11568 22802 11620
rect 24394 11568 24400 11620
rect 24452 11608 24458 11620
rect 25317 11611 25375 11617
rect 25317 11608 25329 11611
rect 24452 11580 25329 11608
rect 24452 11568 24458 11580
rect 25317 11577 25329 11580
rect 25363 11577 25375 11611
rect 25317 11571 25375 11577
rect 17828 11512 18644 11540
rect 17828 11500 17834 11512
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 20070 11540 20076 11552
rect 18748 11512 20076 11540
rect 18748 11500 18754 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 22097 11543 22155 11549
rect 22097 11509 22109 11543
rect 22143 11540 22155 11543
rect 22186 11540 22192 11552
rect 22143 11512 22192 11540
rect 22143 11509 22155 11512
rect 22097 11503 22155 11509
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 22833 11543 22891 11549
rect 22833 11509 22845 11543
rect 22879 11540 22891 11543
rect 23658 11540 23664 11552
rect 22879 11512 23664 11540
rect 22879 11509 22891 11512
rect 22833 11503 22891 11509
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 6178 11336 6184 11348
rect 5767 11308 6184 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 11330 11336 11336 11348
rect 8619 11308 11336 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 14550 11336 14556 11348
rect 13096 11308 14556 11336
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 10873 11271 10931 11277
rect 10873 11268 10885 11271
rect 10836 11240 10885 11268
rect 10836 11228 10842 11240
rect 10873 11237 10885 11240
rect 10919 11237 10931 11271
rect 10873 11231 10931 11237
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8628 11172 9505 11200
rect 8628 11160 8634 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 13096 11200 13124 11308
rect 14550 11296 14556 11308
rect 14608 11336 14614 11348
rect 14967 11339 15025 11345
rect 14967 11336 14979 11339
rect 14608 11308 14979 11336
rect 14608 11296 14614 11308
rect 14967 11305 14979 11308
rect 15013 11305 15025 11339
rect 14967 11299 15025 11305
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 16908 11308 18000 11336
rect 16908 11296 16914 11308
rect 13449 11271 13507 11277
rect 13449 11237 13461 11271
rect 13495 11268 13507 11271
rect 13998 11268 14004 11280
rect 13495 11240 14004 11268
rect 13495 11237 13507 11240
rect 13449 11231 13507 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 17865 11271 17923 11277
rect 17865 11237 17877 11271
rect 17911 11237 17923 11271
rect 17972 11268 18000 11308
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 19886 11336 19892 11348
rect 19668 11308 19892 11336
rect 19668 11296 19674 11308
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 21634 11336 21640 11348
rect 20312 11308 21128 11336
rect 21595 11308 21640 11336
rect 20312 11296 20318 11308
rect 20993 11271 21051 11277
rect 20993 11268 21005 11271
rect 17972 11240 21005 11268
rect 17865 11231 17923 11237
rect 20993 11237 21005 11240
rect 21039 11237 21051 11271
rect 21100 11268 21128 11308
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23937 11339 23995 11345
rect 23937 11305 23949 11339
rect 23983 11336 23995 11339
rect 24670 11336 24676 11348
rect 23983 11308 24676 11336
rect 23983 11305 23995 11308
rect 23937 11299 23995 11305
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 24854 11336 24860 11348
rect 24780 11308 24860 11336
rect 24780 11268 24808 11308
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25130 11336 25136 11348
rect 25091 11308 25136 11336
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 25685 11271 25743 11277
rect 25685 11268 25697 11271
rect 21100 11240 24808 11268
rect 24872 11240 25697 11268
rect 20993 11231 21051 11237
rect 12023 11172 13124 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 15286 11200 15292 11212
rect 13228 11172 15292 11200
rect 13228 11160 13234 11172
rect 15286 11160 15292 11172
rect 15344 11200 15350 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15344 11172 15669 11200
rect 15344 11160 15350 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 8386 11132 8392 11144
rect 8299 11104 8392 11132
rect 8386 11092 8392 11104
rect 8444 11132 8450 11144
rect 8444 11104 9904 11132
rect 8444 11092 8450 11104
rect 9876 11076 9904 11104
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11112 11104 11713 11132
rect 11112 11092 11118 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11132 15255 11135
rect 17880 11132 17908 11231
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 18012 11172 18429 11200
rect 18012 11160 18018 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 19978 11200 19984 11212
rect 19939 11172 19984 11200
rect 18417 11163 18475 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 23106 11200 23112 11212
rect 20088 11172 23112 11200
rect 15243 11104 17908 11132
rect 15243 11101 15255 11104
rect 15197 11095 15255 11101
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 18104 11104 18245 11132
rect 18104 11092 18110 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 20088 11132 20116 11172
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 23492 11200 23520 11240
rect 23566 11200 23572 11212
rect 23492 11172 23572 11200
rect 18371 11104 20116 11132
rect 20165 11135 20223 11141
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 20165 11101 20177 11135
rect 20211 11132 20223 11135
rect 20254 11132 20260 11144
rect 20211 11104 20260 11132
rect 20211 11101 20223 11104
rect 20165 11095 20223 11101
rect 3329 11067 3387 11073
rect 3329 11033 3341 11067
rect 3375 11064 3387 11067
rect 4608 11067 4666 11073
rect 3375 11036 4568 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 4540 10996 4568 11036
rect 4608 11033 4620 11067
rect 4654 11064 4666 11067
rect 4706 11064 4712 11076
rect 4654 11036 4712 11064
rect 4654 11033 4666 11036
rect 4608 11027 4666 11033
rect 4706 11024 4712 11036
rect 4764 11024 4770 11076
rect 6181 11067 6239 11073
rect 6181 11033 6193 11067
rect 6227 11064 6239 11067
rect 6730 11064 6736 11076
rect 6227 11036 6736 11064
rect 6227 11033 6239 11036
rect 6181 11027 6239 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 7300 11036 7604 11064
rect 5258 10996 5264 11008
rect 4540 10968 5264 10996
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6546 10956 6552 11008
rect 6604 10996 6610 11008
rect 7300 10996 7328 11036
rect 7466 10996 7472 11008
rect 6604 10968 7328 10996
rect 7427 10968 7472 10996
rect 6604 10956 6610 10968
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7576 10996 7604 11036
rect 8128 11036 8616 11064
rect 8128 10996 8156 11036
rect 7576 10968 8156 10996
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8386 10996 8392 11008
rect 8260 10968 8392 10996
rect 8260 10956 8266 10968
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 8588 10996 8616 11036
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9738 11067 9796 11073
rect 9738 11064 9750 11067
rect 8720 11036 9750 11064
rect 8720 11024 8726 11036
rect 9738 11033 9750 11036
rect 9784 11033 9796 11067
rect 9738 11027 9796 11033
rect 9858 11024 9864 11076
rect 9916 11024 9922 11076
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 10836 11036 11928 11064
rect 10836 11024 10842 11036
rect 10502 10996 10508 11008
rect 8588 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 11900 10996 11928 11036
rect 12084 11036 12466 11064
rect 12084 10996 12112 11036
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 17405 11067 17463 11073
rect 14700 11036 17356 11064
rect 14700 11024 14706 11036
rect 11900 10968 12112 10996
rect 17328 10996 17356 11036
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 17954 11064 17960 11076
rect 17451 11036 17960 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 19150 11064 19156 11076
rect 18064 11036 19156 11064
rect 18064 10996 18092 11036
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 19242 11024 19248 11076
rect 19300 11064 19306 11076
rect 19794 11064 19800 11076
rect 19300 11036 19800 11064
rect 19300 11024 19306 11036
rect 19794 11024 19800 11036
rect 19852 11064 19858 11076
rect 19889 11067 19947 11073
rect 19889 11064 19901 11067
rect 19852 11036 19901 11064
rect 19852 11024 19858 11036
rect 19889 11033 19901 11036
rect 19935 11033 19947 11067
rect 20180 11064 20208 11095
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21266 11132 21272 11144
rect 21131 11104 21272 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 21508 11104 21557 11132
rect 21508 11092 21514 11104
rect 21545 11101 21557 11104
rect 21591 11101 21603 11135
rect 21545 11095 21603 11101
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 21744 11064 21772 11095
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22189 11135 22247 11141
rect 22189 11132 22201 11135
rect 22152 11104 22201 11132
rect 22152 11092 22158 11104
rect 22189 11101 22201 11104
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11132 22431 11135
rect 23492 11132 23520 11172
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 24302 11160 24308 11212
rect 24360 11200 24366 11212
rect 24872 11209 24900 11240
rect 25685 11237 25697 11240
rect 25731 11237 25743 11271
rect 25685 11231 25743 11237
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24360 11172 24869 11200
rect 24360 11160 24366 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 23658 11132 23664 11144
rect 22419 11104 23520 11132
rect 23619 11104 23664 11132
rect 22419 11101 22431 11104
rect 22373 11095 22431 11101
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11132 23995 11135
rect 24394 11132 24400 11144
rect 23983 11104 24400 11132
rect 23983 11101 23995 11104
rect 23937 11095 23995 11101
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24762 11132 24768 11144
rect 24723 11104 24768 11132
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 25130 11092 25136 11144
rect 25188 11132 25194 11144
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 25188 11104 25605 11132
rect 25188 11092 25194 11104
rect 25593 11101 25605 11104
rect 25639 11132 25651 11135
rect 25682 11132 25688 11144
rect 25639 11104 25688 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 25682 11092 25688 11104
rect 25740 11092 25746 11144
rect 25777 11135 25835 11141
rect 25777 11101 25789 11135
rect 25823 11132 25835 11135
rect 25866 11132 25872 11144
rect 25823 11104 25872 11132
rect 25823 11101 25835 11104
rect 25777 11095 25835 11101
rect 25866 11092 25872 11104
rect 25924 11132 25930 11144
rect 26789 11135 26847 11141
rect 26789 11132 26801 11135
rect 25924 11104 26801 11132
rect 25924 11092 25930 11104
rect 26789 11101 26801 11104
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 19889 11027 19947 11033
rect 19996 11036 20208 11064
rect 20364 11036 24164 11064
rect 17328 10968 18092 10996
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19996 10996 20024 11036
rect 19484 10968 20024 10996
rect 19484 10956 19490 10968
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 20364 11005 20392 11036
rect 20349 10999 20407 11005
rect 20349 10996 20361 10999
rect 20220 10968 20361 10996
rect 20220 10956 20226 10968
rect 20349 10965 20361 10968
rect 20395 10965 20407 10999
rect 20349 10959 20407 10965
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 21450 10996 21456 11008
rect 20772 10968 21456 10996
rect 20772 10956 20778 10968
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 22278 10996 22284 11008
rect 22239 10968 22284 10996
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 23750 10996 23756 11008
rect 23711 10968 23756 10996
rect 23750 10956 23756 10968
rect 23808 10956 23814 11008
rect 24136 10996 24164 11036
rect 24210 11024 24216 11076
rect 24268 11064 24274 11076
rect 26237 11067 26295 11073
rect 26237 11064 26249 11067
rect 24268 11036 26249 11064
rect 24268 11024 24274 11036
rect 26237 11033 26249 11036
rect 26283 11033 26295 11067
rect 26237 11027 26295 11033
rect 25130 10996 25136 11008
rect 24136 10968 25136 10996
rect 25130 10956 25136 10968
rect 25188 10956 25194 11008
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 4338 10792 4344 10804
rect 3099 10764 4344 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4890 10792 4896 10804
rect 4764 10764 4896 10792
rect 4764 10752 4770 10764
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5442 10792 5448 10804
rect 5031 10764 5448 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5718 10792 5724 10804
rect 5583 10764 5724 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5902 10792 5908 10804
rect 5863 10764 5908 10792
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7282 10792 7288 10804
rect 7055 10764 7288 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7432 10764 7573 10792
rect 7432 10752 7438 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 12710 10792 12716 10804
rect 9824 10764 12716 10792
rect 9824 10752 9830 10764
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 12851 10764 16896 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 1765 10727 1823 10733
rect 1765 10693 1777 10727
rect 1811 10724 1823 10727
rect 2774 10724 2780 10736
rect 1811 10696 2780 10724
rect 1811 10693 1823 10696
rect 1765 10687 1823 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 7466 10724 7472 10736
rect 4356 10696 7472 10724
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 3602 10656 3608 10668
rect 1995 10628 3608 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4356 10665 4384 10696
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 5074 10656 5080 10668
rect 5035 10628 5080 10656
rect 4893 10619 4951 10625
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 4908 10588 4936 10619
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5368 10600 5396 10696
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 8696 10727 8754 10733
rect 8696 10693 8708 10727
rect 8742 10724 8754 10727
rect 10962 10724 10968 10736
rect 8742 10696 10968 10724
rect 8742 10693 8754 10696
rect 8696 10687 8754 10693
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11149 10727 11207 10733
rect 11149 10693 11161 10727
rect 11195 10724 11207 10727
rect 11238 10724 11244 10736
rect 11195 10696 11244 10724
rect 11195 10693 11207 10696
rect 11149 10687 11207 10693
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 16868 10733 16896 10764
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 17460 10764 19625 10792
rect 17460 10752 17466 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 11388 10696 13277 10724
rect 11388 10684 11394 10696
rect 13265 10693 13277 10696
rect 13311 10693 13323 10727
rect 13265 10687 13323 10693
rect 16853 10727 16911 10733
rect 16853 10693 16865 10727
rect 16899 10693 16911 10727
rect 16853 10687 16911 10693
rect 5718 10656 5724 10668
rect 5679 10628 5724 10656
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 5997 10619 6055 10625
rect 3936 10560 4936 10588
rect 3936 10548 3942 10560
rect 4908 10520 4936 10560
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 6012 10588 6040 10619
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 8846 10656 8852 10668
rect 7944 10628 8852 10656
rect 7116 10588 7144 10616
rect 6012 10560 7144 10588
rect 7944 10520 7972 10628
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9030 10656 9036 10668
rect 8987 10628 9036 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9030 10616 9036 10628
rect 9088 10656 9094 10668
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 9088 10628 9413 10656
rect 9088 10616 9094 10628
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 10560 10628 11713 10656
rect 10560 10616 10566 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 11882 10656 11888 10668
rect 11839 10628 11888 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12066 10656 12072 10668
rect 12023 10628 12072 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12216 10628 12633 10656
rect 12216 10616 12222 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 18874 10616 18880 10668
rect 18932 10656 18938 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18932 10628 19073 10656
rect 18932 10616 18938 10628
rect 19061 10625 19073 10628
rect 19107 10625 19119 10659
rect 19426 10656 19432 10668
rect 19387 10628 19432 10656
rect 19061 10619 19119 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19628 10656 19656 10755
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20898 10792 20904 10804
rect 19944 10764 20904 10792
rect 19944 10752 19950 10764
rect 20898 10752 20904 10764
rect 20956 10792 20962 10804
rect 20993 10795 21051 10801
rect 20993 10792 21005 10795
rect 20956 10764 21005 10792
rect 20956 10752 20962 10764
rect 20993 10761 21005 10764
rect 21039 10761 21051 10795
rect 20993 10755 21051 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21453 10795 21511 10801
rect 21453 10792 21465 10795
rect 21140 10764 21465 10792
rect 21140 10752 21146 10764
rect 21453 10761 21465 10764
rect 21499 10761 21511 10795
rect 21453 10755 21511 10761
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 21818 10792 21824 10804
rect 21600 10764 21824 10792
rect 21600 10752 21606 10764
rect 21818 10752 21824 10764
rect 21876 10792 21882 10804
rect 24305 10795 24363 10801
rect 21876 10764 24256 10792
rect 21876 10752 21882 10764
rect 20180 10696 22232 10724
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19628 10628 20085 10656
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 8864 10588 8892 10616
rect 10042 10588 10048 10600
rect 8864 10560 10048 10588
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15344 10560 16037 10588
rect 15344 10548 15350 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 16666 10588 16672 10600
rect 16347 10560 16672 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 4908 10492 7972 10520
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 12032 10492 12173 10520
rect 12032 10480 12038 10492
rect 12161 10489 12173 10492
rect 12207 10489 12219 10523
rect 20180 10520 20208 10696
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20530 10656 20536 10668
rect 20303 10628 20536 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10656 21146 10668
rect 22204 10665 22232 10696
rect 22922 10684 22928 10736
rect 22980 10724 22986 10736
rect 23477 10727 23535 10733
rect 23477 10724 23489 10727
rect 22980 10696 23489 10724
rect 22980 10684 22986 10696
rect 23477 10693 23489 10696
rect 23523 10724 23535 10727
rect 24118 10724 24124 10736
rect 23523 10696 24124 10724
rect 23523 10693 23535 10696
rect 23477 10687 23535 10693
rect 24118 10684 24124 10696
rect 24176 10684 24182 10736
rect 24228 10724 24256 10764
rect 24305 10761 24317 10795
rect 24351 10792 24363 10795
rect 24578 10792 24584 10804
rect 24351 10764 24584 10792
rect 24351 10761 24363 10764
rect 24305 10755 24363 10761
rect 24578 10752 24584 10764
rect 24636 10752 24642 10804
rect 25501 10727 25559 10733
rect 25501 10724 25513 10727
rect 24228 10696 25513 10724
rect 25501 10693 25513 10696
rect 25547 10724 25559 10727
rect 26142 10724 26148 10736
rect 25547 10696 26148 10724
rect 25547 10693 25559 10696
rect 25501 10687 25559 10693
rect 26142 10684 26148 10696
rect 26200 10684 26206 10736
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21140 10628 22017 10656
rect 21140 10616 21146 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22370 10656 22376 10668
rect 22235 10628 22376 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22370 10616 22376 10628
rect 22428 10616 22434 10668
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 23385 10659 23443 10665
rect 23385 10656 23397 10659
rect 23348 10628 23397 10656
rect 23348 10616 23354 10628
rect 23385 10625 23397 10628
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 12161 10483 12219 10489
rect 19352 10492 20208 10520
rect 20916 10520 20944 10551
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 23750 10588 23756 10600
rect 21048 10560 23756 10588
rect 21048 10548 21054 10560
rect 23750 10548 23756 10560
rect 23808 10588 23814 10600
rect 24044 10588 24072 10619
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24728 10628 25053 10656
rect 24728 10616 24734 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 24302 10588 24308 10600
rect 23808 10560 24072 10588
rect 24263 10560 24308 10588
rect 23808 10548 23814 10560
rect 24302 10548 24308 10560
rect 24360 10548 24366 10600
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 24636 10560 24777 10588
rect 24636 10548 24642 10560
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 22278 10520 22284 10532
rect 20916 10492 22284 10520
rect 19352 10464 19380 10492
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 22646 10480 22652 10532
rect 22704 10520 22710 10532
rect 22741 10523 22799 10529
rect 22741 10520 22753 10523
rect 22704 10492 22753 10520
rect 22704 10480 22710 10492
rect 22741 10489 22753 10492
rect 22787 10520 22799 10523
rect 22787 10492 23612 10520
rect 22787 10489 22799 10492
rect 22741 10483 22799 10489
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 10502 10452 10508 10464
rect 7432 10424 10508 10452
rect 7432 10412 7438 10424
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 13964 10424 14565 10452
rect 13964 10412 13970 10424
rect 14553 10421 14565 10424
rect 14599 10421 14611 10455
rect 14553 10415 14611 10421
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 18012 10424 18153 10452
rect 18012 10412 18018 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 19334 10452 19340 10464
rect 19295 10424 19340 10452
rect 18141 10415 18199 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19576 10424 20085 10452
rect 19576 10412 19582 10424
rect 20073 10421 20085 10424
rect 20119 10421 20131 10455
rect 20073 10415 20131 10421
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 21174 10452 21180 10464
rect 20312 10424 21180 10452
rect 20312 10412 20318 10424
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21600 10424 22017 10452
rect 21600 10412 21606 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 23584 10452 23612 10492
rect 23658 10480 23664 10532
rect 23716 10520 23722 10532
rect 24121 10523 24179 10529
rect 24121 10520 24133 10523
rect 23716 10492 24133 10520
rect 23716 10480 23722 10492
rect 24121 10489 24133 10492
rect 24167 10489 24179 10523
rect 26053 10523 26111 10529
rect 26053 10520 26065 10523
rect 24121 10483 24179 10489
rect 24228 10492 26065 10520
rect 24228 10452 24256 10492
rect 26053 10489 26065 10492
rect 26099 10489 26111 10523
rect 26053 10483 26111 10489
rect 24854 10452 24860 10464
rect 23584 10424 24256 10452
rect 24815 10424 24860 10452
rect 22005 10415 22063 10421
rect 24854 10412 24860 10424
rect 24912 10412 24918 10464
rect 24946 10412 24952 10464
rect 25004 10452 25010 10464
rect 25004 10424 25049 10452
rect 25004 10412 25010 10424
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 2740 10220 4261 10248
rect 2740 10208 2746 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 5592 10220 6561 10248
rect 5592 10208 5598 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 9582 10248 9588 10260
rect 7699 10220 9588 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 12066 10248 12072 10260
rect 9732 10220 12072 10248
rect 9732 10208 9738 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 12216 10220 12449 10248
rect 12216 10208 12222 10220
rect 12437 10217 12449 10220
rect 12483 10217 12495 10251
rect 16666 10248 16672 10260
rect 12437 10211 12495 10217
rect 14292 10220 16528 10248
rect 16627 10220 16672 10248
rect 8018 10180 8024 10192
rect 6564 10152 8024 10180
rect 6564 10124 6592 10152
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 8113 10183 8171 10189
rect 8113 10149 8125 10183
rect 8159 10180 8171 10183
rect 8294 10180 8300 10192
rect 8159 10152 8300 10180
rect 8159 10149 8171 10152
rect 8113 10143 8171 10149
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 9217 10183 9275 10189
rect 9217 10149 9229 10183
rect 9263 10180 9275 10183
rect 10410 10180 10416 10192
rect 9263 10152 10416 10180
rect 9263 10149 9275 10152
rect 9217 10143 9275 10149
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 6362 10112 6368 10124
rect 4448 10084 6368 10112
rect 3326 10044 3332 10056
rect 3287 10016 3332 10044
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4448 10053 4476 10084
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6546 10072 6552 10124
rect 6604 10072 6610 10124
rect 10594 10112 10600 10124
rect 7668 10084 10600 10112
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4212 10016 4445 10044
rect 4212 10004 4218 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 4709 10007 4767 10013
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 4617 9979 4675 9985
rect 4617 9976 4629 9979
rect 4304 9948 4629 9976
rect 4304 9936 4310 9948
rect 4617 9945 4629 9948
rect 4663 9945 4675 9979
rect 4617 9939 4675 9945
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 4724 9908 4752 10007
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 7469 10046 7527 10049
rect 7668 10046 7696 10084
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 7469 10043 7696 10046
rect 7469 10009 7481 10043
rect 7515 10018 7696 10043
rect 7515 10009 7527 10018
rect 7469 10003 7527 10009
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8076 10016 8309 10044
rect 8076 10004 8082 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8938 10044 8944 10056
rect 8619 10016 8944 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 13725 10047 13783 10053
rect 9171 10016 10732 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 7098 9976 7104 9988
rect 5092 9948 7104 9976
rect 5092 9920 5120 9948
rect 7098 9936 7104 9948
rect 7156 9976 7162 9988
rect 7374 9976 7380 9988
rect 7156 9948 7380 9976
rect 7156 9936 7162 9948
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 7558 9936 7564 9988
rect 7616 9976 7622 9988
rect 8481 9979 8539 9985
rect 8481 9976 8493 9979
rect 7616 9948 8493 9976
rect 7616 9936 7622 9948
rect 8481 9945 8493 9948
rect 8527 9945 8539 9979
rect 9766 9976 9772 9988
rect 9727 9948 9772 9976
rect 8481 9939 8539 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 5074 9908 5080 9920
rect 1728 9880 5080 9908
rect 1728 9868 1734 9880
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 9582 9908 9588 9920
rect 6880 9880 9588 9908
rect 6880 9868 6886 9880
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10704 9908 10732 10016
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 13906 10044 13912 10056
rect 13771 10016 13912 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 13814 9976 13820 9988
rect 11563 9948 13820 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 12802 9908 12808 9920
rect 10704 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9908 12866 9920
rect 14292 9908 14320 10220
rect 16500 10180 16528 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 21085 10251 21143 10257
rect 21085 10217 21097 10251
rect 21131 10248 21143 10251
rect 21542 10248 21548 10260
rect 21131 10220 21548 10248
rect 21131 10217 21143 10220
rect 21085 10211 21143 10217
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 21821 10251 21879 10257
rect 21821 10248 21833 10251
rect 21784 10220 21833 10248
rect 21784 10208 21790 10220
rect 21821 10217 21833 10220
rect 21867 10217 21879 10251
rect 21821 10211 21879 10217
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 24581 10251 24639 10257
rect 22704 10220 23336 10248
rect 22704 10208 22710 10220
rect 17402 10180 17408 10192
rect 16500 10152 17408 10180
rect 17402 10140 17408 10152
rect 17460 10140 17466 10192
rect 21637 10183 21695 10189
rect 21637 10180 21649 10183
rect 21100 10152 21649 10180
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10112 14427 10115
rect 15194 10112 15200 10124
rect 14415 10084 15200 10112
rect 14415 10081 14427 10084
rect 14369 10075 14427 10081
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 17218 10112 17224 10124
rect 16163 10084 17224 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 17328 10084 18337 10112
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17328 10044 17356 10084
rect 18325 10081 18337 10084
rect 18371 10081 18383 10115
rect 21100 10112 21128 10152
rect 21637 10149 21649 10152
rect 21683 10149 21695 10183
rect 21637 10143 21695 10149
rect 23017 10183 23075 10189
rect 23017 10149 23029 10183
rect 23063 10180 23075 10183
rect 23106 10180 23112 10192
rect 23063 10152 23112 10180
rect 23063 10149 23075 10152
rect 23017 10143 23075 10149
rect 23106 10140 23112 10152
rect 23164 10140 23170 10192
rect 23308 10180 23336 10220
rect 24581 10217 24593 10251
rect 24627 10248 24639 10251
rect 24670 10248 24676 10260
rect 24627 10220 24676 10248
rect 24627 10217 24639 10220
rect 24581 10211 24639 10217
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 24765 10251 24823 10257
rect 24765 10217 24777 10251
rect 24811 10248 24823 10251
rect 25130 10248 25136 10260
rect 24811 10220 25136 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 25130 10208 25136 10220
rect 25188 10208 25194 10260
rect 26142 10208 26148 10260
rect 26200 10248 26206 10260
rect 26697 10251 26755 10257
rect 26697 10248 26709 10251
rect 26200 10220 26709 10248
rect 26200 10208 26206 10220
rect 26697 10217 26709 10220
rect 26743 10217 26755 10251
rect 26697 10211 26755 10217
rect 25409 10183 25467 10189
rect 25409 10180 25421 10183
rect 23308 10152 25421 10180
rect 25409 10149 25421 10152
rect 25455 10149 25467 10183
rect 25409 10143 25467 10149
rect 25866 10140 25872 10192
rect 25924 10180 25930 10192
rect 27249 10183 27307 10189
rect 27249 10180 27261 10183
rect 25924 10152 27261 10180
rect 25924 10140 25930 10152
rect 27249 10149 27261 10152
rect 27295 10149 27307 10183
rect 27249 10143 27307 10149
rect 18325 10075 18383 10081
rect 20824 10084 21128 10112
rect 18046 10044 18052 10056
rect 17092 10016 17356 10044
rect 18007 10016 18052 10044
rect 17092 10004 17098 10016
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 19886 10044 19892 10056
rect 19847 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20824 10053 20852 10084
rect 23474 10072 23480 10124
rect 23532 10112 23538 10124
rect 23569 10115 23627 10121
rect 23569 10112 23581 10115
rect 23532 10084 23581 10112
rect 23532 10072 23538 10084
rect 23569 10081 23581 10084
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10044 20131 10047
rect 20809 10047 20867 10053
rect 20119 10016 20760 10044
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 14645 9979 14703 9985
rect 14645 9945 14657 9979
rect 14691 9945 14703 9979
rect 14645 9939 14703 9945
rect 12860 9880 14320 9908
rect 14660 9908 14688 9939
rect 14734 9936 14740 9988
rect 14792 9976 14798 9988
rect 17129 9979 17187 9985
rect 14792 9948 15134 9976
rect 14792 9936 14798 9948
rect 17129 9945 17141 9979
rect 17175 9976 17187 9979
rect 18690 9976 18696 9988
rect 17175 9948 18696 9976
rect 17175 9945 17187 9948
rect 17129 9939 17187 9945
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 20162 9976 20168 9988
rect 20123 9948 20168 9976
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 16022 9908 16028 9920
rect 14660 9880 16028 9908
rect 12860 9868 12866 9880
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17037 9911 17095 9917
rect 17037 9908 17049 9911
rect 16724 9880 17049 9908
rect 16724 9868 16730 9880
rect 17037 9877 17049 9880
rect 17083 9908 17095 9911
rect 19794 9908 19800 9920
rect 17083 9880 19800 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 19794 9868 19800 9880
rect 19852 9868 19858 9920
rect 20254 9868 20260 9920
rect 20312 9908 20318 9920
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20312 9880 20637 9908
rect 20312 9868 20318 9880
rect 20625 9877 20637 9880
rect 20671 9877 20683 9911
rect 20732 9908 20760 10016
rect 20809 10013 20821 10047
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 20898 10004 20904 10056
rect 20956 10044 20962 10056
rect 21174 10044 21180 10056
rect 20956 10016 21001 10044
rect 21135 10016 21180 10044
rect 20956 10004 20962 10016
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21818 10044 21824 10056
rect 21779 10016 21824 10044
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10044 22799 10047
rect 22830 10044 22836 10056
rect 22787 10016 22836 10044
rect 22787 10013 22799 10016
rect 22741 10007 22799 10013
rect 20990 9936 20996 9988
rect 21048 9976 21054 9988
rect 21634 9976 21640 9988
rect 21048 9948 21640 9976
rect 21048 9936 21054 9948
rect 21634 9936 21640 9948
rect 21692 9976 21698 9988
rect 21928 9976 21956 10007
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 23382 10004 23388 10056
rect 23440 10044 23446 10056
rect 23661 10047 23719 10053
rect 23661 10044 23673 10047
rect 23440 10016 23673 10044
rect 23440 10004 23446 10016
rect 23661 10013 23673 10016
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 24912 10016 25697 10044
rect 24912 10004 24918 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 21692 9948 21956 9976
rect 22097 9979 22155 9985
rect 21692 9936 21698 9948
rect 22097 9945 22109 9979
rect 22143 9976 22155 9979
rect 22462 9976 22468 9988
rect 22143 9948 22468 9976
rect 22143 9945 22155 9948
rect 22097 9939 22155 9945
rect 22462 9936 22468 9948
rect 22520 9936 22526 9988
rect 23017 9979 23075 9985
rect 23017 9945 23029 9979
rect 23063 9976 23075 9979
rect 23934 9976 23940 9988
rect 23063 9948 23940 9976
rect 23063 9945 23075 9948
rect 23017 9939 23075 9945
rect 23934 9936 23940 9948
rect 23992 9936 23998 9988
rect 24762 9985 24768 9988
rect 24749 9979 24768 9985
rect 24749 9976 24761 9979
rect 24044 9948 24761 9976
rect 22186 9908 22192 9920
rect 20732 9880 22192 9908
rect 20625 9871 20683 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22833 9911 22891 9917
rect 22833 9908 22845 9911
rect 22428 9880 22845 9908
rect 22428 9868 22434 9880
rect 22833 9877 22845 9880
rect 22879 9908 22891 9911
rect 23382 9908 23388 9920
rect 22879 9880 23388 9908
rect 22879 9877 22891 9880
rect 22833 9871 22891 9877
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 24044 9917 24072 9948
rect 24749 9945 24761 9948
rect 24749 9939 24768 9945
rect 24762 9936 24768 9939
rect 24820 9936 24826 9988
rect 24949 9979 25007 9985
rect 24949 9945 24961 9979
rect 24995 9976 25007 9979
rect 25038 9976 25044 9988
rect 24995 9948 25044 9976
rect 24995 9945 25007 9948
rect 24949 9939 25007 9945
rect 25038 9936 25044 9948
rect 25096 9936 25102 9988
rect 25409 9979 25467 9985
rect 25409 9945 25421 9979
rect 25455 9945 25467 9979
rect 25409 9939 25467 9945
rect 24029 9911 24087 9917
rect 24029 9877 24041 9911
rect 24075 9877 24087 9911
rect 24029 9871 24087 9877
rect 24118 9868 24124 9920
rect 24176 9908 24182 9920
rect 25424 9908 25452 9939
rect 25590 9908 25596 9920
rect 24176 9880 25452 9908
rect 25551 9880 25596 9908
rect 24176 9868 24182 9880
rect 25590 9868 25596 9880
rect 25648 9868 25654 9920
rect 26234 9908 26240 9920
rect 26195 9880 26240 9908
rect 26234 9868 26240 9880
rect 26292 9868 26298 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 6822 9704 6828 9716
rect 2004 9676 6828 9704
rect 2004 9664 2010 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 7929 9707 7987 9713
rect 7929 9673 7941 9707
rect 7975 9673 7987 9707
rect 7929 9667 7987 9673
rect 4617 9639 4675 9645
rect 4617 9605 4629 9639
rect 4663 9636 4675 9639
rect 4706 9636 4712 9648
rect 4663 9608 4712 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5166 9636 5172 9648
rect 5031 9608 5172 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5813 9639 5871 9645
rect 5813 9605 5825 9639
rect 5859 9605 5871 9639
rect 5813 9599 5871 9605
rect 5997 9639 6055 9645
rect 5997 9605 6009 9639
rect 6043 9636 6055 9639
rect 6086 9636 6092 9648
rect 6043 9608 6092 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2308 9571 2366 9577
rect 2308 9537 2320 9571
rect 2354 9568 2366 9571
rect 3326 9568 3332 9580
rect 2354 9540 3332 9568
rect 2354 9537 2366 9540
rect 2308 9531 2366 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 4798 9568 4804 9580
rect 4759 9540 4804 9568
rect 3973 9531 4031 9537
rect 3988 9500 4016 9531
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5828 9568 5856 9599
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 7944 9636 7972 9667
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 14645 9707 14703 9713
rect 14645 9704 14657 9707
rect 13872 9676 14657 9704
rect 13872 9664 13878 9676
rect 14645 9673 14657 9676
rect 14691 9673 14703 9707
rect 14645 9667 14703 9673
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17862 9704 17868 9716
rect 17276 9676 17868 9704
rect 17276 9664 17282 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 18104 9676 18337 9704
rect 18104 9664 18110 9676
rect 18325 9673 18337 9676
rect 18371 9673 18383 9707
rect 18325 9667 18383 9673
rect 18693 9707 18751 9713
rect 18693 9673 18705 9707
rect 18739 9704 18751 9707
rect 18739 9676 19196 9704
rect 18739 9673 18751 9676
rect 18693 9667 18751 9673
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 6420 9608 7880 9636
rect 7944 9608 8769 9636
rect 6420 9596 6426 9608
rect 6454 9568 6460 9580
rect 5828 9540 6460 9568
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6816 9571 6874 9577
rect 6816 9537 6828 9571
rect 6862 9568 6874 9571
rect 7852 9568 7880 9608
rect 8757 9605 8769 9608
rect 8803 9636 8815 9639
rect 9398 9636 9404 9648
rect 8803 9608 9404 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 11698 9636 11704 9648
rect 10902 9608 11704 9636
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 14366 9636 14372 9648
rect 12728 9608 14372 9636
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 6862 9540 7604 9568
rect 7852 9540 8585 9568
rect 6862 9537 6874 9540
rect 6816 9531 6874 9537
rect 3988 9472 5948 9500
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 4062 9432 4068 9444
rect 3467 9404 4068 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 5718 9432 5724 9444
rect 4203 9404 5724 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 5626 9364 5632 9376
rect 5587 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 5920 9364 5948 9472
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6144 9472 6561 9500
rect 6144 9460 6150 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 7576 9432 7604 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8864 9500 8892 9531
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11020 9540 11805 9568
rect 11020 9528 11026 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12158 9568 12164 9580
rect 12115 9540 12164 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12728 9577 12756 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 17497 9639 17555 9645
rect 17497 9605 17509 9639
rect 17543 9605 17555 9639
rect 17880 9636 17908 9664
rect 19168 9648 19196 9676
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 21542 9704 21548 9716
rect 19852 9676 21548 9704
rect 19852 9664 19858 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 21634 9664 21640 9716
rect 21692 9704 21698 9716
rect 21692 9676 23520 9704
rect 21692 9664 21698 9676
rect 18785 9639 18843 9645
rect 17880 9608 18736 9636
rect 17497 9599 17555 9605
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13170 9568 13176 9580
rect 12943 9540 13176 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13354 9568 13360 9580
rect 13315 9540 13360 9568
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 13780 9540 16129 9568
rect 13780 9528 13786 9540
rect 16117 9537 16129 9540
rect 16163 9568 16175 9571
rect 17512 9568 17540 9599
rect 16163 9540 17540 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 7708 9472 8892 9500
rect 9401 9503 9459 9509
rect 7708 9460 7714 9472
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 10226 9500 10232 9512
rect 9723 9472 10232 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 8389 9435 8447 9441
rect 8389 9432 8401 9435
rect 7576 9404 8401 9432
rect 8389 9401 8401 9404
rect 8435 9401 8447 9435
rect 8389 9395 8447 9401
rect 9416 9376 9444 9463
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11606 9500 11612 9512
rect 11195 9472 11612 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11606 9460 11612 9472
rect 11664 9500 11670 9512
rect 15838 9500 15844 9512
rect 11664 9472 12112 9500
rect 15799 9472 15844 9500
rect 11664 9460 11670 9472
rect 7190 9364 7196 9376
rect 5920 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 9398 9364 9404 9376
rect 9311 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9364 9462 9376
rect 11054 9364 11060 9376
rect 9456 9336 11060 9364
rect 9456 9324 9462 9336
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11974 9364 11980 9376
rect 11935 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12084 9364 12112 9472
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 17512 9500 17540 9540
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17828 9540 17877 9568
rect 17828 9528 17834 9540
rect 17865 9537 17877 9540
rect 17911 9568 17923 9571
rect 18598 9568 18604 9580
rect 17911 9540 18604 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18708 9568 18736 9608
rect 18785 9605 18797 9639
rect 18831 9636 18843 9639
rect 19058 9636 19064 9648
rect 18831 9608 19064 9636
rect 18831 9605 18843 9608
rect 18785 9599 18843 9605
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 19150 9596 19156 9648
rect 19208 9596 19214 9648
rect 21177 9639 21235 9645
rect 21177 9605 21189 9639
rect 21223 9636 21235 9639
rect 22646 9636 22652 9648
rect 21223 9608 22652 9636
rect 21223 9605 21235 9608
rect 21177 9599 21235 9605
rect 22646 9596 22652 9608
rect 22704 9596 22710 9648
rect 23492 9645 23520 9676
rect 24670 9664 24676 9716
rect 24728 9664 24734 9716
rect 25038 9664 25044 9716
rect 25096 9704 25102 9716
rect 25866 9704 25872 9716
rect 25096 9676 25872 9704
rect 25096 9664 25102 9676
rect 25866 9664 25872 9676
rect 25924 9704 25930 9716
rect 26053 9707 26111 9713
rect 26053 9704 26065 9707
rect 25924 9676 26065 9704
rect 25924 9664 25930 9676
rect 26053 9673 26065 9676
rect 26099 9673 26111 9707
rect 26053 9667 26111 9673
rect 23477 9639 23535 9645
rect 23477 9605 23489 9639
rect 23523 9636 23535 9639
rect 24118 9636 24124 9648
rect 23523 9608 24124 9636
rect 23523 9605 23535 9608
rect 23477 9599 23535 9605
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 24688 9636 24716 9664
rect 24412 9608 24716 9636
rect 18708 9540 18920 9568
rect 18892 9509 18920 9540
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 22189 9571 22247 9577
rect 19024 9540 20102 9568
rect 19024 9528 19030 9540
rect 22189 9537 22201 9571
rect 22235 9568 22247 9571
rect 22554 9568 22560 9580
rect 22235 9540 22560 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 22922 9568 22928 9580
rect 22756 9540 22928 9568
rect 18877 9503 18935 9509
rect 17512 9472 18828 9500
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 15010 9432 15016 9444
rect 12851 9404 15016 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 15933 9435 15991 9441
rect 15933 9401 15945 9435
rect 15979 9432 15991 9435
rect 18800 9432 18828 9472
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21082 9500 21088 9512
rect 19751 9472 21088 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21453 9503 21511 9509
rect 21453 9469 21465 9503
rect 21499 9500 21511 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21499 9472 22109 9500
rect 21499 9469 21511 9472
rect 21453 9463 21511 9469
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22278 9500 22284 9512
rect 22239 9472 22284 9500
rect 22097 9463 22155 9469
rect 19886 9432 19892 9444
rect 15979 9404 18736 9432
rect 18800 9404 19892 9432
rect 15979 9401 15991 9404
rect 15933 9395 15991 9401
rect 13170 9364 13176 9376
rect 12084 9336 13176 9364
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 16301 9367 16359 9373
rect 16301 9333 16313 9367
rect 16347 9364 16359 9367
rect 16390 9364 16396 9376
rect 16347 9336 16396 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 18138 9364 18144 9376
rect 17543 9336 18144 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18708 9364 18736 9404
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 22112 9432 22140 9463
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 22373 9503 22431 9509
rect 22373 9469 22385 9503
rect 22419 9500 22431 9503
rect 22756 9500 22784 9540
rect 22922 9528 22928 9540
rect 22980 9528 22986 9580
rect 23106 9568 23112 9580
rect 23067 9540 23112 9568
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9568 23443 9571
rect 23569 9571 23627 9577
rect 23431 9540 23520 9568
rect 23431 9537 23443 9540
rect 23385 9531 23443 9537
rect 22419 9472 22784 9500
rect 22419 9469 22431 9472
rect 22373 9463 22431 9469
rect 23216 9444 23244 9531
rect 23492 9512 23520 9540
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 24026 9568 24032 9580
rect 23615 9540 24032 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 23474 9460 23480 9512
rect 23532 9460 23538 9512
rect 22557 9435 22615 9441
rect 22112 9404 22232 9432
rect 22204 9376 22232 9404
rect 22557 9401 22569 9435
rect 22603 9432 22615 9435
rect 22738 9432 22744 9444
rect 22603 9404 22744 9432
rect 22603 9401 22615 9404
rect 22557 9395 22615 9401
rect 22738 9392 22744 9404
rect 22796 9392 22802 9444
rect 22830 9392 22836 9444
rect 22888 9392 22894 9444
rect 23198 9392 23204 9444
rect 23256 9392 23262 9444
rect 23584 9432 23612 9531
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24412 9577 24440 9608
rect 24397 9571 24455 9577
rect 24397 9537 24409 9571
rect 24443 9537 24455 9571
rect 24578 9568 24584 9580
rect 24539 9540 24584 9568
rect 24397 9531 24455 9537
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 24728 9540 24773 9568
rect 24728 9528 24734 9540
rect 25130 9528 25136 9580
rect 25188 9568 25194 9580
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 25188 9540 25421 9568
rect 25188 9528 25194 9540
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 23934 9460 23940 9512
rect 23992 9500 23998 9512
rect 24762 9500 24768 9512
rect 23992 9472 24768 9500
rect 23992 9460 23998 9472
rect 24762 9460 24768 9472
rect 24820 9500 24826 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 24820 9472 25237 9500
rect 24820 9460 24826 9472
rect 25225 9469 25237 9472
rect 25271 9469 25283 9503
rect 25225 9463 25283 9469
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 26234 9500 26240 9512
rect 25639 9472 26240 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 23400 9404 23612 9432
rect 20070 9364 20076 9376
rect 18708 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21818 9364 21824 9376
rect 21140 9336 21824 9364
rect 21140 9324 21146 9336
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 22186 9324 22192 9376
rect 22244 9324 22250 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 22848 9364 22876 9392
rect 23400 9364 23428 9404
rect 24118 9392 24124 9444
rect 24176 9432 24182 9444
rect 24489 9435 24547 9441
rect 24176 9404 24440 9432
rect 24176 9392 24182 9404
rect 22704 9336 23428 9364
rect 22704 9324 22710 9336
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23753 9367 23811 9373
rect 23753 9364 23765 9367
rect 23532 9336 23765 9364
rect 23532 9324 23538 9336
rect 23753 9333 23765 9336
rect 23799 9333 23811 9367
rect 23753 9327 23811 9333
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 24213 9367 24271 9373
rect 24213 9364 24225 9367
rect 23900 9336 24225 9364
rect 23900 9324 23906 9336
rect 24213 9333 24225 9336
rect 24259 9333 24271 9367
rect 24412 9364 24440 9404
rect 24489 9401 24501 9435
rect 24535 9432 24547 9435
rect 24946 9432 24952 9444
rect 24535 9404 24952 9432
rect 24535 9401 24547 9404
rect 24489 9395 24547 9401
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 25608 9364 25636 9463
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 24412 9336 25636 9364
rect 24213 9327 24271 9333
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2924 9132 2973 9160
rect 2924 9120 2930 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 4890 9160 4896 9172
rect 4851 9132 4896 9160
rect 2961 9123 3019 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 7006 9160 7012 9172
rect 5316 9132 7012 9160
rect 5316 9120 5322 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7340 9132 7481 9160
rect 7340 9120 7346 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 10318 9160 10324 9172
rect 7708 9132 10324 9160
rect 7708 9120 7714 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 12805 9163 12863 9169
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 12986 9160 12992 9172
rect 12851 9132 12992 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 15838 9160 15844 9172
rect 13587 9132 15844 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 15838 9120 15844 9132
rect 15896 9160 15902 9172
rect 18874 9160 18880 9172
rect 15896 9132 18880 9160
rect 15896 9120 15902 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 20898 9160 20904 9172
rect 19208 9132 20904 9160
rect 19208 9120 19214 9132
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 21453 9163 21511 9169
rect 21453 9129 21465 9163
rect 21499 9160 21511 9163
rect 22278 9160 22284 9172
rect 21499 9132 22284 9160
rect 21499 9129 21511 9132
rect 21453 9123 21511 9129
rect 22278 9120 22284 9132
rect 22336 9160 22342 9172
rect 22738 9160 22744 9172
rect 22336 9132 22744 9160
rect 22336 9120 22342 9132
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 24670 9160 24676 9172
rect 23256 9132 24676 9160
rect 23256 9120 23262 9132
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 25590 9120 25596 9172
rect 25648 9160 25654 9172
rect 25685 9163 25743 9169
rect 25685 9160 25697 9163
rect 25648 9132 25697 9160
rect 25648 9120 25654 9132
rect 25685 9129 25697 9132
rect 25731 9129 25743 9163
rect 25685 9123 25743 9129
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 3970 9092 3976 9104
rect 1903 9064 3976 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 5442 9092 5448 9104
rect 4448 9064 5448 9092
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 4246 9024 4252 9036
rect 3016 8996 4252 9024
rect 3016 8984 3022 8996
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 3436 8965 3464 8996
rect 4246 8984 4252 8996
rect 4304 9024 4310 9036
rect 4448 9024 4476 9064
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 7024 9092 7052 9120
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 7024 9064 10149 9092
rect 10137 9061 10149 9064
rect 10183 9061 10195 9095
rect 10137 9055 10195 9061
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 18782 9092 18788 9104
rect 18196 9064 18788 9092
rect 18196 9052 18202 9064
rect 18782 9052 18788 9064
rect 18840 9092 18846 9104
rect 19242 9092 19248 9104
rect 18840 9064 19248 9092
rect 18840 9052 18846 9064
rect 19242 9052 19248 9064
rect 19300 9092 19306 9104
rect 21637 9095 21695 9101
rect 19300 9064 20852 9092
rect 19300 9052 19306 9064
rect 4304 8996 4476 9024
rect 4304 8984 4310 8996
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 2682 8888 2688 8900
rect 2004 8860 2688 8888
rect 2004 8848 2010 8860
rect 2682 8848 2688 8860
rect 2740 8888 2746 8900
rect 3160 8888 3188 8919
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3752 8928 3985 8956
rect 3752 8916 3758 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 4154 8956 4160 8968
rect 4115 8928 4160 8956
rect 3973 8919 4031 8925
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4448 8965 4476 8996
rect 4798 8984 4804 9036
rect 4856 9024 4862 9036
rect 4856 8996 6224 9024
rect 4856 8984 4862 8996
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 2740 8860 3188 8888
rect 3252 8860 4353 8888
rect 2740 8848 2746 8860
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 3252 8820 3280 8860
rect 4341 8857 4353 8860
rect 4387 8857 4399 8891
rect 4341 8851 4399 8857
rect 2464 8792 3280 8820
rect 3329 8823 3387 8829
rect 2464 8780 2470 8792
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 3510 8820 3516 8832
rect 3375 8792 3516 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 4816 8820 4844 8984
rect 5092 8965 5120 8996
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 5224 8928 5365 8956
rect 5224 8916 5230 8928
rect 5353 8925 5365 8928
rect 5399 8956 5411 8959
rect 5810 8956 5816 8968
rect 5399 8928 5816 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6196 8956 6224 8996
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 7156 8996 8217 9024
rect 7156 8984 7162 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 8570 9024 8576 9036
rect 8435 8996 8576 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 10686 9024 10692 9036
rect 10244 8996 10692 9024
rect 6356 8959 6414 8965
rect 6196 8928 6316 8956
rect 5261 8891 5319 8897
rect 5261 8857 5273 8891
rect 5307 8888 5319 8891
rect 6178 8888 6184 8900
rect 5307 8860 6184 8888
rect 5307 8857 5319 8860
rect 5261 8851 5319 8857
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 6288 8888 6316 8928
rect 6356 8925 6368 8959
rect 6402 8952 6414 8959
rect 6638 8956 6644 8968
rect 6472 8952 6644 8956
rect 6402 8928 6644 8952
rect 6402 8925 6500 8928
rect 6356 8924 6500 8925
rect 6356 8919 6414 8924
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7616 8928 8125 8956
rect 7616 8916 7622 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8588 8956 8616 8984
rect 8754 8956 8760 8968
rect 8588 8928 8760 8956
rect 8297 8919 8355 8925
rect 6288 8860 6776 8888
rect 3660 8792 4844 8820
rect 3660 8780 3666 8792
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 6638 8820 6644 8832
rect 5776 8792 6644 8820
rect 5776 8780 5782 8792
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 6748 8820 6776 8860
rect 7466 8848 7472 8900
rect 7524 8888 7530 8900
rect 8312 8888 8340 8919
rect 8754 8916 8760 8928
rect 8812 8956 8818 8968
rect 10244 8965 10272 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11054 9024 11060 9036
rect 11015 8996 11060 9024
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 13596 8996 14565 9024
rect 13596 8984 13602 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 17037 9027 17095 9033
rect 17037 9024 17049 9027
rect 15804 8996 17049 9024
rect 15804 8984 15810 8996
rect 17037 8993 17049 8996
rect 17083 8993 17095 9027
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17037 8987 17095 8993
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 17644 8996 18061 9024
rect 17644 8984 17650 8996
rect 18049 8993 18061 8996
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8812 8928 9229 8956
rect 8812 8916 8818 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10870 8956 10876 8968
rect 10459 8928 10876 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8956 20223 8959
rect 20254 8956 20260 8968
rect 20211 8928 20260 8956
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 20824 8965 20852 9064
rect 21637 9061 21649 9095
rect 21683 9092 21695 9095
rect 21726 9092 21732 9104
rect 21683 9064 21732 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 22554 9092 22560 9104
rect 21876 9064 22560 9092
rect 21876 9052 21882 9064
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 23382 9052 23388 9104
rect 23440 9092 23446 9104
rect 23440 9064 23704 9092
rect 23440 9052 23446 9064
rect 21450 8984 21456 9036
rect 21508 9024 21514 9036
rect 22189 9027 22247 9033
rect 22189 9024 22201 9027
rect 21508 8996 22201 9024
rect 21508 8984 21514 8996
rect 22189 8993 22201 8996
rect 22235 8993 22247 9027
rect 22189 8987 22247 8993
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 7524 8860 8340 8888
rect 7524 8848 7530 8860
rect 11238 8848 11244 8900
rect 11296 8888 11302 8900
rect 11333 8891 11391 8897
rect 11333 8888 11345 8891
rect 11296 8860 11345 8888
rect 11296 8848 11302 8860
rect 11333 8857 11345 8860
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 11974 8848 11980 8900
rect 12032 8848 12038 8900
rect 13722 8888 13728 8900
rect 12605 8860 13492 8888
rect 13683 8860 13728 8888
rect 7650 8820 7656 8832
rect 6748 8792 7656 8820
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7800 8792 7941 8820
rect 7800 8780 7806 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 9180 8792 9321 8820
rect 9180 8780 9186 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9309 8783 9367 8789
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 12605 8820 12633 8860
rect 10652 8792 12633 8820
rect 10652 8780 10658 8792
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 12952 8792 13369 8820
rect 12952 8780 12958 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 13464 8820 13492 8860
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 15010 8848 15016 8900
rect 15068 8848 15074 8900
rect 15930 8848 15936 8900
rect 15988 8888 15994 8900
rect 15988 8860 17080 8888
rect 15988 8848 15994 8860
rect 13525 8823 13583 8829
rect 13525 8820 13537 8823
rect 13464 8792 13537 8820
rect 13357 8783 13415 8789
rect 13525 8789 13537 8792
rect 13571 8820 13583 8823
rect 15378 8820 15384 8832
rect 13571 8792 15384 8820
rect 13571 8789 13583 8792
rect 13525 8783 13583 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15528 8792 16037 8820
rect 15528 8780 15534 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 17052 8820 17080 8860
rect 17126 8848 17132 8900
rect 17184 8888 17190 8900
rect 17184 8860 19748 8888
rect 17184 8848 17190 8860
rect 19334 8820 19340 8832
rect 17052 8792 19340 8820
rect 16025 8783 16083 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19521 8823 19579 8829
rect 19521 8789 19533 8823
rect 19567 8820 19579 8823
rect 19610 8820 19616 8832
rect 19567 8792 19616 8820
rect 19567 8789 19579 8792
rect 19521 8783 19579 8789
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 19720 8820 19748 8860
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 20364 8888 20392 8919
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 23382 8956 23388 8968
rect 22152 8928 22197 8956
rect 23343 8928 23388 8956
rect 22152 8916 22158 8928
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 23474 8916 23480 8968
rect 23532 8956 23538 8968
rect 23676 8956 23704 9064
rect 24762 9052 24768 9104
rect 24820 9052 24826 9104
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 24026 8984 24032 9036
rect 24084 9024 24090 9036
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24084 8996 24685 9024
rect 24084 8984 24090 8996
rect 24673 8993 24685 8996
rect 24719 8993 24731 9027
rect 24780 9024 24808 9052
rect 24780 8996 25636 9024
rect 24673 8987 24731 8993
rect 25608 8965 25636 8996
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 23532 8928 23577 8956
rect 23676 8928 24777 8956
rect 23532 8916 23538 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25777 8919 25835 8925
rect 20036 8860 20392 8888
rect 20036 8848 20042 8860
rect 21082 8848 21088 8900
rect 21140 8888 21146 8900
rect 21269 8891 21327 8897
rect 21269 8888 21281 8891
rect 21140 8860 21281 8888
rect 21140 8848 21146 8860
rect 21269 8857 21281 8860
rect 21315 8857 21327 8891
rect 21269 8851 21327 8857
rect 21358 8848 21364 8900
rect 21416 8888 21422 8900
rect 21469 8891 21527 8897
rect 21469 8888 21481 8891
rect 21416 8860 21481 8888
rect 21416 8848 21422 8860
rect 21469 8857 21481 8860
rect 21515 8857 21527 8891
rect 21469 8851 21527 8857
rect 23753 8891 23811 8897
rect 23753 8857 23765 8891
rect 23799 8888 23811 8891
rect 24854 8888 24860 8900
rect 23799 8860 24860 8888
rect 23799 8857 23811 8860
rect 23753 8851 23811 8857
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 22646 8820 22652 8832
rect 19720 8792 22652 8820
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 23198 8820 23204 8832
rect 23159 8792 23204 8820
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 25130 8820 25136 8832
rect 25043 8792 25136 8820
rect 25130 8780 25136 8792
rect 25188 8820 25194 8832
rect 25792 8820 25820 8919
rect 25188 8792 25820 8820
rect 25188 8780 25194 8792
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 1728 8588 4077 8616
rect 1728 8576 1734 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 5258 8616 5264 8628
rect 4295 8588 5264 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5534 8616 5540 8628
rect 5495 8588 5540 8616
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5902 8616 5908 8628
rect 5863 8588 5908 8616
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 6638 8616 6644 8628
rect 6599 8588 6644 8616
rect 6638 8576 6644 8588
rect 6696 8616 6702 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 6696 8588 7757 8616
rect 6696 8576 6702 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 12894 8616 12900 8628
rect 7745 8579 7803 8585
rect 8772 8588 12900 8616
rect 1946 8548 1952 8560
rect 1907 8520 1952 8548
rect 1946 8508 1952 8520
rect 2004 8508 2010 8560
rect 3050 8548 3056 8560
rect 3011 8520 3056 8548
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 3418 8548 3424 8560
rect 3379 8520 3424 8548
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 5442 8548 5448 8560
rect 4479 8520 5448 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 5442 8508 5448 8520
rect 5500 8548 5506 8560
rect 6012 8548 6040 8576
rect 5500 8520 6040 8548
rect 5500 8508 5506 8520
rect 2958 8480 2964 8492
rect 2919 8452 2964 8480
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3602 8480 3608 8492
rect 3283 8452 3608 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5776 8452 5821 8480
rect 5776 8440 5782 8452
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5960 8452 6009 8480
rect 5960 8440 5966 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7098 8480 7104 8492
rect 6871 8452 7104 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 6564 8412 6592 8443
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 8772 8489 8800 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 14642 8616 14648 8628
rect 13832 8588 14648 8616
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 12329 8551 12387 8557
rect 9732 8520 10166 8548
rect 9732 8508 9738 8520
rect 12329 8517 12341 8551
rect 12375 8548 12387 8551
rect 12529 8551 12587 8557
rect 12375 8517 12388 8548
rect 12329 8511 12388 8517
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 13832 8548 13860 8588
rect 14642 8576 14648 8588
rect 14700 8616 14706 8628
rect 15930 8616 15936 8628
rect 14700 8588 15936 8616
rect 14700 8576 14706 8588
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 16080 8588 16129 8616
rect 16080 8576 16086 8588
rect 16117 8585 16129 8588
rect 16163 8585 16175 8619
rect 16117 8579 16175 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 17184 8588 17325 8616
rect 17184 8576 17190 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17770 8616 17776 8628
rect 17460 8588 17505 8616
rect 17731 8588 17776 8616
rect 17460 8576 17466 8588
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 19944 8588 20729 8616
rect 19944 8576 19950 8588
rect 12575 8520 13860 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7708 8452 7849 8480
rect 7708 8440 7714 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 8757 8443 8815 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 12360 8480 12388 8511
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 13964 8520 14749 8548
rect 13964 8508 13970 8520
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 15197 8551 15255 8557
rect 15197 8548 15209 8551
rect 15160 8520 15209 8548
rect 15160 8508 15166 8520
rect 15197 8517 15209 8520
rect 15243 8517 15255 8551
rect 15197 8511 15255 8517
rect 18601 8551 18659 8557
rect 18601 8517 18613 8551
rect 18647 8548 18659 8551
rect 18966 8548 18972 8560
rect 18647 8520 18972 8548
rect 18647 8517 18659 8520
rect 18601 8511 18659 8517
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 19058 8508 19064 8560
rect 19116 8548 19122 8560
rect 20272 8557 20300 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 22186 8616 22192 8628
rect 22147 8588 22192 8616
rect 20717 8579 20775 8585
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 24118 8616 24124 8628
rect 24079 8588 24124 8616
rect 24118 8576 24124 8588
rect 24176 8616 24182 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 24176 8588 25697 8616
rect 24176 8576 24182 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 20041 8551 20099 8557
rect 20041 8548 20053 8551
rect 19116 8520 20053 8548
rect 19116 8508 19122 8520
rect 20041 8517 20053 8520
rect 20087 8548 20099 8551
rect 20257 8551 20315 8557
rect 20087 8520 20208 8548
rect 20087 8517 20099 8520
rect 20041 8511 20099 8517
rect 15381 8483 15439 8489
rect 10980 8452 12434 8480
rect 7558 8412 7564 8424
rect 6564 8384 7564 8412
rect 2498 8344 2504 8356
rect 2411 8316 2504 8344
rect 2498 8304 2504 8316
rect 2556 8344 2562 8356
rect 4985 8347 5043 8353
rect 2556 8316 4292 8344
rect 2556 8304 2562 8316
rect 4264 8285 4292 8316
rect 4985 8313 4997 8347
rect 5031 8344 5043 8347
rect 6564 8344 6592 8384
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 10980 8412 11008 8452
rect 11146 8412 11152 8424
rect 8352 8384 11008 8412
rect 11107 8384 11152 8412
rect 8352 8372 8358 8384
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 12406 8412 12434 8452
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15470 8480 15476 8492
rect 15427 8452 15476 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16301 8483 16359 8489
rect 15611 8452 15792 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 13262 8412 13268 8424
rect 12406 8384 13268 8412
rect 13262 8372 13268 8384
rect 13320 8412 13326 8424
rect 15654 8412 15660 8424
rect 13320 8384 15660 8412
rect 13320 8372 13326 8384
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15764 8412 15792 8452
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 18046 8480 18052 8492
rect 16347 8452 18052 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18156 8452 18245 8480
rect 16574 8412 16580 8424
rect 15764 8384 16580 8412
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 17218 8412 17224 8424
rect 17179 8384 17224 8412
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 5031 8316 6592 8344
rect 8205 8347 8263 8353
rect 5031 8313 5043 8316
rect 4985 8307 5043 8313
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 9306 8344 9312 8356
rect 8251 8316 9312 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9398 8304 9404 8356
rect 9456 8304 9462 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 10744 8316 12173 8344
rect 10744 8304 10750 8316
rect 12161 8313 12173 8316
rect 12207 8313 12219 8347
rect 13446 8344 13452 8356
rect 13359 8316 13452 8344
rect 12161 8307 12219 8313
rect 13446 8304 13452 8316
rect 13504 8344 13510 8356
rect 18156 8344 18184 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18380 8452 18429 8480
rect 18380 8440 18386 8452
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 18417 8443 18475 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19426 8480 19432 8492
rect 19387 8452 19432 8480
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19058 8412 19064 8424
rect 19019 8384 19064 8412
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 20180 8412 20208 8520
rect 20257 8517 20269 8551
rect 20303 8517 20315 8551
rect 20257 8511 20315 8517
rect 23008 8551 23066 8557
rect 23008 8517 23020 8551
rect 23054 8548 23066 8551
rect 23198 8548 23204 8560
rect 23054 8520 23204 8548
rect 23054 8517 23066 8520
rect 23008 8511 23066 8517
rect 23198 8508 23204 8520
rect 23256 8508 23262 8560
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20680 8452 20913 8480
rect 20680 8440 20686 8452
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21174 8480 21180 8492
rect 21131 8452 21180 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21692 8452 22017 8480
rect 21692 8440 21698 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8480 22799 8483
rect 22830 8480 22836 8492
rect 22787 8452 22836 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25041 8483 25099 8489
rect 25041 8480 25053 8483
rect 24820 8452 25053 8480
rect 24820 8440 24826 8452
rect 25041 8449 25053 8452
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 20714 8412 20720 8424
rect 20180 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 24673 8415 24731 8421
rect 24673 8412 24685 8415
rect 24636 8384 24685 8412
rect 24636 8372 24642 8384
rect 24673 8381 24685 8384
rect 24719 8381 24731 8415
rect 25130 8412 25136 8424
rect 25091 8384 25136 8412
rect 24673 8375 24731 8381
rect 25130 8372 25136 8384
rect 25188 8372 25194 8424
rect 13504 8316 18184 8344
rect 13504 8304 13510 8316
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 21174 8344 21180 8356
rect 19392 8316 21180 8344
rect 19392 8304 19398 8316
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4798 8276 4804 8288
rect 4295 8248 4804 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4798 8236 4804 8248
rect 4856 8276 4862 8288
rect 5534 8276 5540 8288
rect 4856 8248 5540 8276
rect 4856 8236 4862 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 7009 8279 7067 8285
rect 7009 8245 7021 8279
rect 7055 8276 7067 8279
rect 7282 8276 7288 8288
rect 7055 8248 7288 8276
rect 7055 8245 7067 8248
rect 7009 8239 7067 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9416 8276 9444 8304
rect 8987 8248 9444 8276
rect 9664 8279 9722 8285
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9664 8245 9676 8279
rect 9710 8276 9722 8279
rect 9858 8276 9864 8288
rect 9710 8248 9864 8276
rect 9710 8245 9722 8248
rect 9664 8239 9722 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 12345 8279 12403 8285
rect 12345 8245 12357 8279
rect 12391 8276 12403 8279
rect 16850 8276 16856 8288
rect 12391 8248 16856 8276
rect 12391 8245 12403 8248
rect 12345 8239 12403 8245
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17126 8236 17132 8288
rect 17184 8276 17190 8288
rect 19150 8276 19156 8288
rect 17184 8248 19156 8276
rect 17184 8236 17190 8248
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 19886 8276 19892 8288
rect 19847 8248 19892 8276
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 20070 8236 20076 8288
rect 20128 8276 20134 8288
rect 21450 8276 21456 8288
rect 20128 8248 21456 8276
rect 20128 8236 20134 8248
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 2958 8072 2964 8084
rect 2915 8044 2964 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3326 8032 3332 8084
rect 3384 8072 3390 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3384 8044 3985 8072
rect 3384 8032 3390 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6144 8044 6561 8072
rect 6144 8032 6150 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 7432 8044 9321 8072
rect 7432 8032 7438 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 10134 8072 10140 8084
rect 10095 8044 10140 8072
rect 9309 8035 9367 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10778 8072 10784 8084
rect 10739 8044 10784 8072
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 11238 8072 11244 8084
rect 10888 8044 11244 8072
rect 2041 8007 2099 8013
rect 2041 7973 2053 8007
rect 2087 8004 2099 8007
rect 4338 8004 4344 8016
rect 2087 7976 4344 8004
rect 2087 7973 2099 7976
rect 2041 7967 2099 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 7248 7976 9137 8004
rect 7248 7964 7254 7976
rect 9125 7973 9137 7976
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10888 8004 10916 8044
rect 11238 8032 11244 8044
rect 11296 8072 11302 8084
rect 12250 8072 12256 8084
rect 11296 8044 12256 8072
rect 11296 8032 11302 8044
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 18230 8072 18236 8084
rect 14700 8044 18236 8072
rect 14700 8032 14706 8044
rect 10100 7976 10916 8004
rect 12713 8007 12771 8013
rect 10100 7964 10106 7976
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 12894 8004 12900 8016
rect 12759 7976 12900 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 13630 7964 13636 8016
rect 13688 8004 13694 8016
rect 17126 8004 17132 8016
rect 13688 7976 17132 8004
rect 13688 7964 13694 7976
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 17954 8004 17960 8016
rect 17880 7976 17960 8004
rect 3418 7936 3424 7948
rect 3379 7908 3424 7936
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 5718 7936 5724 7948
rect 4172 7908 5724 7936
rect 4172 7877 4200 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 10594 7936 10600 7948
rect 8312 7908 10600 7936
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4304 7840 4445 7868
rect 4304 7828 4310 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7466 7868 7472 7880
rect 7248 7840 7472 7868
rect 7248 7828 7254 7840
rect 7466 7828 7472 7840
rect 7524 7868 7530 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7524 7840 7849 7868
rect 7524 7828 7530 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4341 7803 4399 7809
rect 4341 7800 4353 7803
rect 4120 7772 4353 7800
rect 4120 7760 4126 7772
rect 4341 7769 4353 7772
rect 4387 7769 4399 7803
rect 4341 7763 4399 7769
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 8113 7803 8171 7809
rect 8113 7800 8125 7803
rect 4948 7772 8125 7800
rect 4948 7760 4954 7772
rect 8113 7769 8125 7772
rect 8159 7800 8171 7803
rect 8312 7800 8340 7908
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 10704 7908 11652 7936
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9180 7840 9689 7868
rect 9180 7828 9186 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9306 7800 9312 7812
rect 8159 7772 8340 7800
rect 9267 7772 9312 7800
rect 8159 7769 8171 7772
rect 8113 7763 8171 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9692 7800 9720 7831
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10704 7877 10732 7908
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 9916 7840 10701 7868
rect 9916 7828 9922 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11054 7868 11060 7880
rect 11011 7840 11060 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 10980 7800 11008 7831
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 9692 7772 11008 7800
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7732 7622 7744
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7616 7704 7941 7732
rect 7616 7692 7622 7704
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 7929 7695 7987 7701
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 9272 7704 11529 7732
rect 9272 7692 9278 7704
rect 11517 7701 11529 7704
rect 11563 7701 11575 7735
rect 11624 7732 11652 7908
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12299 7939 12357 7945
rect 12299 7936 12311 7939
rect 12032 7908 12311 7936
rect 12032 7896 12038 7908
rect 12299 7905 12311 7908
rect 12345 7905 12357 7939
rect 12618 7936 12624 7948
rect 12299 7899 12357 7905
rect 12452 7908 12624 7936
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12452 7877 12480 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13044 7908 13369 7936
rect 13044 7896 13050 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 14366 7896 14372 7948
rect 14424 7936 14430 7948
rect 14921 7939 14979 7945
rect 14921 7936 14933 7939
rect 14424 7908 14933 7936
rect 14424 7896 14430 7908
rect 14921 7905 14933 7908
rect 14967 7936 14979 7939
rect 15102 7936 15108 7948
rect 14967 7908 15108 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 12437 7871 12495 7877
rect 12216 7840 12261 7868
rect 12216 7828 12222 7840
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13188 7800 13216 7831
rect 14642 7828 14648 7880
rect 14700 7868 14706 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14700 7840 14749 7868
rect 14700 7828 14706 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7868 17463 7871
rect 17880 7868 17908 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18064 7877 18092 8044
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 18874 8072 18880 8084
rect 18835 8044 18880 8072
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 22925 8075 22983 8081
rect 19260 8044 20484 8072
rect 19260 8016 19288 8044
rect 18138 7964 18144 8016
rect 18196 8004 18202 8016
rect 19242 8004 19248 8016
rect 18196 7976 19248 8004
rect 18196 7964 18202 7976
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 19334 7964 19340 8016
rect 19392 8004 19398 8016
rect 20349 8007 20407 8013
rect 20349 8004 20361 8007
rect 19392 7976 20361 8004
rect 19392 7964 19398 7976
rect 20349 7973 20361 7976
rect 20395 7973 20407 8007
rect 20349 7967 20407 7973
rect 19426 7936 19432 7948
rect 18156 7908 19432 7936
rect 18156 7877 18184 7908
rect 19426 7896 19432 7908
rect 19484 7936 19490 7948
rect 19484 7908 19748 7936
rect 19484 7896 19490 7908
rect 17451 7840 17908 7868
rect 18049 7871 18107 7877
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18141 7831 18199 7837
rect 16666 7800 16672 7812
rect 13188 7772 13584 7800
rect 12710 7732 12716 7744
rect 11624 7704 12716 7732
rect 11517 7695 11575 7701
rect 12710 7692 12716 7704
rect 12768 7732 12774 7744
rect 13446 7732 13452 7744
rect 12768 7704 13452 7732
rect 12768 7692 12774 7704
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13556 7732 13584 7772
rect 16040 7772 16672 7800
rect 16040 7732 16068 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 16758 7760 16764 7812
rect 16816 7800 16822 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 16816 7772 17877 7800
rect 16816 7760 16822 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 13556 7704 16068 7732
rect 16117 7735 16175 7741
rect 16117 7701 16129 7735
rect 16163 7732 16175 7735
rect 18156 7732 18184 7831
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 19720 7877 19748 7908
rect 20456 7877 20484 8044
rect 22925 8041 22937 8075
rect 22971 8072 22983 8075
rect 23382 8072 23388 8084
rect 22971 8044 23388 8072
rect 22971 8041 22983 8044
rect 22925 8035 22983 8041
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 24176 8044 24593 8072
rect 24176 8032 24182 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 24581 8035 24639 8041
rect 21266 8004 21272 8016
rect 21100 7976 21272 8004
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 21100 7945 21128 7976
rect 21266 7964 21272 7976
rect 21324 8004 21330 8016
rect 23477 8007 23535 8013
rect 23477 8004 23489 8007
rect 21324 7976 23489 8004
rect 21324 7964 21330 7976
rect 23477 7973 23489 7976
rect 23523 8004 23535 8007
rect 24029 8007 24087 8013
rect 24029 8004 24041 8007
rect 23523 7976 24041 8004
rect 23523 7973 23535 7976
rect 23477 7967 23535 7973
rect 24029 7973 24041 7976
rect 24075 8004 24087 8007
rect 24210 8004 24216 8016
rect 24075 7976 24216 8004
rect 24075 7973 24087 7976
rect 24029 7967 24087 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 21085 7939 21143 7945
rect 21085 7936 21097 7939
rect 20772 7908 21097 7936
rect 20772 7896 20778 7908
rect 21085 7905 21097 7908
rect 21131 7905 21143 7939
rect 23290 7936 23296 7948
rect 21085 7899 21143 7905
rect 21284 7908 22140 7936
rect 18877 7871 18935 7877
rect 18877 7868 18889 7871
rect 18840 7840 18889 7868
rect 18840 7828 18846 7840
rect 18877 7837 18889 7840
rect 18923 7837 18935 7871
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 18877 7831 18935 7837
rect 18984 7840 19533 7868
rect 18230 7760 18236 7812
rect 18288 7800 18294 7812
rect 18984 7800 19012 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 19751 7840 20269 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 21174 7868 21180 7880
rect 21135 7840 21180 7868
rect 20441 7831 20499 7837
rect 19426 7800 19432 7812
rect 18288 7772 19012 7800
rect 19387 7772 19432 7800
rect 18288 7760 18294 7772
rect 19426 7760 19432 7772
rect 19484 7760 19490 7812
rect 20456 7800 20484 7831
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21082 7800 21088 7812
rect 20456 7772 21088 7800
rect 21082 7760 21088 7772
rect 21140 7800 21146 7812
rect 21284 7800 21312 7908
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7868 21511 7871
rect 21542 7868 21548 7880
rect 21499 7840 21548 7868
rect 21499 7837 21511 7840
rect 21453 7831 21511 7837
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 22112 7877 22140 7908
rect 22756 7908 23296 7936
rect 22756 7877 22784 7908
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 21140 7772 21312 7800
rect 21140 7760 21146 7772
rect 16163 7704 18184 7732
rect 16163 7701 16175 7704
rect 16117 7695 16175 7701
rect 20990 7692 20996 7744
rect 21048 7732 21054 7744
rect 21928 7732 21956 7831
rect 22278 7800 22284 7812
rect 22239 7772 22284 7800
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 22940 7800 22968 7831
rect 22704 7772 22968 7800
rect 22704 7760 22710 7772
rect 21048 7704 21956 7732
rect 21048 7692 21054 7704
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1820 7500 2053 7528
rect 1820 7488 1826 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 4154 7528 4160 7540
rect 3743 7500 4160 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4982 7528 4988 7540
rect 4295 7500 4988 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5445 7531 5503 7537
rect 5445 7497 5457 7531
rect 5491 7528 5503 7531
rect 6730 7528 6736 7540
rect 5491 7500 6736 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7466 7528 7472 7540
rect 7156 7500 7472 7528
rect 7156 7488 7162 7500
rect 7466 7488 7472 7500
rect 7524 7528 7530 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7524 7500 7757 7528
rect 7524 7488 7530 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 8478 7528 8484 7540
rect 8439 7500 8484 7528
rect 7745 7491 7803 7497
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 10962 7528 10968 7540
rect 9456 7500 10968 7528
rect 9456 7488 9462 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11149 7531 11207 7537
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 12618 7528 12624 7540
rect 11195 7500 12624 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 13372 7500 16313 7528
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 5905 7463 5963 7469
rect 5905 7460 5917 7463
rect 4396 7432 5917 7460
rect 4396 7420 4402 7432
rect 5905 7429 5917 7432
rect 5951 7429 5963 7463
rect 7374 7460 7380 7472
rect 7335 7432 7380 7460
rect 5905 7423 5963 7429
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 11790 7460 11796 7472
rect 8312 7432 10180 7460
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 4890 7392 4896 7404
rect 3191 7364 4896 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5626 7392 5632 7404
rect 5307 7364 5632 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 7098 7392 7104 7404
rect 6687 7364 7104 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7282 7392 7288 7404
rect 7243 7364 7288 7392
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7742 7392 7748 7404
rect 7607 7364 7748 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 8312 7401 8340 7432
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 8297 7355 8355 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9858 7392 9864 7404
rect 9355 7364 9864 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10042 7401 10048 7404
rect 10036 7392 10048 7401
rect 10003 7364 10048 7392
rect 10036 7355 10048 7364
rect 10042 7352 10048 7355
rect 10100 7352 10106 7404
rect 10152 7392 10180 7432
rect 10336 7432 11796 7460
rect 10336 7392 10364 7432
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 10152 7364 10364 7392
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 13372 7401 13400 7500
rect 16301 7497 16313 7500
rect 16347 7528 16359 7531
rect 16482 7528 16488 7540
rect 16347 7500 16488 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 17402 7528 17408 7540
rect 16908 7500 17408 7528
rect 16908 7488 16914 7500
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 19426 7528 19432 7540
rect 17512 7500 19432 7528
rect 13998 7420 14004 7472
rect 14056 7420 14062 7472
rect 17512 7460 17540 7500
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 23566 7528 23572 7540
rect 23523 7500 23572 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 19058 7460 19064 7472
rect 15502 7432 17540 7460
rect 18354 7432 19064 7460
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 22278 7460 22284 7472
rect 20746 7432 22284 7460
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11020 7364 11713 7392
rect 11020 7352 11026 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 11701 7355 11759 7361
rect 13188 7364 13369 7392
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9640 7296 9781 7324
rect 9640 7284 9646 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12216 7296 12357 7324
rect 12216 7284 12222 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12434 7284 12440 7336
rect 12492 7333 12498 7336
rect 12492 7327 12541 7333
rect 12492 7293 12495 7327
rect 12529 7293 12541 7327
rect 12492 7287 12541 7293
rect 12492 7284 12498 7287
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 12676 7296 12721 7324
rect 12676 7284 12682 7296
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7256 4859 7259
rect 9217 7259 9275 7265
rect 4847 7228 8616 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 8478 7188 8484 7200
rect 6871 7160 8484 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 8588 7188 8616 7228
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 9674 7256 9680 7268
rect 9263 7228 9680 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 12894 7256 12900 7268
rect 11624 7228 11836 7256
rect 12855 7228 12900 7256
rect 11624 7188 11652 7228
rect 8588 7160 11652 7188
rect 11808 7188 11836 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13188 7188 13216 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 14016 7392 14044 7420
rect 13587 7364 14044 7392
rect 19245 7395 19303 7401
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 19245 7361 19257 7395
rect 19291 7392 19303 7395
rect 19886 7392 19892 7404
rect 19291 7364 19892 7392
rect 19291 7361 19303 7364
rect 19245 7355 19303 7361
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22554 7392 22560 7404
rect 22235 7364 22560 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22554 7352 22560 7364
rect 22612 7352 22618 7404
rect 22738 7392 22744 7404
rect 22699 7364 22744 7392
rect 22738 7352 22744 7364
rect 22796 7352 22802 7404
rect 13998 7324 14004 7336
rect 13959 7296 14004 7324
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 14108 7296 14289 7324
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 14108 7256 14136 7296
rect 14277 7293 14289 7296
rect 14323 7324 14335 7327
rect 15286 7324 15292 7336
rect 14323 7296 15292 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 17126 7324 17132 7336
rect 17087 7296 17132 7324
rect 16853 7287 16911 7293
rect 13780 7228 14136 7256
rect 15749 7259 15807 7265
rect 13780 7216 13786 7228
rect 15749 7225 15761 7259
rect 15795 7256 15807 7259
rect 16666 7256 16672 7268
rect 15795 7228 16672 7256
rect 15795 7225 15807 7228
rect 15749 7219 15807 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 11808 7160 13216 7188
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 16868 7188 16896 7287
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 17552 7296 19717 7324
rect 17552 7284 17558 7296
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7324 21235 7327
rect 21453 7327 21511 7333
rect 21223 7296 21404 7324
rect 21223 7293 21235 7296
rect 21177 7287 21235 7293
rect 19061 7259 19119 7265
rect 19061 7256 19073 7259
rect 18156 7228 19073 7256
rect 17126 7188 17132 7200
rect 14148 7160 17132 7188
rect 14148 7148 14154 7160
rect 17126 7148 17132 7160
rect 17184 7188 17190 7200
rect 18156 7188 18184 7228
rect 19061 7225 19073 7228
rect 19107 7225 19119 7259
rect 19061 7219 19119 7225
rect 17184 7160 18184 7188
rect 18601 7191 18659 7197
rect 17184 7148 17190 7160
rect 18601 7157 18613 7191
rect 18647 7188 18659 7191
rect 18690 7188 18696 7200
rect 18647 7160 18696 7188
rect 18647 7157 18659 7160
rect 18601 7151 18659 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 19720 7188 19748 7287
rect 21376 7256 21404 7296
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 22005 7327 22063 7333
rect 22005 7324 22017 7327
rect 21499 7296 22017 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 22005 7293 22017 7296
rect 22051 7293 22063 7327
rect 22005 7287 22063 7293
rect 21542 7256 21548 7268
rect 21376 7228 21548 7256
rect 21542 7216 21548 7228
rect 21600 7256 21606 7268
rect 22833 7259 22891 7265
rect 22833 7256 22845 7259
rect 21600 7228 22845 7256
rect 21600 7216 21606 7228
rect 22833 7225 22845 7228
rect 22879 7225 22891 7259
rect 22833 7219 22891 7225
rect 22738 7188 22744 7200
rect 19720 7160 22744 7188
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7156 6956 7389 6984
rect 7156 6944 7162 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7524 6956 7573 6984
rect 7524 6944 7530 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 7800 6956 8401 6984
rect 7800 6944 7806 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 11057 6987 11115 6993
rect 9732 6956 10732 6984
rect 9732 6944 9738 6956
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 8294 6916 8300 6928
rect 4856 6888 8300 6916
rect 4856 6876 4862 6888
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2498 6848 2504 6860
rect 1995 6820 2504 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3878 6848 3884 6860
rect 3467 6820 3884 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4338 6848 4344 6860
rect 4299 6820 4344 6848
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4982 6848 4988 6860
rect 4943 6820 4988 6848
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 5868 6820 9137 6848
rect 5868 6808 5874 6820
rect 9125 6817 9137 6820
rect 9171 6848 9183 6851
rect 10704 6848 10732 6956
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11882 6984 11888 6996
rect 11103 6956 11888 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12676 6956 12909 6984
rect 12676 6944 12682 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 16574 6916 16580 6928
rect 13924 6888 14412 6916
rect 16487 6888 16580 6916
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 9171 6820 9812 6848
rect 10704 6820 11529 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 9784 6792 9812 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 13538 6848 13544 6860
rect 13499 6820 13544 6848
rect 11517 6811 11575 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6638 6780 6644 6792
rect 6135 6752 6644 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7558 6780 7564 6792
rect 6963 6752 7564 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 9582 6780 9588 6792
rect 8536 6752 9588 6780
rect 8536 6740 8542 6752
rect 9582 6740 9588 6752
rect 9640 6780 9646 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9640 6752 9689 6780
rect 9640 6740 9646 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 10686 6780 10692 6792
rect 9876 6752 10692 6780
rect 2682 6672 2688 6724
rect 2740 6712 2746 6724
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 2740 6684 5549 6712
rect 2740 6672 2746 6684
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 5537 6675 5595 6681
rect 6825 6715 6883 6721
rect 6825 6681 6837 6715
rect 6871 6712 6883 6715
rect 7374 6712 7380 6724
rect 6871 6684 7380 6712
rect 6871 6681 6883 6684
rect 6825 6675 6883 6681
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 7484 6684 7757 6712
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 3326 6644 3332 6656
rect 2547 6616 3332 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 6181 6647 6239 6653
rect 6181 6613 6193 6647
rect 6227 6644 6239 6647
rect 7190 6644 7196 6656
rect 6227 6616 7196 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 7190 6604 7196 6616
rect 7248 6644 7254 6656
rect 7484 6644 7512 6684
rect 7745 6681 7757 6684
rect 7791 6712 7803 6715
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 7791 6684 8217 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 8662 6712 8668 6724
rect 8205 6675 8263 6681
rect 8404 6684 8668 6712
rect 8404 6653 8432 6684
rect 8662 6672 8668 6684
rect 8720 6712 8726 6724
rect 9876 6712 9904 6752
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13320 6752 13461 6780
rect 13320 6740 13326 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13924 6780 13952 6888
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14148 6820 14289 6848
rect 14148 6808 14154 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14384 6848 14412 6888
rect 16574 6876 16580 6888
rect 16632 6876 16638 6928
rect 22373 6919 22431 6925
rect 22373 6885 22385 6919
rect 22419 6885 22431 6919
rect 22373 6879 22431 6885
rect 16592 6848 16620 6876
rect 17126 6848 17132 6860
rect 14384 6820 16620 6848
rect 17087 6820 17132 6848
rect 14277 6811 14335 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 22388 6848 22416 6879
rect 19444 6820 22416 6848
rect 13679 6752 13952 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 15988 6752 16497 6780
rect 15988 6740 15994 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 16850 6780 16856 6792
rect 16715 6752 16856 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 19444 6789 19472 6820
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 20073 6783 20131 6789
rect 20073 6780 20085 6783
rect 19429 6743 19487 6749
rect 19628 6752 20085 6780
rect 8720 6684 9904 6712
rect 9944 6715 10002 6721
rect 8720 6672 8726 6684
rect 9944 6681 9956 6715
rect 9990 6712 10002 6715
rect 10042 6712 10048 6724
rect 9990 6684 10048 6712
rect 9990 6681 10002 6684
rect 9944 6675 10002 6681
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 11422 6672 11428 6724
rect 11480 6712 11486 6724
rect 11762 6715 11820 6721
rect 11762 6712 11774 6715
rect 11480 6684 11774 6712
rect 11480 6672 11486 6684
rect 11762 6681 11774 6684
rect 11808 6712 11820 6715
rect 14550 6712 14556 6724
rect 11808 6684 14556 6712
rect 11808 6681 11820 6684
rect 11762 6675 11820 6681
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 16758 6712 16764 6724
rect 15778 6684 16764 6712
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 17402 6712 17408 6724
rect 17363 6684 17408 6712
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 19334 6712 19340 6724
rect 18630 6684 19340 6712
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 7248 6616 7512 6644
rect 7545 6647 7603 6653
rect 7248 6604 7254 6616
rect 7545 6613 7557 6647
rect 7591 6644 7603 6647
rect 8404 6647 8463 6653
rect 8404 6644 8417 6647
rect 7591 6616 8417 6644
rect 7591 6613 7603 6616
rect 7545 6607 7603 6613
rect 8405 6613 8417 6616
rect 8451 6613 8463 6647
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8405 6607 8463 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 16022 6644 16028 6656
rect 15983 6616 16028 6644
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 18874 6644 18880 6656
rect 18835 6616 18880 6644
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 19628 6653 19656 6752
rect 20073 6749 20085 6752
rect 20119 6749 20131 6783
rect 20438 6780 20444 6792
rect 20399 6752 20444 6780
rect 20073 6743 20131 6749
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 22554 6780 22560 6792
rect 22515 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 20806 6672 20812 6724
rect 20864 6672 20870 6724
rect 19613 6647 19671 6653
rect 19613 6613 19625 6647
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21867 6647 21925 6653
rect 21867 6644 21879 6647
rect 20772 6616 21879 6644
rect 20772 6604 20778 6616
rect 21867 6613 21879 6616
rect 21913 6613 21925 6647
rect 21867 6607 21925 6613
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 3326 6440 3332 6452
rect 3239 6412 3332 6440
rect 3326 6400 3332 6412
rect 3384 6440 3390 6452
rect 5442 6440 5448 6452
rect 3384 6412 5448 6440
rect 3384 6400 3390 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 7009 6443 7067 6449
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7742 6440 7748 6452
rect 7055 6412 7748 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 8352 6412 9229 6440
rect 8352 6400 8358 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 12434 6440 12440 6452
rect 11195 6412 12440 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 14642 6440 14648 6452
rect 12912 6412 14648 6440
rect 4338 6372 4344 6384
rect 4299 6344 4344 6372
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 8386 6332 8392 6384
rect 8444 6372 8450 6384
rect 10036 6375 10094 6381
rect 8444 6344 9996 6372
rect 8444 6332 8450 6344
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2682 6304 2688 6316
rect 2363 6276 2688 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3660 6276 3801 6304
rect 3660 6264 3666 6276
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7466 6304 7472 6316
rect 6963 6276 7472 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8662 6304 8668 6316
rect 8619 6276 8668 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9582 6304 9588 6316
rect 9364 6276 9588 6304
rect 9364 6264 9370 6276
rect 9582 6264 9588 6276
rect 9640 6304 9646 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9640 6276 9781 6304
rect 9640 6264 9646 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9968 6304 9996 6344
rect 10036 6341 10048 6375
rect 10082 6372 10094 6375
rect 11422 6372 11428 6384
rect 10082 6344 11428 6372
rect 10082 6341 10094 6344
rect 10036 6335 10094 6341
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 11698 6372 11704 6384
rect 11659 6344 11704 6372
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 12912 6372 12940 6412
rect 14642 6400 14648 6412
rect 14700 6440 14706 6452
rect 15010 6440 15016 6452
rect 14700 6412 15016 6440
rect 14700 6400 14706 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 18138 6440 18144 6452
rect 16347 6412 18144 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 19242 6440 19248 6452
rect 19203 6412 19248 6440
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 20956 6412 21281 6440
rect 20956 6400 20962 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 11900 6344 12940 6372
rect 12989 6375 13047 6381
rect 9968 6276 11008 6304
rect 9769 6267 9827 6273
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 6696 6208 8401 6236
rect 6696 6196 6702 6208
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 10980 6236 11008 6276
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11900 6313 11928 6344
rect 12989 6341 13001 6375
rect 13035 6372 13047 6375
rect 13814 6372 13820 6384
rect 13035 6344 13820 6372
rect 13035 6341 13047 6344
rect 12989 6335 13047 6341
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 16758 6372 16764 6384
rect 15764 6344 16764 6372
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11112 6276 11897 6304
rect 11112 6264 11118 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12710 6304 12716 6316
rect 12115 6276 12716 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12710 6264 12716 6276
rect 12768 6304 12774 6316
rect 14826 6304 14832 6316
rect 12768 6276 14832 6304
rect 12768 6264 12774 6276
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 10980 6208 12434 6236
rect 8389 6199 8447 6205
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 7282 6168 7288 6180
rect 4212 6140 7288 6168
rect 4212 6128 4218 6140
rect 7282 6128 7288 6140
rect 7340 6168 7346 6180
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7340 6140 7849 6168
rect 7340 6128 7346 6140
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 8757 6171 8815 6177
rect 8757 6137 8769 6171
rect 8803 6168 8815 6171
rect 12406 6168 12434 6208
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 15764 6245 15792 6344
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 16942 6332 16948 6384
rect 17000 6372 17006 6384
rect 17865 6375 17923 6381
rect 17865 6372 17877 6375
rect 17000 6344 17877 6372
rect 17000 6332 17006 6344
rect 17865 6341 17877 6344
rect 17911 6341 17923 6375
rect 18874 6372 18880 6384
rect 17865 6335 17923 6341
rect 18340 6344 18880 6372
rect 15930 6304 15936 6316
rect 15891 6276 15936 6304
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16080 6276 17049 6304
rect 16080 6264 16086 6276
rect 17037 6273 17049 6276
rect 17083 6304 17095 6307
rect 18230 6304 18236 6316
rect 17083 6276 18236 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 18340 6313 18368 6344
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 19058 6332 19064 6384
rect 19116 6372 19122 6384
rect 20438 6372 20444 6384
rect 19116 6344 20444 6372
rect 19116 6332 19122 6344
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 20806 6372 20812 6384
rect 20767 6344 20812 6372
rect 20806 6332 20812 6344
rect 20864 6332 20870 6384
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6304 18567 6307
rect 18690 6304 18696 6316
rect 18555 6276 18696 6304
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 18800 6276 19349 6304
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 14332 6208 14749 6236
rect 14332 6196 14338 6208
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 13630 6168 13636 6180
rect 8803 6140 9812 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 2866 6100 2872 6112
rect 1811 6072 2872 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 2866 6060 2872 6072
rect 2924 6100 2930 6112
rect 3602 6100 3608 6112
rect 2924 6072 3608 6100
rect 2924 6060 2930 6072
rect 3602 6060 3608 6072
rect 3660 6100 3666 6112
rect 5166 6100 5172 6112
rect 3660 6072 5172 6100
rect 3660 6060 3666 6072
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5868 6072 5917 6100
rect 5868 6060 5874 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 9784 6100 9812 6140
rect 11072 6140 11284 6168
rect 12406 6140 13636 6168
rect 11072 6100 11100 6140
rect 9784 6072 11100 6100
rect 11256 6100 11284 6140
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 14752 6168 14780 6199
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 15896 6208 15941 6236
rect 15896 6196 15902 6208
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 16724 6208 16957 6236
rect 16724 6196 16730 6208
rect 16945 6205 16957 6208
rect 16991 6205 17003 6239
rect 16945 6199 17003 6205
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 17276 6208 17509 6236
rect 17276 6196 17282 6208
rect 17497 6205 17509 6208
rect 17543 6236 17555 6239
rect 18800 6236 18828 6276
rect 19337 6273 19349 6276
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 21082 6304 21088 6316
rect 20763 6276 21088 6304
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 19058 6236 19064 6248
rect 17543 6208 18828 6236
rect 19019 6208 19064 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 19426 6236 19432 6248
rect 19300 6208 19432 6236
rect 19300 6196 19306 6208
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 20548 6236 20576 6267
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 20990 6236 20996 6248
rect 20548 6208 20996 6236
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 22186 6168 22192 6180
rect 14752 6140 18552 6168
rect 16022 6100 16028 6112
rect 11256 6072 16028 6100
rect 5905 6063 5963 6069
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6100 17463 6103
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 17451 6072 18429 6100
rect 17451 6069 17463 6072
rect 17405 6063 17463 6069
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 18524 6100 18552 6140
rect 19306 6140 22192 6168
rect 19306 6100 19334 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 19702 6100 19708 6112
rect 18524 6072 19334 6100
rect 19663 6072 19708 6100
rect 18417 6063 18475 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 14 5856 20 5908
rect 72 5896 78 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 72 5868 7849 5896
rect 72 5856 78 5868
rect 7837 5865 7849 5868
rect 7883 5896 7895 5899
rect 13354 5896 13360 5908
rect 7883 5868 13360 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14458 5896 14464 5908
rect 14415 5868 14464 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14792 5868 14933 5896
rect 14792 5856 14798 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 17865 5899 17923 5905
rect 17865 5896 17877 5899
rect 15988 5868 17877 5896
rect 15988 5856 15994 5868
rect 17865 5865 17877 5868
rect 17911 5865 17923 5899
rect 17865 5859 17923 5865
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 19058 5896 19064 5908
rect 18012 5868 19064 5896
rect 18012 5856 18018 5868
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 20717 5899 20775 5905
rect 20717 5896 20729 5899
rect 20496 5868 20729 5896
rect 20496 5856 20502 5868
rect 20717 5865 20729 5868
rect 20763 5865 20775 5899
rect 20717 5859 20775 5865
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 2777 5831 2835 5837
rect 2777 5828 2789 5831
rect 2740 5800 2789 5828
rect 2740 5788 2746 5800
rect 2777 5797 2789 5800
rect 2823 5797 2835 5831
rect 2777 5791 2835 5797
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4522 5828 4528 5840
rect 4212 5800 4528 5828
rect 4212 5788 4218 5800
rect 4522 5788 4528 5800
rect 4580 5788 4586 5840
rect 5074 5828 5080 5840
rect 5035 5800 5080 5828
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5718 5828 5724 5840
rect 5679 5800 5724 5828
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 8573 5831 8631 5837
rect 8573 5797 8585 5831
rect 8619 5828 8631 5831
rect 10873 5831 10931 5837
rect 8619 5800 9536 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2866 5760 2872 5772
rect 2363 5732 2872 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3467 5732 4077 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4246 5760 4252 5772
rect 4111 5732 4252 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 7742 5760 7748 5772
rect 6319 5732 7748 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 7742 5720 7748 5732
rect 7800 5760 7806 5772
rect 8754 5760 8760 5772
rect 7800 5732 8760 5760
rect 7800 5720 7806 5732
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 4264 5692 4292 5720
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 4264 5664 7297 5692
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8570 5692 8576 5704
rect 8435 5664 8576 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 9508 5701 9536 5800
rect 10873 5797 10885 5831
rect 10919 5797 10931 5831
rect 10873 5791 10931 5797
rect 10888 5760 10916 5791
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 19518 5828 19524 5840
rect 15896 5800 19524 5828
rect 15896 5788 15902 5800
rect 19518 5788 19524 5800
rect 19576 5788 19582 5840
rect 20070 5788 20076 5840
rect 20128 5828 20134 5840
rect 21361 5831 21419 5837
rect 21361 5828 21373 5831
rect 20128 5800 21373 5828
rect 20128 5788 20134 5800
rect 21361 5797 21373 5800
rect 21407 5797 21419 5831
rect 21361 5791 21419 5797
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 10888 5732 12541 5760
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 12894 5760 12900 5772
rect 12851 5732 12900 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 12894 5720 12900 5732
rect 12952 5760 12958 5772
rect 12952 5732 15148 5760
rect 12952 5720 12958 5732
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 9582 5692 9588 5704
rect 9539 5664 9588 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12434 5701 12440 5704
rect 12412 5695 12440 5701
rect 12308 5664 12353 5692
rect 12308 5652 12314 5664
rect 12412 5661 12424 5695
rect 12412 5655 12440 5661
rect 12434 5652 12440 5655
rect 12492 5652 12498 5704
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13354 5692 13360 5704
rect 13311 5664 13360 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 14826 5692 14832 5704
rect 14787 5664 14832 5692
rect 13449 5655 13507 5661
rect 6825 5627 6883 5633
rect 6825 5593 6837 5627
rect 6871 5624 6883 5627
rect 8294 5624 8300 5636
rect 6871 5596 8300 5624
rect 6871 5593 6883 5596
rect 6825 5587 6883 5593
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 9760 5627 9818 5633
rect 9760 5593 9772 5627
rect 9806 5624 9818 5627
rect 9858 5624 9864 5636
rect 9806 5596 9864 5624
rect 9806 5593 9818 5596
rect 9760 5587 9818 5593
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 11146 5584 11152 5636
rect 11204 5624 11210 5636
rect 11204 5596 11744 5624
rect 11204 5584 11210 5596
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 11020 5528 11621 5556
rect 11020 5516 11026 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 11716 5556 11744 5596
rect 13464 5556 13492 5655
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 15010 5692 15016 5704
rect 14971 5664 15016 5692
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15120 5692 15148 5732
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 15712 5732 18337 5760
rect 15712 5720 15718 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 19610 5760 19616 5772
rect 18472 5732 19616 5760
rect 18472 5720 18478 5732
rect 19610 5720 19616 5732
rect 19668 5760 19674 5772
rect 19978 5760 19984 5772
rect 19668 5732 19984 5760
rect 19668 5720 19674 5732
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 20162 5720 20168 5772
rect 20220 5760 20226 5772
rect 20220 5732 21588 5760
rect 20220 5720 20226 5732
rect 17954 5692 17960 5704
rect 15120 5664 17960 5692
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 18932 5664 19809 5692
rect 18932 5652 18938 5664
rect 19797 5661 19809 5664
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 21560 5701 21588 5732
rect 20717 5695 20775 5701
rect 20717 5692 20729 5695
rect 20680 5664 20729 5692
rect 20680 5652 20686 5664
rect 20717 5661 20729 5664
rect 20763 5661 20775 5695
rect 20717 5655 20775 5661
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 15657 5627 15715 5633
rect 15657 5593 15669 5627
rect 15703 5624 15715 5627
rect 16482 5624 16488 5636
rect 15703 5596 16488 5624
rect 15703 5593 15715 5596
rect 15657 5587 15715 5593
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 20990 5624 20996 5636
rect 16960 5596 20996 5624
rect 11716 5528 13492 5556
rect 11609 5519 11667 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 16960 5565 16988 5596
rect 20990 5584 20996 5596
rect 21048 5584 21054 5636
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 15528 5528 16957 5556
rect 15528 5516 15534 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 16945 5519 17003 5525
rect 19886 5516 19892 5568
rect 19944 5556 19950 5568
rect 22097 5559 22155 5565
rect 19944 5528 19989 5556
rect 19944 5516 19950 5528
rect 22097 5525 22109 5559
rect 22143 5556 22155 5559
rect 22278 5556 22284 5568
rect 22143 5528 22284 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22278 5516 22284 5528
rect 22336 5516 22342 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2372 5324 2605 5352
rect 2372 5312 2378 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4065 5355 4123 5361
rect 4065 5352 4077 5355
rect 3559 5324 4077 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4065 5321 4077 5324
rect 4111 5352 4123 5355
rect 4246 5352 4252 5364
rect 4111 5324 4252 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 2608 5284 2636 5315
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4522 5352 4528 5364
rect 4483 5324 4528 5352
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5166 5352 5172 5364
rect 5127 5324 5172 5352
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5905 5355 5963 5361
rect 5905 5352 5917 5355
rect 5500 5324 5917 5352
rect 5500 5312 5506 5324
rect 5905 5321 5917 5324
rect 5951 5321 5963 5355
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 5905 5315 5963 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 12342 5352 12348 5364
rect 10735 5324 12348 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 15565 5355 15623 5361
rect 12492 5324 15516 5352
rect 12492 5312 12498 5324
rect 5810 5284 5816 5296
rect 2608 5256 5816 5284
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 10962 5284 10968 5296
rect 8864 5256 10968 5284
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6638 5216 6644 5228
rect 5776 5188 6644 5216
rect 5776 5176 5782 5188
rect 6638 5176 6644 5188
rect 6696 5216 6702 5228
rect 8864 5225 8892 5256
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 14452 5287 14510 5293
rect 14452 5253 14464 5287
rect 14498 5284 14510 5287
rect 15286 5284 15292 5296
rect 14498 5256 15292 5284
rect 14498 5253 14510 5256
rect 14452 5247 14510 5253
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6696 5188 7021 5216
rect 6696 5176 6702 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5185 8907 5219
rect 9306 5216 9312 5228
rect 9267 5188 9312 5216
rect 8849 5179 8907 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9576 5219 9634 5225
rect 9576 5185 9588 5219
rect 9622 5216 9634 5219
rect 9858 5216 9864 5228
rect 9622 5188 9864 5216
rect 9622 5185 9634 5188
rect 9576 5179 9634 5185
rect 9858 5176 9864 5188
rect 9916 5216 9922 5228
rect 10410 5216 10416 5228
rect 9916 5188 10416 5216
rect 9916 5176 9922 5188
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13228 5188 13553 5216
rect 13228 5176 13234 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 12158 5108 12164 5160
rect 12216 5148 12222 5160
rect 12345 5151 12403 5157
rect 12345 5148 12357 5151
rect 12216 5120 12357 5148
rect 12216 5108 12222 5120
rect 12345 5117 12357 5120
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 12434 5108 12440 5160
rect 12492 5157 12498 5160
rect 12492 5151 12541 5157
rect 12492 5117 12495 5151
rect 12529 5117 12541 5151
rect 12492 5111 12541 5117
rect 12492 5108 12498 5111
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12894 5148 12900 5160
rect 12676 5120 12721 5148
rect 12855 5120 12900 5148
rect 12676 5108 12682 5120
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5117 13415 5151
rect 14182 5148 14188 5160
rect 14143 5120 14188 5148
rect 13357 5111 13415 5117
rect 7653 5083 7711 5089
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 7926 5080 7932 5092
rect 7699 5052 7932 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 7926 5040 7932 5052
rect 7984 5080 7990 5092
rect 7984 5052 8800 5080
rect 7984 5040 7990 5052
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 8536 4984 8677 5012
rect 8536 4972 8542 4984
rect 8665 4981 8677 4984
rect 8711 4981 8723 5015
rect 8772 5012 8800 5052
rect 10244 5052 11836 5080
rect 10244 5012 10272 5052
rect 8772 4984 10272 5012
rect 8665 4975 8723 4981
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 10836 4984 11713 5012
rect 10836 4972 10842 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11808 5012 11836 5052
rect 12802 5012 12808 5024
rect 11808 4984 12808 5012
rect 11701 4975 11759 4981
rect 12802 4972 12808 4984
rect 12860 5012 12866 5024
rect 13372 5012 13400 5111
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 15488 5148 15516 5324
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 17129 5355 17187 5361
rect 17129 5352 17141 5355
rect 15611 5324 17141 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 17129 5321 17141 5324
rect 17175 5321 17187 5355
rect 17129 5315 17187 5321
rect 19429 5355 19487 5361
rect 19429 5321 19441 5355
rect 19475 5352 19487 5355
rect 19886 5352 19892 5364
rect 19475 5324 19892 5352
rect 19475 5321 19487 5324
rect 19429 5315 19487 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 22278 5352 22284 5364
rect 22020 5324 22284 5352
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 17221 5287 17279 5293
rect 17221 5284 17233 5287
rect 16724 5256 17233 5284
rect 16724 5244 16730 5256
rect 17221 5253 17233 5256
rect 17267 5253 17279 5287
rect 17221 5247 17279 5253
rect 17586 5244 17592 5296
rect 17644 5284 17650 5296
rect 18294 5287 18352 5293
rect 18294 5284 18306 5287
rect 17644 5256 18306 5284
rect 17644 5244 17650 5256
rect 18294 5253 18306 5256
rect 18340 5253 18352 5287
rect 18294 5247 18352 5253
rect 18414 5244 18420 5296
rect 18472 5244 18478 5296
rect 16022 5216 16028 5228
rect 15983 5188 16028 5216
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 18432 5216 18460 5244
rect 16960 5188 18460 5216
rect 16960 5157 16988 5188
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 18748 5188 19901 5216
rect 18748 5176 18754 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 21048 5188 21097 5216
rect 21048 5176 21054 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 21634 5176 21640 5228
rect 21692 5216 21698 5228
rect 22020 5225 22048 5324
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22189 5287 22247 5293
rect 22189 5253 22201 5287
rect 22235 5284 22247 5287
rect 22462 5284 22468 5296
rect 22235 5256 22468 5284
rect 22235 5253 22247 5256
rect 22189 5247 22247 5253
rect 22462 5244 22468 5256
rect 22520 5244 22526 5296
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21692 5188 22017 5216
rect 21692 5176 21698 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5216 22431 5219
rect 23477 5219 23535 5225
rect 23477 5216 23489 5219
rect 22419 5188 23489 5216
rect 22419 5185 22431 5188
rect 22373 5179 22431 5185
rect 23477 5185 23489 5188
rect 23523 5185 23535 5219
rect 23477 5179 23535 5185
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 15488 5120 16957 5148
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 18064 5080 18092 5111
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 20165 5151 20223 5157
rect 20165 5148 20177 5151
rect 19484 5120 20177 5148
rect 19484 5108 19490 5120
rect 20165 5117 20177 5120
rect 20211 5148 20223 5151
rect 20622 5148 20628 5160
rect 20211 5120 20628 5148
rect 20211 5117 20223 5120
rect 20165 5111 20223 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 16224 5052 18092 5080
rect 16224 5024 16252 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 20993 5083 21051 5089
rect 20993 5080 21005 5083
rect 19392 5052 21005 5080
rect 19392 5040 19398 5052
rect 20993 5049 21005 5052
rect 21039 5049 21051 5083
rect 20993 5043 21051 5049
rect 12860 4984 13400 5012
rect 12860 4972 12866 4984
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 16206 5012 16212 5024
rect 14240 4984 16212 5012
rect 14240 4972 14246 4984
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17276 4984 17601 5012
rect 17276 4972 17282 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 17589 4975 17647 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 5012 20499 5015
rect 20622 5012 20628 5024
rect 20487 4984 20628 5012
rect 20487 4981 20499 4984
rect 20441 4975 20499 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 23293 5015 23351 5021
rect 23293 5012 23305 5015
rect 22336 4984 23305 5012
rect 22336 4972 22342 4984
rect 23293 4981 23305 4984
rect 23339 4981 23351 5015
rect 23293 4975 23351 4981
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 4617 4811 4675 4817
rect 4617 4777 4629 4811
rect 4663 4808 4675 4811
rect 4798 4808 4804 4820
rect 4663 4780 4804 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4948 4780 5181 4808
rect 4948 4768 4954 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 6638 4808 6644 4820
rect 6599 4780 6644 4808
rect 5169 4771 5227 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 12618 4808 12624 4820
rect 10827 4780 12624 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 12912 4780 16160 4808
rect 4816 4740 4844 4768
rect 6089 4743 6147 4749
rect 6089 4740 6101 4743
rect 4816 4712 6101 4740
rect 6089 4709 6101 4712
rect 6135 4709 6147 4743
rect 6089 4703 6147 4709
rect 10410 4700 10416 4752
rect 10468 4740 10474 4752
rect 12912 4740 12940 4780
rect 10468 4712 12940 4740
rect 10468 4700 10474 4712
rect 12986 4700 12992 4752
rect 13044 4740 13050 4752
rect 13044 4712 13089 4740
rect 13044 4700 13050 4712
rect 10502 4632 10508 4684
rect 10560 4672 10566 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 10560 4644 11253 4672
rect 10560 4632 10566 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4672 12495 4675
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 12483 4644 13553 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 13541 4641 13553 4644
rect 13587 4672 13599 4675
rect 14642 4672 14648 4684
rect 13587 4644 14648 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9490 4604 9496 4616
rect 9447 4576 9496 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 12986 4604 12992 4616
rect 9600 4576 12992 4604
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 9600 4536 9628 4576
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14734 4604 14740 4616
rect 14323 4576 14740 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 16132 4604 16160 4780
rect 18877 4743 18935 4749
rect 18877 4709 18889 4743
rect 18923 4740 18935 4743
rect 19521 4743 19579 4749
rect 19521 4740 19533 4743
rect 18923 4712 19533 4740
rect 18923 4709 18935 4712
rect 18877 4703 18935 4709
rect 19521 4709 19533 4712
rect 19567 4709 19579 4743
rect 19521 4703 19579 4709
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 16264 4644 17509 4672
rect 16264 4632 16270 4644
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17497 4635 17555 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19978 4672 19984 4684
rect 19751 4644 19984 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 17034 4604 17040 4616
rect 16132 4576 17040 4604
rect 17034 4564 17040 4576
rect 17092 4604 17098 4616
rect 17753 4607 17811 4613
rect 17753 4604 17765 4607
rect 17092 4576 17765 4604
rect 17092 4564 17098 4576
rect 17753 4573 17765 4576
rect 17799 4573 17811 4607
rect 19426 4604 19432 4616
rect 19387 4576 19432 4604
rect 17753 4567 17811 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 22244 4576 22845 4604
rect 22244 4564 22250 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 22922 4564 22928 4616
rect 22980 4604 22986 4616
rect 23477 4607 23535 4613
rect 23477 4604 23489 4607
rect 22980 4576 23489 4604
rect 22980 4564 22986 4576
rect 23477 4573 23489 4576
rect 23523 4573 23535 4607
rect 23477 4567 23535 4573
rect 8352 4508 9628 4536
rect 9668 4539 9726 4545
rect 8352 4496 8358 4508
rect 9668 4505 9680 4539
rect 9714 4536 9726 4539
rect 9858 4536 9864 4548
rect 9714 4508 9864 4536
rect 9714 4505 9726 4508
rect 9668 4499 9726 4505
rect 9858 4496 9864 4508
rect 9916 4536 9922 4548
rect 10226 4536 10232 4548
rect 9916 4508 10232 4536
rect 9916 4496 9922 4508
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 11204 4508 13461 4536
rect 11204 4496 11210 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13449 4499 13507 4505
rect 15197 4539 15255 4545
rect 15197 4505 15209 4539
rect 15243 4505 15255 4539
rect 15197 4499 15255 4505
rect 19705 4539 19763 4545
rect 19705 4505 19717 4539
rect 19751 4536 19763 4539
rect 20530 4536 20536 4548
rect 19751 4508 20536 4536
rect 19751 4505 19763 4508
rect 19705 4499 19763 4505
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4468 8539 4471
rect 10410 4468 10416 4480
rect 8527 4440 10416 4468
rect 8527 4437 8539 4440
rect 8481 4431 8539 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11330 4428 11336 4480
rect 11388 4468 11394 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 11388 4440 11805 4468
rect 11388 4428 11394 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 11940 4440 12173 4468
rect 11940 4428 11946 4440
rect 12161 4437 12173 4440
rect 12207 4437 12219 4471
rect 12161 4431 12219 4437
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 13354 4468 13360 4480
rect 12308 4440 12353 4468
rect 13315 4440 13360 4468
rect 12308 4428 12314 4440
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 14461 4471 14519 4477
rect 14461 4437 14473 4471
rect 14507 4468 14519 4471
rect 15212 4468 15240 4499
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 22588 4539 22646 4545
rect 22588 4505 22600 4539
rect 22634 4536 22646 4539
rect 24486 4536 24492 4548
rect 22634 4508 24492 4536
rect 22634 4505 22646 4508
rect 22588 4499 22646 4505
rect 24486 4496 24492 4508
rect 24544 4496 24550 4548
rect 16482 4468 16488 4480
rect 14507 4440 15240 4468
rect 16443 4440 16488 4468
rect 14507 4437 14519 4440
rect 14461 4431 14519 4437
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 20165 4471 20223 4477
rect 20165 4468 20177 4471
rect 16632 4440 20177 4468
rect 16632 4428 16638 4440
rect 20165 4437 20177 4440
rect 20211 4437 20223 4471
rect 20898 4468 20904 4480
rect 20859 4440 20904 4468
rect 20165 4431 20223 4437
rect 20898 4428 20904 4440
rect 20956 4428 20962 4480
rect 21450 4468 21456 4480
rect 21411 4440 21456 4468
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 22738 4428 22744 4480
rect 22796 4468 22802 4480
rect 23293 4471 23351 4477
rect 23293 4468 23305 4471
rect 22796 4440 23305 4468
rect 22796 4428 22802 4440
rect 23293 4437 23305 4440
rect 23339 4437 23351 4471
rect 23293 4431 23351 4437
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 5718 4264 5724 4276
rect 4663 4236 5724 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 17218 4264 17224 4276
rect 8312 4236 12434 4264
rect 17179 4236 17224 4264
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 7742 4088 7748 4100
rect 7800 4128 7806 4140
rect 8312 4128 8340 4236
rect 10778 4196 10784 4208
rect 9508 4168 10784 4196
rect 7800 4100 8340 4128
rect 8849 4131 8907 4137
rect 7800 4088 7806 4100
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9508 4128 9536 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 12406 4196 12434 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 20441 4267 20499 4273
rect 19260 4236 20392 4264
rect 19260 4196 19288 4236
rect 19426 4196 19432 4208
rect 12406 4168 19288 4196
rect 19352 4168 19432 4196
rect 8895 4100 9536 4128
rect 9576 4131 9634 4137
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9576 4097 9588 4131
rect 9622 4128 9634 4131
rect 9858 4128 9864 4140
rect 9622 4100 9864 4128
rect 9622 4097 9634 4100
rect 9576 4091 9634 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12693 4131 12751 4137
rect 12693 4128 12705 4131
rect 12032 4100 12705 4128
rect 12032 4088 12038 4100
rect 12693 4097 12705 4100
rect 12739 4097 12751 4131
rect 12693 4091 12751 4097
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14550 4137 14556 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 14240 4100 14289 4128
rect 14240 4088 14246 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14544 4128 14556 4137
rect 14511 4100 14556 4128
rect 14277 4091 14335 4097
rect 14544 4091 14556 4100
rect 14550 4088 14556 4091
rect 14608 4088 14614 4140
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 16448 4100 17325 4128
rect 16448 4088 16454 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 19352 4128 19380 4168
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 19978 4156 19984 4208
rect 20036 4196 20042 4208
rect 20257 4199 20315 4205
rect 20257 4196 20269 4199
rect 20036 4168 20269 4196
rect 20036 4156 20042 4168
rect 20257 4165 20269 4168
rect 20303 4165 20315 4199
rect 20364 4196 20392 4236
rect 20441 4233 20453 4267
rect 20487 4264 20499 4267
rect 20622 4264 20628 4276
rect 20487 4236 20628 4264
rect 20487 4233 20499 4236
rect 20441 4227 20499 4233
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 22066 4236 23428 4264
rect 20714 4196 20720 4208
rect 20364 4168 20720 4196
rect 20257 4159 20315 4165
rect 20714 4156 20720 4168
rect 20772 4196 20778 4208
rect 20993 4199 21051 4205
rect 20993 4196 21005 4199
rect 20772 4168 21005 4196
rect 20772 4156 20778 4168
rect 20993 4165 21005 4168
rect 21039 4196 21051 4199
rect 21634 4196 21640 4208
rect 21039 4168 21640 4196
rect 21039 4165 21051 4168
rect 20993 4159 21051 4165
rect 21634 4156 21640 4168
rect 21692 4196 21698 4208
rect 22066 4196 22094 4236
rect 22278 4205 22284 4208
rect 22272 4196 22284 4205
rect 21692 4168 22094 4196
rect 22239 4168 22284 4196
rect 21692 4156 21698 4168
rect 22272 4159 22284 4168
rect 22278 4156 22284 4159
rect 22336 4156 22342 4208
rect 17313 4091 17371 4097
rect 17420 4100 19380 4128
rect 19541 4131 19599 4137
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 10468 4032 12449 4060
rect 10468 4020 10474 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 17420 4069 17448 4100
rect 19541 4097 19553 4131
rect 19587 4128 19599 4131
rect 20070 4128 20076 4140
rect 19587 4100 20076 4128
rect 19587 4097 19599 4100
rect 19541 4091 19599 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 23400 4128 23428 4236
rect 22112 4100 23152 4128
rect 23400 4100 23980 4128
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 16816 4032 17417 4060
rect 16816 4020 16822 4032
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 20898 4060 20904 4072
rect 19843 4032 20904 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 20898 4020 20904 4032
rect 20956 4020 20962 4072
rect 22112 4060 22140 4100
rect 21376 4032 22140 4060
rect 21376 4004 21404 4032
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 12342 3992 12348 4004
rect 10735 3964 12348 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 15344 3964 16865 3992
rect 15344 3952 15350 3964
rect 16853 3961 16865 3964
rect 16899 3961 16911 3995
rect 21358 3992 21364 4004
rect 21319 3964 21364 3992
rect 16853 3955 16911 3961
rect 21358 3952 21364 3964
rect 21416 3952 21422 4004
rect 23124 3992 23152 4100
rect 23198 3992 23204 4004
rect 23111 3964 23204 3992
rect 23198 3952 23204 3964
rect 23256 3992 23262 4004
rect 23382 3992 23388 4004
rect 23256 3964 23388 3992
rect 23256 3952 23262 3964
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 23952 3936 23980 4100
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 9306 3924 9312 3936
rect 8711 3896 9312 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 11974 3924 11980 3936
rect 11935 3896 11980 3924
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 15562 3924 15568 3936
rect 13863 3896 15568 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 16114 3924 16120 3936
rect 15712 3896 15757 3924
rect 16075 3896 16120 3924
rect 15712 3884 15718 3896
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 18417 3927 18475 3933
rect 18417 3893 18429 3927
rect 18463 3924 18475 3927
rect 19610 3924 19616 3936
rect 18463 3896 19616 3924
rect 18463 3893 18475 3896
rect 18417 3887 18475 3893
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 20254 3924 20260 3936
rect 20215 3896 20260 3924
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 21453 3927 21511 3933
rect 21453 3893 21465 3927
rect 21499 3924 21511 3927
rect 22922 3924 22928 3936
rect 21499 3896 22928 3924
rect 21499 3893 21511 3896
rect 21453 3887 21511 3893
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9582 3720 9588 3732
rect 9263 3692 9588 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9582 3680 9588 3692
rect 9640 3720 9646 3732
rect 11698 3720 11704 3732
rect 9640 3692 11704 3720
rect 9640 3680 9646 3692
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 11885 3723 11943 3729
rect 11885 3689 11897 3723
rect 11931 3720 11943 3723
rect 12250 3720 12256 3732
rect 11931 3692 12256 3720
rect 11931 3689 11943 3692
rect 11885 3683 11943 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 13354 3720 13360 3732
rect 12360 3692 13360 3720
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 12360 3652 12388 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 16298 3720 16304 3732
rect 15519 3692 16304 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 20346 3720 20352 3732
rect 18555 3692 20352 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 22186 3680 22192 3732
rect 22244 3720 22250 3732
rect 23106 3720 23112 3732
rect 22244 3692 22600 3720
rect 23067 3692 23112 3720
rect 22244 3680 22250 3692
rect 20162 3652 20168 3664
rect 11572 3624 12388 3652
rect 20123 3624 20168 3652
rect 11572 3612 11578 3624
rect 20162 3612 20168 3624
rect 20220 3612 20226 3664
rect 8294 3584 8300 3596
rect 7760 3556 8300 3584
rect 7760 3525 7788 3556
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 8527 3556 10517 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14642 3584 14648 3596
rect 13872 3556 14648 3584
rect 13872 3544 13878 3556
rect 14642 3544 14648 3556
rect 14700 3584 14706 3596
rect 14829 3587 14887 3593
rect 14829 3584 14841 3587
rect 14700 3556 14841 3584
rect 14700 3544 14706 3556
rect 14829 3553 14841 3556
rect 14875 3553 14887 3587
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 14829 3547 14887 3553
rect 16960 3556 17969 3584
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 7745 3479 7803 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 9398 3516 9404 3528
rect 9359 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 11698 3476 11704 3528
rect 11756 3516 11762 3528
rect 12345 3519 12403 3525
rect 12345 3516 12357 3519
rect 11756 3488 12357 3516
rect 11756 3476 11762 3488
rect 12345 3485 12357 3488
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 10750 3451 10808 3457
rect 10750 3448 10762 3451
rect 9732 3420 10762 3448
rect 9732 3408 9738 3420
rect 10750 3417 10762 3420
rect 10796 3417 10808 3451
rect 12158 3448 12164 3460
rect 10750 3411 10808 3417
rect 11808 3420 12164 3448
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3380 7987 3383
rect 9122 3380 9128 3392
rect 7975 3352 9128 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9953 3383 10011 3389
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 11808 3380 11836 3420
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 12590 3451 12648 3457
rect 12590 3448 12602 3451
rect 12406 3420 12602 3448
rect 9999 3352 11836 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 12406 3380 12434 3420
rect 12590 3417 12602 3420
rect 12636 3417 12648 3451
rect 14844 3448 14872 3547
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15286 3516 15292 3528
rect 15151 3488 15292 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15930 3516 15936 3528
rect 15891 3488 15936 3516
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16200 3519 16258 3525
rect 16200 3485 16212 3519
rect 16246 3516 16258 3519
rect 16574 3516 16580 3528
rect 16246 3488 16580 3516
rect 16246 3485 16258 3488
rect 16200 3479 16258 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16960 3448 16988 3556
rect 17957 3553 17969 3556
rect 18003 3584 18015 3587
rect 19518 3584 19524 3596
rect 18003 3556 19524 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 22572 3593 22600 3692
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 23569 3723 23627 3729
rect 23569 3720 23581 3723
rect 23216 3692 23581 3720
rect 22557 3587 22615 3593
rect 22557 3553 22569 3587
rect 22603 3553 22615 3587
rect 22557 3547 22615 3553
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 19702 3476 19708 3528
rect 19760 3516 19766 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 19760 3488 19809 3516
rect 19760 3476 19766 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 22301 3519 22359 3525
rect 22301 3485 22313 3519
rect 22347 3516 22359 3519
rect 22738 3516 22744 3528
rect 22347 3488 22744 3516
rect 22347 3485 22359 3488
rect 22301 3479 22359 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 23216 3460 23244 3692
rect 23569 3689 23581 3692
rect 23615 3689 23627 3723
rect 23569 3683 23627 3689
rect 23477 3655 23535 3661
rect 23477 3621 23489 3655
rect 23523 3621 23535 3655
rect 23477 3615 23535 3621
rect 23382 3584 23388 3596
rect 23343 3556 23388 3584
rect 23382 3544 23388 3556
rect 23440 3544 23446 3596
rect 23492 3584 23520 3615
rect 23566 3584 23572 3596
rect 23492 3556 23572 3584
rect 23566 3544 23572 3556
rect 23624 3544 23630 3596
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23937 3519 23995 3525
rect 23937 3516 23949 3519
rect 23532 3488 23949 3516
rect 23532 3476 23538 3488
rect 23937 3485 23949 3488
rect 23983 3485 23995 3519
rect 23937 3479 23995 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 14844 3420 16988 3448
rect 12590 3411 12648 3417
rect 21450 3408 21456 3460
rect 21508 3448 21514 3460
rect 23198 3448 23204 3460
rect 21508 3420 23204 3448
rect 21508 3408 21514 3420
rect 23198 3408 23204 3420
rect 23256 3408 23262 3460
rect 24780 3448 24808 3479
rect 23308 3420 24808 3448
rect 23308 3392 23336 3420
rect 11940 3352 12434 3380
rect 11940 3340 11946 3352
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13725 3383 13783 3389
rect 13725 3380 13737 3383
rect 13044 3352 13737 3380
rect 13044 3340 13050 3352
rect 13725 3349 13737 3352
rect 13771 3349 13783 3383
rect 13725 3343 13783 3349
rect 15013 3383 15071 3389
rect 15013 3349 15025 3383
rect 15059 3380 15071 3383
rect 16298 3380 16304 3392
rect 15059 3352 16304 3380
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 17310 3380 17316 3392
rect 17223 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3380 17374 3392
rect 18049 3383 18107 3389
rect 18049 3380 18061 3383
rect 17368 3352 18061 3380
rect 17368 3340 17374 3352
rect 18049 3349 18061 3352
rect 18095 3349 18107 3383
rect 18049 3343 18107 3349
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 19705 3383 19763 3389
rect 19705 3380 19717 3383
rect 19668 3352 19717 3380
rect 19668 3340 19674 3352
rect 19705 3349 19717 3352
rect 19751 3349 19763 3383
rect 19705 3343 19763 3349
rect 20990 3340 20996 3392
rect 21048 3380 21054 3392
rect 21177 3383 21235 3389
rect 21177 3380 21189 3383
rect 21048 3352 21189 3380
rect 21048 3340 21054 3352
rect 21177 3349 21189 3352
rect 21223 3380 21235 3383
rect 22370 3380 22376 3392
rect 21223 3352 22376 3380
rect 21223 3349 21235 3352
rect 21177 3343 21235 3349
rect 22370 3340 22376 3352
rect 22428 3340 22434 3392
rect 23290 3340 23296 3392
rect 23348 3340 23354 3392
rect 24578 3380 24584 3392
rect 24539 3352 24584 3380
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 11146 3176 11152 3188
rect 9180 3148 9996 3176
rect 11107 3148 11152 3176
rect 9180 3136 9186 3148
rect 8386 3068 8392 3120
rect 8444 3108 8450 3120
rect 9858 3108 9864 3120
rect 8444 3080 9864 3108
rect 8444 3068 8450 3080
rect 8496 3049 8524 3080
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 9968 3108 9996 3148
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 15197 3179 15255 3185
rect 15197 3176 15209 3179
rect 11848 3148 15209 3176
rect 11848 3136 11854 3148
rect 15197 3145 15209 3148
rect 15243 3145 15255 3179
rect 15197 3139 15255 3145
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15620 3148 15669 3176
rect 15620 3136 15626 3148
rect 15657 3145 15669 3148
rect 15703 3176 15715 3179
rect 16022 3176 16028 3188
rect 15703 3148 16028 3176
rect 15703 3145 15715 3148
rect 15657 3139 15715 3145
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19978 3176 19984 3188
rect 19576 3148 19984 3176
rect 19576 3136 19582 3148
rect 19978 3136 19984 3148
rect 20036 3176 20042 3188
rect 20165 3179 20223 3185
rect 20165 3176 20177 3179
rect 20036 3148 20177 3176
rect 20036 3136 20042 3148
rect 20165 3145 20177 3148
rect 20211 3145 20223 3179
rect 20165 3139 20223 3145
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3145 20867 3179
rect 22462 3176 22468 3188
rect 20809 3139 20867 3145
rect 22066 3148 22468 3176
rect 10025 3111 10083 3117
rect 10025 3108 10037 3111
rect 9968 3080 10037 3108
rect 10025 3077 10037 3080
rect 10071 3077 10083 3111
rect 10025 3071 10083 3077
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11882 3108 11888 3120
rect 11112 3080 11888 3108
rect 11112 3068 11118 3080
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 14737 3111 14795 3117
rect 14737 3077 14749 3111
rect 14783 3108 14795 3111
rect 16482 3108 16488 3120
rect 14783 3080 16488 3108
rect 14783 3077 14795 3080
rect 14737 3071 14795 3077
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 8481 3043 8539 3049
rect 1903 3012 2774 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2746 2904 2774 3012
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 9272 3012 9321 3040
rect 9272 3000 9278 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 11793 3043 11851 3049
rect 9456 3012 10824 3040
rect 9456 3000 9462 3012
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 8619 2944 9781 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 9125 2907 9183 2913
rect 9125 2904 9137 2907
rect 2746 2876 9137 2904
rect 9125 2873 9137 2876
rect 9171 2873 9183 2907
rect 10796 2904 10824 3012
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 12066 3040 12072 3052
rect 11839 3012 12072 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 15565 3003 15623 3009
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 11020 2944 13001 2972
rect 11020 2932 11026 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 15580 2904 15608 3003
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 18874 3040 18880 3052
rect 18932 3049 18938 3052
rect 18844 3012 18880 3040
rect 18874 3000 18880 3012
rect 18932 3003 18944 3049
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19334 3040 19340 3052
rect 19199 3012 19340 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 18932 3000 18938 3003
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 20824 3040 20852 3139
rect 22066 3108 22094 3148
rect 22462 3136 22468 3148
rect 22520 3176 22526 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 22520 3148 23397 3176
rect 22520 3136 22526 3148
rect 23385 3145 23397 3148
rect 23431 3176 23443 3179
rect 23566 3176 23572 3188
rect 23431 3148 23572 3176
rect 23431 3145 23443 3148
rect 23385 3139 23443 3145
rect 23566 3136 23572 3148
rect 23624 3176 23630 3188
rect 23842 3176 23848 3188
rect 23624 3148 23848 3176
rect 23624 3136 23630 3148
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 23934 3136 23940 3188
rect 23992 3176 23998 3188
rect 25225 3179 25283 3185
rect 25225 3176 25237 3179
rect 23992 3148 25237 3176
rect 23992 3136 23998 3148
rect 25225 3145 25237 3148
rect 25271 3145 25283 3179
rect 25225 3139 25283 3145
rect 21192 3080 22094 3108
rect 22272 3111 22330 3117
rect 20990 3040 20996 3052
rect 20395 3012 20852 3040
rect 20951 3012 20996 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21192 3049 21220 3080
rect 22272 3077 22284 3111
rect 22318 3108 22330 3111
rect 24578 3108 24584 3120
rect 22318 3080 24584 3108
rect 22318 3077 22330 3080
rect 22272 3071 22330 3077
rect 24578 3068 24584 3080
rect 24636 3068 24642 3120
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3009 21235 3043
rect 21450 3040 21456 3052
rect 21411 3012 21456 3040
rect 21177 3003 21235 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 22005 3043 22063 3049
rect 22005 3009 22017 3043
rect 22051 3040 22063 3043
rect 22094 3040 22100 3052
rect 22051 3012 22100 3040
rect 22051 3009 22063 3012
rect 22005 3003 22063 3009
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 23198 3000 23204 3052
rect 23256 3040 23262 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23256 3012 23857 3040
rect 23256 3000 23262 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 23845 3003 23903 3009
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 10796 2876 15608 2904
rect 15672 2944 15761 2972
rect 9125 2867 9183 2873
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 624 2808 1685 2836
rect 624 2796 630 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 6086 2796 6092 2848
rect 6144 2836 6150 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6144 2808 6561 2836
rect 6144 2796 6150 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 7190 2836 7196 2848
rect 7151 2808 7196 2836
rect 6549 2799 6607 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 8294 2836 8300 2848
rect 8067 2808 8300 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 9140 2836 9168 2867
rect 11514 2836 11520 2848
rect 9140 2808 11520 2836
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 12710 2836 12716 2848
rect 12483 2808 12716 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 14642 2796 14648 2848
rect 14700 2836 14706 2848
rect 15672 2836 15700 2944
rect 15749 2941 15761 2944
rect 15795 2941 15807 2975
rect 15749 2935 15807 2941
rect 28353 2975 28411 2981
rect 28353 2941 28365 2975
rect 28399 2972 28411 2975
rect 29270 2972 29276 2984
rect 28399 2944 29276 2972
rect 28399 2941 28411 2944
rect 28353 2935 28411 2941
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 24029 2907 24087 2913
rect 24029 2904 24041 2907
rect 22940 2876 24041 2904
rect 17126 2836 17132 2848
rect 14700 2808 15700 2836
rect 17087 2808 17132 2836
rect 14700 2796 14706 2808
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17773 2839 17831 2845
rect 17773 2805 17785 2839
rect 17819 2836 17831 2839
rect 18138 2836 18144 2848
rect 17819 2808 18144 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 21358 2836 21364 2848
rect 21319 2808 21364 2836
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 22940 2836 22968 2876
rect 24029 2873 24041 2876
rect 24075 2873 24087 2907
rect 24029 2867 24087 2873
rect 24486 2864 24492 2916
rect 24544 2904 24550 2916
rect 24581 2907 24639 2913
rect 24581 2904 24593 2907
rect 24544 2876 24593 2904
rect 24544 2864 24550 2876
rect 24581 2873 24593 2876
rect 24627 2873 24639 2907
rect 24581 2867 24639 2873
rect 22704 2808 22968 2836
rect 22704 2796 22710 2808
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 8478 2632 8484 2644
rect 6886 2604 8484 2632
rect 6886 2564 6914 2604
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9674 2632 9680 2644
rect 8619 2604 9680 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 11698 2632 11704 2644
rect 10367 2604 11704 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 12529 2635 12587 2641
rect 12529 2632 12541 2635
rect 12360 2604 12541 2632
rect 3160 2536 6914 2564
rect 7929 2567 7987 2573
rect 3160 2437 3188 2536
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 10502 2564 10508 2576
rect 7975 2536 10508 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 7285 2499 7343 2505
rect 4264 2468 7236 2496
rect 4264 2437 4292 2468
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 2056 2360 2084 2391
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 5040 2400 5089 2428
rect 5040 2388 5046 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 7208 2360 7236 2468
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 9398 2496 9404 2508
rect 7331 2468 9404 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 12360 2496 12388 2604
rect 12529 2601 12541 2604
rect 12575 2601 12587 2635
rect 12529 2595 12587 2601
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 15930 2632 15936 2644
rect 14415 2604 15936 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16298 2632 16304 2644
rect 16259 2604 16304 2632
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 18874 2632 18880 2644
rect 18371 2604 18880 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 21542 2592 21548 2644
rect 21600 2632 21606 2644
rect 23845 2635 23903 2641
rect 23845 2632 23857 2635
rect 21600 2604 23857 2632
rect 21600 2592 21606 2604
rect 23845 2601 23857 2604
rect 23891 2601 23903 2635
rect 23845 2595 23903 2601
rect 12820 2536 14964 2564
rect 9600 2468 12388 2496
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 9600 2437 9628 2468
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12820 2496 12848 2536
rect 12986 2496 12992 2508
rect 12584 2468 12848 2496
rect 12947 2468 12992 2496
rect 12584 2456 12590 2468
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13814 2496 13820 2508
rect 13219 2468 13820 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 14936 2505 14964 2536
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 16080 2536 17632 2564
rect 16080 2524 16086 2536
rect 14921 2499 14979 2505
rect 14921 2465 14933 2499
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9916 2400 10241 2428
rect 9916 2388 9922 2400
rect 10229 2397 10241 2400
rect 10275 2428 10287 2431
rect 10778 2428 10784 2440
rect 10275 2400 10784 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11146 2428 11152 2440
rect 11107 2400 11152 2428
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 13004 2428 13032 2456
rect 12115 2400 13032 2428
rect 14461 2431 14519 2437
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 15470 2428 15476 2440
rect 14507 2400 15476 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 17604 2437 17632 2536
rect 18524 2536 19196 2564
rect 18524 2437 18552 2536
rect 19168 2496 19196 2536
rect 19334 2524 19340 2576
rect 19392 2564 19398 2576
rect 20349 2567 20407 2573
rect 20349 2564 20361 2567
rect 19392 2536 20361 2564
rect 19392 2524 19398 2536
rect 20349 2533 20361 2536
rect 20395 2533 20407 2567
rect 20349 2527 20407 2533
rect 21361 2567 21419 2573
rect 21361 2533 21373 2567
rect 21407 2564 21419 2567
rect 21450 2564 21456 2576
rect 21407 2536 21456 2564
rect 21407 2533 21419 2536
rect 21361 2527 21419 2533
rect 21450 2524 21456 2536
rect 21508 2524 21514 2576
rect 22370 2564 22376 2576
rect 22283 2536 22376 2564
rect 22370 2524 22376 2536
rect 22428 2564 22434 2576
rect 22922 2564 22928 2576
rect 22428 2536 22928 2564
rect 22428 2524 22434 2536
rect 22922 2524 22928 2536
rect 22980 2524 22986 2576
rect 23017 2567 23075 2573
rect 23017 2533 23029 2567
rect 23063 2533 23075 2567
rect 23017 2527 23075 2533
rect 20254 2496 20260 2508
rect 19168 2468 20260 2496
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 23032 2496 23060 2527
rect 23750 2524 23756 2576
rect 23808 2564 23814 2576
rect 24765 2567 24823 2573
rect 24765 2564 24777 2567
rect 23808 2536 24777 2564
rect 23808 2524 23814 2536
rect 24765 2533 24777 2536
rect 24811 2533 24823 2567
rect 24765 2527 24823 2533
rect 20496 2468 23060 2496
rect 20496 2456 20502 2468
rect 23106 2456 23112 2508
rect 23164 2496 23170 2508
rect 23164 2468 23428 2496
rect 23164 2456 23170 2468
rect 23400 2440 23428 2468
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17589 2431 17647 2437
rect 17589 2397 17601 2431
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 18509 2431 18567 2437
rect 18509 2397 18521 2431
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 19150 2428 19156 2440
rect 18831 2400 19156 2428
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19300 2400 19441 2428
rect 19300 2388 19306 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19610 2388 19616 2440
rect 19668 2428 19674 2440
rect 20165 2431 20223 2437
rect 20165 2428 20177 2431
rect 19668 2400 20177 2428
rect 19668 2388 19674 2400
rect 20165 2397 20177 2400
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20772 2400 21005 2428
rect 20772 2388 20778 2400
rect 20993 2397 21005 2400
rect 21039 2428 21051 2431
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21039 2400 22017 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 23198 2428 23204 2440
rect 23159 2400 23204 2428
rect 22005 2391 22063 2397
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 23440 2400 23673 2428
rect 23440 2388 23446 2400
rect 23661 2397 23673 2400
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23900 2400 24593 2428
rect 23900 2388 23906 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25317 2431 25375 2437
rect 25317 2428 25329 2431
rect 24912 2400 25329 2428
rect 24912 2388 24918 2400
rect 25317 2397 25329 2400
rect 25363 2397 25375 2431
rect 25317 2391 25375 2397
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 26016 2400 26065 2428
rect 26016 2388 26022 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 28166 2428 28172 2440
rect 28127 2400 28172 2428
rect 27157 2391 27215 2397
rect 28166 2388 28172 2400
rect 28224 2388 28230 2440
rect 9306 2360 9312 2372
rect 2056 2332 6914 2360
rect 7208 2332 9312 2360
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 1728 2264 1869 2292
rect 1728 2252 1734 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2832 2264 2973 2292
rect 2832 2252 2838 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 6886 2292 6914 2332
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 11054 2360 11060 2372
rect 9784 2332 11060 2360
rect 9582 2292 9588 2304
rect 6886 2264 9588 2292
rect 4065 2255 4123 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 9784 2301 9812 2332
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 13814 2360 13820 2372
rect 11900 2332 13820 2360
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10965 2295 11023 2301
rect 10965 2261 10977 2295
rect 11011 2292 11023 2295
rect 11606 2292 11612 2304
rect 11011 2264 11612 2292
rect 11011 2261 11023 2264
rect 10965 2255 11023 2261
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 11900 2301 11928 2332
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 15188 2363 15246 2369
rect 15188 2329 15200 2363
rect 15234 2329 15246 2363
rect 15188 2323 15246 2329
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2261 11943 2295
rect 12894 2292 12900 2304
rect 12855 2264 12900 2292
rect 11885 2255 11943 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 15212 2292 15240 2323
rect 15286 2320 15292 2372
rect 15344 2360 15350 2372
rect 15344 2332 17816 2360
rect 15344 2320 15350 2332
rect 16114 2292 16120 2304
rect 15212 2264 16120 2292
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 17788 2301 17816 2332
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 23290 2360 23296 2372
rect 18288 2332 19656 2360
rect 18288 2320 18294 2332
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16448 2264 17049 2292
rect 16448 2252 16454 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17773 2295 17831 2301
rect 17773 2261 17785 2295
rect 17819 2261 17831 2295
rect 17773 2255 17831 2261
rect 18138 2252 18144 2304
rect 18196 2292 18202 2304
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 18196 2264 18705 2292
rect 18196 2252 18202 2264
rect 18693 2261 18705 2264
rect 18739 2292 18751 2295
rect 19242 2292 19248 2304
rect 18739 2264 19248 2292
rect 18739 2261 18751 2264
rect 18693 2255 18751 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19628 2301 19656 2332
rect 22388 2332 23296 2360
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 21453 2295 21511 2301
rect 21453 2261 21465 2295
rect 21499 2292 21511 2295
rect 22388 2292 22416 2332
rect 23290 2320 23296 2332
rect 23348 2320 23354 2372
rect 21499 2264 22416 2292
rect 22465 2295 22523 2301
rect 21499 2261 21511 2264
rect 21453 2255 21511 2261
rect 22465 2261 22477 2295
rect 22511 2292 22523 2295
rect 24762 2292 24768 2304
rect 22511 2264 24768 2292
rect 22511 2261 22523 2264
rect 22465 2255 22523 2261
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 8386 2048 8392 2100
rect 8444 2088 8450 2100
rect 11238 2088 11244 2100
rect 8444 2060 11244 2088
rect 8444 2048 8450 2060
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 8478 1980 8484 2032
rect 8536 2020 8542 2032
rect 12894 2020 12900 2032
rect 8536 1992 12900 2020
rect 8536 1980 8542 1992
rect 12894 1980 12900 1992
rect 12952 1980 12958 2032
<< via1 >>
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 3792 27548 3844 27600
rect 8576 27591 8628 27600
rect 8576 27557 8585 27591
rect 8585 27557 8619 27591
rect 8619 27557 8628 27591
rect 8576 27548 8628 27557
rect 6552 27455 6604 27464
rect 6552 27421 6561 27455
rect 6561 27421 6595 27455
rect 6595 27421 6604 27455
rect 6552 27412 6604 27421
rect 17868 27548 17920 27600
rect 21180 27548 21232 27600
rect 23664 27548 23716 27600
rect 26148 27548 26200 27600
rect 17776 27480 17828 27532
rect 11244 27412 11296 27464
rect 12624 27455 12676 27464
rect 12624 27421 12633 27455
rect 12633 27421 12667 27455
rect 12667 27421 12676 27455
rect 12624 27412 12676 27421
rect 12808 27455 12860 27464
rect 12808 27421 12817 27455
rect 12817 27421 12851 27455
rect 12851 27421 12860 27455
rect 12808 27412 12860 27421
rect 13820 27412 13872 27464
rect 16212 27412 16264 27464
rect 18696 27412 18748 27464
rect 28356 27455 28408 27464
rect 28356 27421 28365 27455
rect 28365 27421 28399 27455
rect 28399 27421 28408 27455
rect 28356 27412 28408 27421
rect 17960 27344 18012 27396
rect 4160 27319 4212 27328
rect 4160 27285 4169 27319
rect 4169 27285 4203 27319
rect 4203 27285 4212 27319
rect 4160 27276 4212 27285
rect 6736 27319 6788 27328
rect 6736 27285 6745 27319
rect 6745 27285 6779 27319
rect 6779 27285 6788 27319
rect 6736 27276 6788 27285
rect 10140 27276 10192 27328
rect 10876 27319 10928 27328
rect 10876 27285 10885 27319
rect 10885 27285 10919 27319
rect 10919 27285 10928 27319
rect 10876 27276 10928 27285
rect 12992 27276 13044 27328
rect 15200 27276 15252 27328
rect 15292 27276 15344 27328
rect 17684 27276 17736 27328
rect 23756 27319 23808 27328
rect 23756 27285 23765 27319
rect 23765 27285 23799 27319
rect 23799 27285 23808 27319
rect 23756 27276 23808 27285
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 9864 27072 9916 27124
rect 10876 27072 10928 27124
rect 8944 27004 8996 27056
rect 12716 27004 12768 27056
rect 12900 27004 12952 27056
rect 14004 27004 14056 27056
rect 8392 26936 8444 26988
rect 9404 26868 9456 26920
rect 10692 26936 10744 26988
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 11796 26936 11848 26988
rect 12808 26936 12860 26988
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 12256 26868 12308 26920
rect 13176 26868 13228 26920
rect 6736 26800 6788 26852
rect 9956 26732 10008 26784
rect 10048 26775 10100 26784
rect 10048 26741 10057 26775
rect 10057 26741 10091 26775
rect 10091 26741 10100 26775
rect 10048 26732 10100 26741
rect 11152 26732 11204 26784
rect 12348 26800 12400 26852
rect 13084 26732 13136 26784
rect 13636 26732 13688 26784
rect 14280 26732 14332 26784
rect 17040 26775 17092 26784
rect 17040 26741 17049 26775
rect 17049 26741 17083 26775
rect 17083 26741 17092 26775
rect 17040 26732 17092 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 10692 26528 10744 26580
rect 11152 26571 11204 26580
rect 11152 26537 11161 26571
rect 11161 26537 11195 26571
rect 11195 26537 11204 26571
rect 11152 26528 11204 26537
rect 12900 26528 12952 26580
rect 13268 26528 13320 26580
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 9312 26324 9364 26376
rect 4068 26299 4120 26308
rect 4068 26265 4077 26299
rect 4077 26265 4111 26299
rect 4111 26265 4120 26299
rect 4068 26256 4120 26265
rect 8484 26299 8536 26308
rect 8484 26265 8493 26299
rect 8493 26265 8527 26299
rect 8527 26265 8536 26299
rect 9956 26324 10008 26376
rect 10600 26367 10652 26376
rect 10600 26333 10609 26367
rect 10609 26333 10643 26367
rect 10643 26333 10652 26367
rect 10600 26324 10652 26333
rect 10968 26324 11020 26376
rect 12256 26460 12308 26512
rect 12624 26392 12676 26444
rect 13084 26460 13136 26512
rect 11796 26324 11848 26376
rect 12348 26367 12400 26376
rect 12348 26333 12357 26367
rect 12357 26333 12391 26367
rect 12391 26333 12400 26367
rect 12348 26324 12400 26333
rect 8484 26256 8536 26265
rect 2136 26231 2188 26240
rect 2136 26197 2145 26231
rect 2145 26197 2179 26231
rect 2179 26197 2188 26231
rect 2136 26188 2188 26197
rect 2596 26231 2648 26240
rect 2596 26197 2605 26231
rect 2605 26197 2639 26231
rect 2639 26197 2648 26231
rect 2596 26188 2648 26197
rect 3148 26188 3200 26240
rect 6460 26188 6512 26240
rect 8300 26188 8352 26240
rect 9772 26231 9824 26240
rect 9772 26197 9781 26231
rect 9781 26197 9815 26231
rect 9815 26197 9824 26231
rect 9772 26188 9824 26197
rect 13912 26392 13964 26444
rect 12900 26367 12952 26376
rect 12900 26333 12909 26367
rect 12909 26333 12943 26367
rect 12943 26333 12952 26367
rect 12900 26324 12952 26333
rect 13176 26367 13228 26376
rect 13176 26333 13185 26367
rect 13185 26333 13219 26367
rect 13219 26333 13228 26367
rect 13176 26324 13228 26333
rect 17040 26528 17092 26580
rect 15200 26392 15252 26444
rect 17776 26435 17828 26444
rect 17776 26401 17785 26435
rect 17785 26401 17819 26435
rect 17819 26401 17828 26435
rect 17776 26392 17828 26401
rect 18052 26392 18104 26444
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 23756 26460 23808 26512
rect 28172 26392 28224 26444
rect 26240 26324 26292 26376
rect 19524 26299 19576 26308
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 24952 26256 25004 26308
rect 14372 26231 14424 26240
rect 14372 26197 14381 26231
rect 14381 26197 14415 26231
rect 14415 26197 14424 26231
rect 14372 26188 14424 26197
rect 15660 26231 15712 26240
rect 15660 26197 15669 26231
rect 15669 26197 15703 26231
rect 15703 26197 15712 26231
rect 15660 26188 15712 26197
rect 16212 26188 16264 26240
rect 17132 26188 17184 26240
rect 18696 26188 18748 26240
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 2228 25848 2280 25900
rect 4068 25984 4120 26036
rect 10600 26027 10652 26036
rect 10600 25993 10609 26027
rect 10609 25993 10643 26027
rect 10643 25993 10652 26027
rect 10600 25984 10652 25993
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 11060 25984 11112 26036
rect 13176 25984 13228 26036
rect 9312 25916 9364 25968
rect 13452 25984 13504 26036
rect 14464 25984 14516 26036
rect 17960 25984 18012 26036
rect 14372 25916 14424 25968
rect 17868 25959 17920 25968
rect 17868 25925 17877 25959
rect 17877 25925 17911 25959
rect 17911 25925 17920 25959
rect 17868 25916 17920 25925
rect 8484 25848 8536 25900
rect 8944 25891 8996 25900
rect 8944 25857 8953 25891
rect 8953 25857 8987 25891
rect 8987 25857 8996 25891
rect 8944 25848 8996 25857
rect 9128 25848 9180 25900
rect 9956 25891 10008 25900
rect 9956 25857 9965 25891
rect 9965 25857 9999 25891
rect 9999 25857 10008 25891
rect 9956 25848 10008 25857
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 2596 25780 2648 25832
rect 6920 25780 6972 25832
rect 2688 25712 2740 25764
rect 12808 25891 12860 25900
rect 11152 25755 11204 25764
rect 11152 25721 11161 25755
rect 11161 25721 11195 25755
rect 11195 25721 11204 25755
rect 11152 25712 11204 25721
rect 3700 25644 3752 25696
rect 5816 25644 5868 25696
rect 7656 25687 7708 25696
rect 7656 25653 7665 25687
rect 7665 25653 7699 25687
rect 7699 25653 7708 25687
rect 7656 25644 7708 25653
rect 9772 25687 9824 25696
rect 9772 25653 9781 25687
rect 9781 25653 9815 25687
rect 9815 25653 9824 25687
rect 12808 25857 12817 25891
rect 12817 25857 12851 25891
rect 12851 25857 12860 25891
rect 12808 25848 12860 25857
rect 13268 25848 13320 25900
rect 14004 25891 14056 25900
rect 14004 25857 14013 25891
rect 14013 25857 14047 25891
rect 14047 25857 14056 25891
rect 14004 25848 14056 25857
rect 14096 25848 14148 25900
rect 16212 25891 16264 25900
rect 16212 25857 16221 25891
rect 16221 25857 16255 25891
rect 16255 25857 16264 25891
rect 16212 25848 16264 25857
rect 12716 25823 12768 25832
rect 12716 25789 12725 25823
rect 12725 25789 12759 25823
rect 12759 25789 12768 25823
rect 12716 25780 12768 25789
rect 13912 25823 13964 25832
rect 13912 25789 13921 25823
rect 13921 25789 13955 25823
rect 13955 25789 13964 25823
rect 13912 25780 13964 25789
rect 18052 25823 18104 25832
rect 18052 25789 18061 25823
rect 18061 25789 18095 25823
rect 18095 25789 18104 25823
rect 18052 25780 18104 25789
rect 18696 25780 18748 25832
rect 13176 25712 13228 25764
rect 16856 25712 16908 25764
rect 12072 25687 12124 25696
rect 9772 25644 9824 25653
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 12072 25644 12124 25653
rect 13360 25644 13412 25696
rect 15752 25644 15804 25696
rect 17224 25644 17276 25696
rect 17592 25644 17644 25696
rect 18696 25687 18748 25696
rect 18696 25653 18705 25687
rect 18705 25653 18739 25687
rect 18739 25653 18748 25687
rect 18696 25644 18748 25653
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 8484 25440 8536 25492
rect 8944 25372 8996 25424
rect 10048 25440 10100 25492
rect 11796 25483 11848 25492
rect 11796 25449 11805 25483
rect 11805 25449 11839 25483
rect 11839 25449 11848 25483
rect 11796 25440 11848 25449
rect 12900 25440 12952 25492
rect 5724 25304 5776 25356
rect 9404 25304 9456 25356
rect 3976 25236 4028 25288
rect 8668 25236 8720 25288
rect 9220 25236 9272 25288
rect 9680 25236 9732 25288
rect 10416 25236 10468 25288
rect 10876 25372 10928 25424
rect 10692 25347 10744 25356
rect 10692 25313 10701 25347
rect 10701 25313 10735 25347
rect 10735 25313 10744 25347
rect 10692 25304 10744 25313
rect 2228 25100 2280 25152
rect 3700 25100 3752 25152
rect 4712 25100 4764 25152
rect 5080 25143 5132 25152
rect 5080 25109 5089 25143
rect 5089 25109 5123 25143
rect 5123 25109 5132 25143
rect 5080 25100 5132 25109
rect 6460 25100 6512 25152
rect 9036 25168 9088 25220
rect 9588 25168 9640 25220
rect 9220 25100 9272 25152
rect 9404 25100 9456 25152
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 12808 25304 12860 25356
rect 13268 25304 13320 25356
rect 11152 25168 11204 25220
rect 11796 25168 11848 25220
rect 12716 25236 12768 25288
rect 13544 25279 13596 25288
rect 13544 25245 13553 25279
rect 13553 25245 13587 25279
rect 13587 25245 13596 25279
rect 13544 25236 13596 25245
rect 13636 25279 13688 25288
rect 13636 25245 13645 25279
rect 13645 25245 13679 25279
rect 13679 25245 13688 25279
rect 13636 25236 13688 25245
rect 15660 25236 15712 25288
rect 17132 25279 17184 25288
rect 17132 25245 17141 25279
rect 17141 25245 17175 25279
rect 17175 25245 17184 25279
rect 17132 25236 17184 25245
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 11060 25100 11112 25152
rect 14464 25100 14516 25152
rect 15936 25100 15988 25152
rect 16488 25100 16540 25152
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 2136 24896 2188 24948
rect 3792 24896 3844 24948
rect 5080 24896 5132 24948
rect 8944 24896 8996 24948
rect 9404 24896 9456 24948
rect 9128 24871 9180 24880
rect 9128 24837 9137 24871
rect 9137 24837 9171 24871
rect 9171 24837 9180 24871
rect 9128 24828 9180 24837
rect 8852 24760 8904 24812
rect 9220 24803 9272 24812
rect 4988 24692 5040 24744
rect 7012 24735 7064 24744
rect 7012 24701 7021 24735
rect 7021 24701 7055 24735
rect 7055 24701 7064 24735
rect 7012 24692 7064 24701
rect 8760 24692 8812 24744
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 9588 24760 9640 24812
rect 12716 24896 12768 24948
rect 11060 24828 11112 24880
rect 10600 24803 10652 24812
rect 9680 24692 9732 24744
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 10968 24760 11020 24812
rect 11796 24760 11848 24812
rect 13268 24803 13320 24812
rect 10876 24692 10928 24744
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13452 24803 13504 24812
rect 13452 24769 13461 24803
rect 13461 24769 13495 24803
rect 13495 24769 13504 24803
rect 13452 24760 13504 24769
rect 14096 24760 14148 24812
rect 17040 24760 17092 24812
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18696 24803 18748 24812
rect 18696 24769 18705 24803
rect 18705 24769 18739 24803
rect 18739 24769 18748 24803
rect 18696 24760 18748 24769
rect 5724 24624 5776 24676
rect 8576 24624 8628 24676
rect 2504 24599 2556 24608
rect 2504 24565 2513 24599
rect 2513 24565 2547 24599
rect 2547 24565 2556 24599
rect 2504 24556 2556 24565
rect 2688 24556 2740 24608
rect 3976 24556 4028 24608
rect 9772 24556 9824 24608
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 12808 24556 12860 24608
rect 14004 24556 14056 24608
rect 18052 24692 18104 24744
rect 19248 24760 19300 24812
rect 19432 24803 19484 24812
rect 19432 24769 19441 24803
rect 19441 24769 19475 24803
rect 19475 24769 19484 24803
rect 19616 24803 19668 24812
rect 19432 24760 19484 24769
rect 19616 24769 19625 24803
rect 19625 24769 19659 24803
rect 19659 24769 19668 24803
rect 19616 24760 19668 24769
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 17408 24624 17460 24676
rect 18236 24624 18288 24676
rect 18880 24624 18932 24676
rect 19432 24624 19484 24676
rect 21548 24692 21600 24744
rect 22284 24692 22336 24744
rect 22468 24803 22520 24812
rect 22468 24769 22480 24803
rect 22480 24769 22514 24803
rect 22514 24769 22520 24803
rect 23296 24803 23348 24812
rect 22468 24760 22520 24769
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 23112 24692 23164 24744
rect 15200 24556 15252 24608
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 18788 24599 18840 24608
rect 18788 24565 18797 24599
rect 18797 24565 18831 24599
rect 18831 24565 18840 24599
rect 18788 24556 18840 24565
rect 18972 24556 19024 24608
rect 22468 24624 22520 24676
rect 24492 24624 24544 24676
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 22100 24599 22152 24608
rect 22100 24565 22109 24599
rect 22109 24565 22143 24599
rect 22143 24565 22152 24599
rect 22100 24556 22152 24565
rect 22744 24556 22796 24608
rect 24676 24556 24728 24608
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 5724 24395 5776 24404
rect 5724 24361 5733 24395
rect 5733 24361 5767 24395
rect 5767 24361 5776 24395
rect 5724 24352 5776 24361
rect 8576 24352 8628 24404
rect 16580 24395 16632 24404
rect 4896 24284 4948 24336
rect 4988 24284 5040 24336
rect 6460 24284 6512 24336
rect 8760 24284 8812 24336
rect 3148 24148 3200 24200
rect 4988 24148 5040 24200
rect 9036 24216 9088 24268
rect 10876 24284 10928 24336
rect 5356 24148 5408 24200
rect 6460 24191 6512 24200
rect 6460 24157 6469 24191
rect 6469 24157 6503 24191
rect 6503 24157 6512 24191
rect 6460 24148 6512 24157
rect 7012 24148 7064 24200
rect 9220 24148 9272 24200
rect 9588 24191 9640 24200
rect 9588 24157 9597 24191
rect 9597 24157 9631 24191
rect 9631 24157 9640 24191
rect 10600 24216 10652 24268
rect 9588 24148 9640 24157
rect 9772 24148 9824 24200
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 17592 24395 17644 24404
rect 16580 24352 16632 24361
rect 17592 24361 17601 24395
rect 17601 24361 17635 24395
rect 17635 24361 17644 24395
rect 17592 24352 17644 24361
rect 19616 24352 19668 24404
rect 23112 24395 23164 24404
rect 23112 24361 23121 24395
rect 23121 24361 23155 24395
rect 23155 24361 23164 24395
rect 23112 24352 23164 24361
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 12808 24284 12860 24336
rect 4252 24080 4304 24132
rect 6276 24123 6328 24132
rect 6276 24089 6285 24123
rect 6285 24089 6319 24123
rect 6319 24089 6328 24123
rect 6276 24080 6328 24089
rect 9036 24080 9088 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 2228 24055 2280 24064
rect 2228 24021 2237 24055
rect 2237 24021 2271 24055
rect 2271 24021 2280 24055
rect 2228 24012 2280 24021
rect 3976 24012 4028 24064
rect 4804 24012 4856 24064
rect 5448 24012 5500 24064
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 8484 24055 8536 24064
rect 8484 24021 8493 24055
rect 8493 24021 8527 24055
rect 8527 24021 8536 24055
rect 8484 24012 8536 24021
rect 9312 24080 9364 24132
rect 10600 24012 10652 24064
rect 10968 24055 11020 24064
rect 10968 24021 10977 24055
rect 10977 24021 11011 24055
rect 11011 24021 11020 24055
rect 13912 24216 13964 24268
rect 22100 24284 22152 24336
rect 21272 24216 21324 24268
rect 22744 24259 22796 24268
rect 12072 24148 12124 24200
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 15200 24191 15252 24200
rect 15200 24157 15209 24191
rect 15209 24157 15243 24191
rect 15243 24157 15252 24191
rect 15200 24148 15252 24157
rect 18052 24148 18104 24200
rect 18696 24148 18748 24200
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 19248 24148 19300 24200
rect 14648 24080 14700 24132
rect 15752 24080 15804 24132
rect 19524 24123 19576 24132
rect 19524 24089 19533 24123
rect 19533 24089 19567 24123
rect 19567 24089 19576 24123
rect 19524 24080 19576 24089
rect 20076 24148 20128 24200
rect 22744 24225 22753 24259
rect 22753 24225 22787 24259
rect 22787 24225 22796 24259
rect 22744 24216 22796 24225
rect 23204 24216 23256 24268
rect 24676 24259 24728 24268
rect 24676 24225 24685 24259
rect 24685 24225 24719 24259
rect 24719 24225 24728 24259
rect 24676 24216 24728 24225
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 22468 24191 22520 24200
rect 10968 24012 11020 24021
rect 12900 24012 12952 24064
rect 13636 24055 13688 24064
rect 13636 24021 13645 24055
rect 13645 24021 13679 24055
rect 13679 24021 13688 24055
rect 13636 24012 13688 24021
rect 13820 24012 13872 24064
rect 17868 24012 17920 24064
rect 18512 24012 18564 24064
rect 19432 24012 19484 24064
rect 21272 24012 21324 24064
rect 22468 24157 22477 24191
rect 22477 24157 22511 24191
rect 22511 24157 22520 24191
rect 22468 24148 22520 24157
rect 22652 24191 22704 24200
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 22192 24080 22244 24132
rect 23480 24148 23532 24200
rect 23388 24080 23440 24132
rect 23756 24080 23808 24132
rect 23572 24012 23624 24064
rect 24860 24012 24912 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 2688 23808 2740 23860
rect 8760 23808 8812 23860
rect 9036 23851 9088 23860
rect 9036 23817 9045 23851
rect 9045 23817 9079 23851
rect 9079 23817 9088 23851
rect 9036 23808 9088 23817
rect 10140 23808 10192 23860
rect 10692 23808 10744 23860
rect 15752 23851 15804 23860
rect 15752 23817 15761 23851
rect 15761 23817 15795 23851
rect 15795 23817 15804 23851
rect 15752 23808 15804 23817
rect 16580 23808 16632 23860
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 18512 23851 18564 23860
rect 17408 23808 17460 23817
rect 1860 23783 1912 23792
rect 1860 23749 1869 23783
rect 1869 23749 1903 23783
rect 1903 23749 1912 23783
rect 1860 23740 1912 23749
rect 8484 23740 8536 23792
rect 9680 23740 9732 23792
rect 15200 23740 15252 23792
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 5356 23672 5408 23724
rect 5816 23715 5868 23724
rect 5816 23681 5825 23715
rect 5825 23681 5859 23715
rect 5859 23681 5868 23715
rect 5816 23672 5868 23681
rect 6368 23672 6420 23724
rect 7472 23672 7524 23724
rect 7288 23604 7340 23656
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 9864 23604 9916 23656
rect 3976 23536 4028 23588
rect 5264 23536 5316 23588
rect 9588 23536 9640 23588
rect 10600 23672 10652 23724
rect 10968 23715 11020 23724
rect 10968 23681 10977 23715
rect 10977 23681 11011 23715
rect 11011 23681 11020 23715
rect 10968 23672 11020 23681
rect 11704 23672 11756 23724
rect 12256 23672 12308 23724
rect 10232 23604 10284 23656
rect 12808 23672 12860 23724
rect 15844 23672 15896 23724
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 15200 23604 15252 23656
rect 2136 23468 2188 23520
rect 2872 23468 2924 23520
rect 4068 23468 4120 23520
rect 6736 23468 6788 23520
rect 9496 23468 9548 23520
rect 11244 23468 11296 23520
rect 12072 23468 12124 23520
rect 14004 23468 14056 23520
rect 16028 23536 16080 23588
rect 16856 23672 16908 23724
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 18512 23817 18521 23851
rect 18521 23817 18555 23851
rect 18555 23817 18564 23851
rect 18512 23808 18564 23817
rect 18696 23808 18748 23860
rect 22284 23808 22336 23860
rect 22376 23808 22428 23860
rect 23204 23808 23256 23860
rect 23296 23808 23348 23860
rect 17960 23740 18012 23792
rect 21456 23783 21508 23792
rect 21456 23749 21465 23783
rect 21465 23749 21499 23783
rect 21499 23749 21508 23783
rect 21456 23740 21508 23749
rect 20076 23715 20128 23724
rect 20076 23681 20085 23715
rect 20085 23681 20119 23715
rect 20119 23681 20128 23715
rect 20076 23672 20128 23681
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20444 23672 20496 23724
rect 18052 23604 18104 23656
rect 19248 23604 19300 23656
rect 18972 23579 19024 23588
rect 18972 23545 18981 23579
rect 18981 23545 19015 23579
rect 19015 23545 19024 23579
rect 18972 23536 19024 23545
rect 16396 23468 16448 23520
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 22744 23672 22796 23724
rect 23572 23715 23624 23724
rect 22284 23604 22336 23656
rect 22652 23604 22704 23656
rect 23572 23681 23581 23715
rect 23581 23681 23615 23715
rect 23615 23681 23624 23715
rect 23572 23672 23624 23681
rect 23756 23672 23808 23724
rect 24492 23715 24544 23724
rect 24492 23681 24501 23715
rect 24501 23681 24535 23715
rect 24535 23681 24544 23715
rect 24492 23672 24544 23681
rect 24584 23672 24636 23724
rect 25596 23672 25648 23724
rect 23480 23647 23532 23656
rect 23480 23613 23489 23647
rect 23489 23613 23523 23647
rect 23523 23613 23532 23647
rect 23480 23604 23532 23613
rect 19524 23511 19576 23520
rect 19524 23477 19533 23511
rect 19533 23477 19567 23511
rect 19567 23477 19576 23511
rect 19524 23468 19576 23477
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 22468 23536 22520 23588
rect 23204 23468 23256 23520
rect 23848 23511 23900 23520
rect 23848 23477 23857 23511
rect 23857 23477 23891 23511
rect 23891 23477 23900 23511
rect 23848 23468 23900 23477
rect 25136 23511 25188 23520
rect 25136 23477 25145 23511
rect 25145 23477 25179 23511
rect 25179 23477 25188 23511
rect 25136 23468 25188 23477
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 7472 23307 7524 23316
rect 7472 23273 7481 23307
rect 7481 23273 7515 23307
rect 7515 23273 7524 23307
rect 7472 23264 7524 23273
rect 8852 23264 8904 23316
rect 15844 23264 15896 23316
rect 16856 23264 16908 23316
rect 17960 23264 18012 23316
rect 18144 23264 18196 23316
rect 19432 23307 19484 23316
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 2136 23060 2188 23112
rect 2596 23128 2648 23180
rect 3056 23128 3108 23180
rect 3700 23060 3752 23112
rect 5080 23128 5132 23180
rect 5356 23128 5408 23180
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 8300 23103 8352 23112
rect 8300 23069 8309 23103
rect 8309 23069 8343 23103
rect 8343 23069 8352 23103
rect 8300 23060 8352 23069
rect 8484 23060 8536 23112
rect 9404 23128 9456 23180
rect 9036 23060 9088 23112
rect 2044 22967 2096 22976
rect 2044 22933 2053 22967
rect 2053 22933 2087 22967
rect 2087 22933 2096 22967
rect 2044 22924 2096 22933
rect 2228 22924 2280 22976
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 2964 22967 3016 22976
rect 2964 22933 2973 22967
rect 2973 22933 3007 22967
rect 3007 22933 3016 22967
rect 2964 22924 3016 22933
rect 3240 22924 3292 22976
rect 5356 22992 5408 23044
rect 9864 23060 9916 23112
rect 10416 23060 10468 23112
rect 11336 23128 11388 23180
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12900 23128 12952 23180
rect 13268 23171 13320 23180
rect 13268 23137 13277 23171
rect 13277 23137 13311 23171
rect 13311 23137 13320 23171
rect 13268 23128 13320 23137
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 19248 23196 19300 23248
rect 18144 23128 18196 23180
rect 19524 23128 19576 23180
rect 17868 23060 17920 23112
rect 19340 23060 19392 23112
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 21088 23196 21140 23248
rect 22744 23264 22796 23316
rect 20536 23128 20588 23180
rect 19708 23060 19760 23069
rect 10048 22992 10100 23044
rect 10876 22992 10928 23044
rect 11888 22992 11940 23044
rect 14556 22992 14608 23044
rect 18696 22992 18748 23044
rect 20996 23060 21048 23112
rect 21916 23103 21968 23112
rect 21916 23069 21925 23103
rect 21925 23069 21959 23103
rect 21959 23069 21968 23103
rect 21916 23060 21968 23069
rect 22284 23060 22336 23112
rect 24584 23128 24636 23180
rect 23204 23103 23256 23112
rect 4988 22924 5040 22976
rect 7748 22924 7800 22976
rect 9128 22924 9180 22976
rect 9312 22924 9364 22976
rect 9404 22924 9456 22976
rect 10324 22967 10376 22976
rect 10324 22933 10333 22967
rect 10333 22933 10367 22967
rect 10367 22933 10376 22967
rect 10324 22924 10376 22933
rect 10784 22924 10836 22976
rect 11152 22924 11204 22976
rect 13452 22924 13504 22976
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 17684 22924 17736 22976
rect 20260 22924 20312 22976
rect 21180 22924 21232 22976
rect 21640 22924 21692 22976
rect 22468 22992 22520 23044
rect 23204 23069 23213 23103
rect 23213 23069 23247 23103
rect 23247 23069 23256 23103
rect 23204 23060 23256 23069
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 23664 22992 23716 23044
rect 24860 23060 24912 23112
rect 25136 22992 25188 23044
rect 25044 22924 25096 22976
rect 25412 22967 25464 22976
rect 25412 22933 25421 22967
rect 25421 22933 25455 22967
rect 25455 22933 25464 22967
rect 25412 22924 25464 22933
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 2412 22720 2464 22772
rect 5724 22720 5776 22772
rect 6276 22720 6328 22772
rect 7472 22720 7524 22772
rect 2044 22652 2096 22704
rect 6644 22652 6696 22704
rect 9036 22720 9088 22772
rect 9128 22763 9180 22772
rect 9128 22729 9137 22763
rect 9137 22729 9171 22763
rect 9171 22729 9180 22763
rect 9128 22720 9180 22729
rect 9404 22720 9456 22772
rect 9588 22720 9640 22772
rect 8576 22652 8628 22704
rect 10600 22652 10652 22704
rect 10968 22695 11020 22704
rect 10968 22661 10977 22695
rect 10977 22661 11011 22695
rect 11011 22661 11020 22695
rect 10968 22652 11020 22661
rect 2228 22584 2280 22636
rect 3056 22584 3108 22636
rect 3516 22627 3568 22636
rect 2780 22516 2832 22568
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 3700 22584 3752 22636
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 6460 22584 6512 22636
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 9220 22584 9272 22593
rect 9312 22627 9364 22636
rect 9312 22593 9321 22627
rect 9321 22593 9355 22627
rect 9355 22593 9364 22627
rect 10140 22627 10192 22636
rect 9312 22584 9364 22593
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 10140 22584 10192 22593
rect 10232 22627 10284 22636
rect 10232 22593 10241 22627
rect 10241 22593 10275 22627
rect 10275 22593 10284 22627
rect 10232 22584 10284 22593
rect 6552 22559 6604 22568
rect 6552 22525 6561 22559
rect 6561 22525 6595 22559
rect 6595 22525 6604 22559
rect 6552 22516 6604 22525
rect 9404 22516 9456 22568
rect 10784 22584 10836 22636
rect 13544 22720 13596 22772
rect 16396 22720 16448 22772
rect 18236 22720 18288 22772
rect 13912 22652 13964 22704
rect 11336 22584 11388 22636
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 13268 22627 13320 22636
rect 11612 22516 11664 22568
rect 13268 22593 13277 22627
rect 13277 22593 13311 22627
rect 13311 22593 13320 22627
rect 13268 22584 13320 22593
rect 13636 22584 13688 22636
rect 14004 22627 14056 22636
rect 14004 22593 14013 22627
rect 14013 22593 14047 22627
rect 14047 22593 14056 22627
rect 14004 22584 14056 22593
rect 16120 22652 16172 22704
rect 18788 22720 18840 22772
rect 19432 22652 19484 22704
rect 15568 22584 15620 22636
rect 17868 22584 17920 22636
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 20996 22720 21048 22772
rect 21272 22720 21324 22772
rect 22560 22720 22612 22772
rect 23388 22720 23440 22772
rect 19708 22652 19760 22704
rect 20536 22652 20588 22704
rect 20628 22652 20680 22704
rect 21180 22652 21232 22704
rect 25412 22652 25464 22704
rect 26056 22652 26108 22704
rect 13360 22516 13412 22568
rect 14924 22559 14976 22568
rect 14924 22525 14933 22559
rect 14933 22525 14967 22559
rect 14967 22525 14976 22559
rect 14924 22516 14976 22525
rect 17408 22516 17460 22568
rect 17684 22516 17736 22568
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 1768 22491 1820 22500
rect 1768 22457 1777 22491
rect 1777 22457 1811 22491
rect 1811 22457 1820 22491
rect 1768 22448 1820 22457
rect 3056 22448 3108 22500
rect 11244 22448 11296 22500
rect 2412 22380 2464 22432
rect 3148 22423 3200 22432
rect 3148 22389 3157 22423
rect 3157 22389 3191 22423
rect 3191 22389 3200 22423
rect 3148 22380 3200 22389
rect 5724 22380 5776 22432
rect 5908 22423 5960 22432
rect 5908 22389 5917 22423
rect 5917 22389 5951 22423
rect 5951 22389 5960 22423
rect 5908 22380 5960 22389
rect 8300 22380 8352 22432
rect 12164 22423 12216 22432
rect 12164 22389 12173 22423
rect 12173 22389 12207 22423
rect 12207 22389 12216 22423
rect 12164 22380 12216 22389
rect 18236 22448 18288 22500
rect 22192 22627 22244 22636
rect 20168 22559 20220 22568
rect 20168 22525 20177 22559
rect 20177 22525 20211 22559
rect 20211 22525 20220 22559
rect 20168 22516 20220 22525
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 21088 22516 21140 22568
rect 23756 22584 23808 22636
rect 23940 22584 23992 22636
rect 24492 22584 24544 22636
rect 25780 22584 25832 22636
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 24860 22516 24912 22568
rect 25596 22516 25648 22568
rect 26240 22516 26292 22568
rect 13912 22380 13964 22432
rect 15292 22380 15344 22432
rect 16304 22423 16356 22432
rect 16304 22389 16313 22423
rect 16313 22389 16347 22423
rect 16347 22389 16356 22423
rect 16304 22380 16356 22389
rect 16764 22380 16816 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 19340 22380 19392 22432
rect 24584 22380 24636 22432
rect 24676 22380 24728 22432
rect 26424 22423 26476 22432
rect 26424 22389 26433 22423
rect 26433 22389 26467 22423
rect 26467 22389 26476 22423
rect 26424 22380 26476 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 8392 22040 8444 22092
rect 9220 22040 9272 22092
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 4804 21972 4856 22024
rect 6552 21972 6604 22024
rect 6736 22015 6788 22024
rect 6736 21981 6770 22015
rect 6770 21981 6788 22015
rect 6736 21972 6788 21981
rect 8576 21972 8628 22024
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 2412 21904 2464 21956
rect 2872 21904 2924 21956
rect 9404 21947 9456 21956
rect 2780 21836 2832 21888
rect 5172 21836 5224 21888
rect 5448 21879 5500 21888
rect 5448 21845 5457 21879
rect 5457 21845 5491 21879
rect 5491 21845 5500 21879
rect 5448 21836 5500 21845
rect 9404 21913 9413 21947
rect 9413 21913 9447 21947
rect 9447 21913 9456 21947
rect 9404 21904 9456 21913
rect 11244 22176 11296 22228
rect 12072 22176 12124 22228
rect 12716 22219 12768 22228
rect 12716 22185 12725 22219
rect 12725 22185 12759 22219
rect 12759 22185 12768 22219
rect 12716 22176 12768 22185
rect 14556 22176 14608 22228
rect 16120 22176 16172 22228
rect 11704 22108 11756 22160
rect 14004 22108 14056 22160
rect 16396 22151 16448 22160
rect 16396 22117 16405 22151
rect 16405 22117 16439 22151
rect 16439 22117 16448 22151
rect 16396 22108 16448 22117
rect 10968 22040 11020 22092
rect 11796 22040 11848 22092
rect 12440 22040 12492 22092
rect 12808 22040 12860 22092
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 13452 21972 13504 22024
rect 13728 21972 13780 22024
rect 14648 22040 14700 22092
rect 18144 22176 18196 22228
rect 19432 22219 19484 22228
rect 19432 22185 19441 22219
rect 19441 22185 19475 22219
rect 19475 22185 19484 22219
rect 19432 22176 19484 22185
rect 19156 22108 19208 22160
rect 19524 22108 19576 22160
rect 19616 22108 19668 22160
rect 20628 22176 20680 22228
rect 21916 22176 21968 22228
rect 22192 22176 22244 22228
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 24860 22176 24912 22228
rect 25044 22176 25096 22228
rect 20260 22108 20312 22160
rect 14740 21972 14792 22024
rect 14924 21972 14976 22024
rect 15292 22015 15344 22024
rect 15292 21981 15326 22015
rect 15326 21981 15344 22015
rect 16856 22015 16908 22024
rect 15292 21972 15344 21981
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 19340 22040 19392 22092
rect 20168 22040 20220 22092
rect 19800 22015 19852 22024
rect 19800 21981 19809 22015
rect 19809 21981 19843 22015
rect 19843 21981 19852 22015
rect 19800 21972 19852 21981
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20536 22015 20588 22024
rect 10416 21904 10468 21956
rect 12532 21904 12584 21956
rect 14096 21904 14148 21956
rect 17868 21904 17920 21956
rect 19340 21904 19392 21956
rect 8852 21836 8904 21888
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 11060 21836 11112 21888
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 12992 21836 13044 21845
rect 14464 21879 14516 21888
rect 14464 21845 14466 21879
rect 14466 21845 14500 21879
rect 14500 21845 14516 21879
rect 14464 21836 14516 21845
rect 17592 21836 17644 21888
rect 20536 21981 20545 22015
rect 20545 21981 20579 22015
rect 20579 21981 20588 22015
rect 20536 21972 20588 21981
rect 20628 21972 20680 22024
rect 20812 21972 20864 22024
rect 21088 21972 21140 22024
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 22100 22108 22152 22160
rect 26424 22108 26476 22160
rect 23572 22040 23624 22092
rect 23940 22040 23992 22092
rect 23664 22015 23716 22024
rect 20352 21904 20404 21956
rect 21916 21904 21968 21956
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 20628 21836 20680 21888
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 25044 22015 25096 22024
rect 25044 21981 25058 22015
rect 25058 21981 25092 22015
rect 25092 21981 25096 22015
rect 25044 21972 25096 21981
rect 25780 21972 25832 22024
rect 26332 21972 26384 22024
rect 24860 21947 24912 21956
rect 24860 21913 24869 21947
rect 24869 21913 24903 21947
rect 24903 21913 24912 21947
rect 24860 21904 24912 21913
rect 25596 21904 25648 21956
rect 24768 21836 24820 21888
rect 27160 21836 27212 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 3424 21632 3476 21684
rect 9312 21675 9364 21684
rect 9312 21641 9321 21675
rect 9321 21641 9355 21675
rect 9355 21641 9364 21675
rect 9312 21632 9364 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11796 21632 11848 21684
rect 14096 21675 14148 21684
rect 14096 21641 14105 21675
rect 14105 21641 14139 21675
rect 14139 21641 14148 21675
rect 14096 21632 14148 21641
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 16304 21632 16356 21684
rect 18236 21632 18288 21684
rect 19800 21632 19852 21684
rect 19892 21632 19944 21684
rect 3516 21564 3568 21616
rect 5080 21564 5132 21616
rect 2136 21496 2188 21548
rect 3056 21496 3108 21548
rect 3700 21496 3752 21548
rect 7104 21496 7156 21548
rect 7380 21539 7432 21548
rect 7012 21428 7064 21480
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 7564 21496 7616 21548
rect 2320 21292 2372 21344
rect 2780 21335 2832 21344
rect 2780 21301 2789 21335
rect 2789 21301 2823 21335
rect 2823 21301 2832 21335
rect 4344 21335 4396 21344
rect 2780 21292 2832 21301
rect 4344 21301 4353 21335
rect 4353 21301 4387 21335
rect 4387 21301 4396 21335
rect 4344 21292 4396 21301
rect 7012 21335 7064 21344
rect 7012 21301 7021 21335
rect 7021 21301 7055 21335
rect 7055 21301 7064 21335
rect 7012 21292 7064 21301
rect 7748 21428 7800 21480
rect 8024 21496 8076 21548
rect 10324 21564 10376 21616
rect 12164 21564 12216 21616
rect 13636 21564 13688 21616
rect 14188 21496 14240 21548
rect 16948 21564 17000 21616
rect 17960 21564 18012 21616
rect 19524 21564 19576 21616
rect 20168 21607 20220 21616
rect 20168 21573 20177 21607
rect 20177 21573 20211 21607
rect 20211 21573 20220 21607
rect 20720 21607 20772 21616
rect 20168 21564 20220 21573
rect 20720 21573 20729 21607
rect 20729 21573 20763 21607
rect 20763 21573 20772 21607
rect 20720 21564 20772 21573
rect 21364 21564 21416 21616
rect 10968 21428 11020 21480
rect 13544 21428 13596 21480
rect 15568 21496 15620 21548
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 15844 21496 15896 21548
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 17408 21496 17460 21548
rect 19432 21496 19484 21548
rect 20628 21539 20680 21548
rect 16672 21428 16724 21480
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 19248 21428 19300 21480
rect 10048 21292 10100 21344
rect 12992 21292 13044 21344
rect 19156 21292 19208 21344
rect 19340 21360 19392 21412
rect 20628 21505 20637 21539
rect 20637 21505 20671 21539
rect 20671 21505 20680 21539
rect 20628 21496 20680 21505
rect 20076 21360 20128 21412
rect 22468 21360 22520 21412
rect 19984 21292 20036 21344
rect 20628 21292 20680 21344
rect 23480 21632 23532 21684
rect 24768 21632 24820 21684
rect 25136 21632 25188 21684
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 23848 21496 23900 21548
rect 24400 21496 24452 21548
rect 25136 21496 25188 21548
rect 23020 21428 23072 21480
rect 24676 21471 24728 21480
rect 24676 21437 24685 21471
rect 24685 21437 24719 21471
rect 24719 21437 24728 21471
rect 24676 21428 24728 21437
rect 23664 21360 23716 21412
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 27252 21496 27304 21548
rect 26240 21403 26292 21412
rect 26240 21369 26249 21403
rect 26249 21369 26283 21403
rect 26283 21369 26292 21403
rect 26240 21360 26292 21369
rect 25596 21292 25648 21344
rect 26332 21292 26384 21344
rect 27712 21292 27764 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 6552 21131 6604 21140
rect 6552 21097 6561 21131
rect 6561 21097 6595 21131
rect 6595 21097 6604 21131
rect 6552 21088 6604 21097
rect 7104 21088 7156 21140
rect 12992 21088 13044 21140
rect 13452 21131 13504 21140
rect 7196 21020 7248 21072
rect 8668 21020 8720 21072
rect 13452 21097 13461 21131
rect 13461 21097 13495 21131
rect 13495 21097 13504 21131
rect 13452 21088 13504 21097
rect 16856 21088 16908 21140
rect 17040 21088 17092 21140
rect 19892 21088 19944 21140
rect 23664 21131 23716 21140
rect 23664 21097 23673 21131
rect 23673 21097 23707 21131
rect 23707 21097 23716 21131
rect 23664 21088 23716 21097
rect 24676 21088 24728 21140
rect 13820 21020 13872 21072
rect 5264 20927 5316 20936
rect 5264 20893 5273 20927
rect 5273 20893 5307 20927
rect 5307 20893 5316 20927
rect 5264 20884 5316 20893
rect 7288 20884 7340 20936
rect 8484 20952 8536 21004
rect 10232 20952 10284 21004
rect 15752 21020 15804 21072
rect 16212 21020 16264 21072
rect 16304 21020 16356 21072
rect 21548 21020 21600 21072
rect 2964 20816 3016 20868
rect 4712 20859 4764 20868
rect 4712 20825 4721 20859
rect 4721 20825 4755 20859
rect 4755 20825 4764 20859
rect 4712 20816 4764 20825
rect 8668 20884 8720 20936
rect 11060 20884 11112 20936
rect 8576 20816 8628 20868
rect 14648 20952 14700 21004
rect 17224 20952 17276 21004
rect 20076 20952 20128 21004
rect 14188 20884 14240 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 18144 20884 18196 20936
rect 18236 20884 18288 20936
rect 20536 20884 20588 20936
rect 21640 20884 21692 20936
rect 23020 20927 23072 20936
rect 23020 20893 23029 20927
rect 23029 20893 23063 20927
rect 23063 20893 23072 20927
rect 23020 20884 23072 20893
rect 23112 20884 23164 20936
rect 23388 20995 23440 21004
rect 23388 20961 23397 20995
rect 23397 20961 23431 20995
rect 23431 20961 23440 20995
rect 23388 20952 23440 20961
rect 23572 20952 23624 21004
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 23480 20927 23532 20936
rect 23480 20893 23489 20927
rect 23489 20893 23523 20927
rect 23523 20893 23532 20927
rect 23480 20884 23532 20893
rect 24860 20884 24912 20936
rect 27160 21088 27212 21140
rect 25596 21020 25648 21072
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 26332 20927 26384 20936
rect 13084 20859 13136 20868
rect 13084 20825 13093 20859
rect 13093 20825 13127 20859
rect 13127 20825 13136 20859
rect 13084 20816 13136 20825
rect 13820 20816 13872 20868
rect 18052 20816 18104 20868
rect 19248 20816 19300 20868
rect 21364 20816 21416 20868
rect 2044 20748 2096 20800
rect 3056 20748 3108 20800
rect 4804 20748 4856 20800
rect 5264 20748 5316 20800
rect 5448 20748 5500 20800
rect 8392 20748 8444 20800
rect 8944 20748 8996 20800
rect 10508 20748 10560 20800
rect 10968 20748 11020 20800
rect 13452 20748 13504 20800
rect 17684 20748 17736 20800
rect 18236 20748 18288 20800
rect 19800 20791 19852 20800
rect 19800 20757 19809 20791
rect 19809 20757 19843 20791
rect 19843 20757 19852 20791
rect 19800 20748 19852 20757
rect 20352 20748 20404 20800
rect 20536 20791 20588 20800
rect 20536 20757 20545 20791
rect 20545 20757 20579 20791
rect 20579 20757 20588 20791
rect 20536 20748 20588 20757
rect 23388 20816 23440 20868
rect 26332 20893 26341 20927
rect 26341 20893 26375 20927
rect 26375 20893 26384 20927
rect 26332 20884 26384 20893
rect 26608 20884 26660 20936
rect 27252 20927 27304 20936
rect 27252 20893 27261 20927
rect 27261 20893 27295 20927
rect 27295 20893 27304 20927
rect 27252 20884 27304 20893
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 27528 20884 27580 20936
rect 28080 20927 28132 20936
rect 28080 20893 28089 20927
rect 28089 20893 28123 20927
rect 28123 20893 28132 20927
rect 28080 20884 28132 20893
rect 23848 20748 23900 20800
rect 27160 20791 27212 20800
rect 27160 20757 27169 20791
rect 27169 20757 27203 20791
rect 27203 20757 27212 20791
rect 27160 20748 27212 20757
rect 27252 20748 27304 20800
rect 27620 20748 27672 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 7656 20544 7708 20596
rect 7840 20544 7892 20596
rect 2688 20519 2740 20528
rect 2688 20485 2697 20519
rect 2697 20485 2731 20519
rect 2731 20485 2740 20519
rect 2688 20476 2740 20485
rect 3332 20476 3384 20528
rect 4160 20476 4212 20528
rect 5540 20476 5592 20528
rect 5724 20476 5776 20528
rect 8484 20544 8536 20596
rect 4896 20408 4948 20460
rect 6460 20408 6512 20460
rect 3056 20340 3108 20392
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 7564 20451 7616 20460
rect 7564 20417 7573 20451
rect 7573 20417 7607 20451
rect 7607 20417 7616 20451
rect 7564 20408 7616 20417
rect 7932 20408 7984 20460
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 9588 20476 9640 20528
rect 10232 20519 10284 20528
rect 10232 20485 10250 20519
rect 10250 20485 10284 20519
rect 10232 20476 10284 20485
rect 8024 20408 8076 20417
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 7656 20340 7708 20392
rect 8944 20340 8996 20392
rect 12624 20544 12676 20596
rect 13176 20544 13228 20596
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 13360 20476 13412 20528
rect 16580 20476 16632 20528
rect 16672 20476 16724 20528
rect 11888 20451 11940 20460
rect 11888 20417 11897 20451
rect 11897 20417 11931 20451
rect 11931 20417 11940 20451
rect 11888 20408 11940 20417
rect 12072 20451 12124 20460
rect 12072 20417 12081 20451
rect 12081 20417 12115 20451
rect 12115 20417 12124 20451
rect 12072 20408 12124 20417
rect 12716 20408 12768 20460
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 15384 20408 15436 20460
rect 15752 20408 15804 20460
rect 16120 20408 16172 20460
rect 19156 20476 19208 20528
rect 23480 20544 23532 20596
rect 23664 20544 23716 20596
rect 24768 20544 24820 20596
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 19616 20408 19668 20460
rect 19892 20451 19944 20460
rect 19892 20417 19901 20451
rect 19901 20417 19935 20451
rect 19935 20417 19944 20451
rect 19892 20408 19944 20417
rect 20444 20408 20496 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20720 20451 20772 20460
rect 20536 20408 20588 20417
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 21548 20408 21600 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 11980 20383 12032 20392
rect 11980 20349 11989 20383
rect 11989 20349 12023 20383
rect 12023 20349 12032 20383
rect 11980 20340 12032 20349
rect 12440 20272 12492 20324
rect 12808 20272 12860 20324
rect 13176 20340 13228 20392
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 14372 20340 14424 20392
rect 14924 20340 14976 20392
rect 20904 20340 20956 20392
rect 23572 20408 23624 20460
rect 24032 20408 24084 20460
rect 24584 20408 24636 20460
rect 27712 20544 27764 20596
rect 27344 20476 27396 20528
rect 23848 20383 23900 20392
rect 23848 20349 23857 20383
rect 23857 20349 23891 20383
rect 23891 20349 23900 20383
rect 23848 20340 23900 20349
rect 26516 20408 26568 20460
rect 26332 20340 26384 20392
rect 13820 20272 13872 20324
rect 15476 20272 15528 20324
rect 17224 20272 17276 20324
rect 20536 20272 20588 20324
rect 21456 20272 21508 20324
rect 21640 20272 21692 20324
rect 27620 20272 27672 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2504 20247 2556 20256
rect 2504 20213 2513 20247
rect 2513 20213 2547 20247
rect 2547 20213 2556 20247
rect 2504 20204 2556 20213
rect 3792 20204 3844 20256
rect 4068 20204 4120 20256
rect 4252 20204 4304 20256
rect 5816 20204 5868 20256
rect 6368 20204 6420 20256
rect 6552 20247 6604 20256
rect 6552 20213 6561 20247
rect 6561 20213 6595 20247
rect 6595 20213 6604 20247
rect 6552 20204 6604 20213
rect 7104 20247 7156 20256
rect 7104 20213 7113 20247
rect 7113 20213 7147 20247
rect 7147 20213 7156 20247
rect 7104 20204 7156 20213
rect 7472 20204 7524 20256
rect 7840 20204 7892 20256
rect 8392 20204 8444 20256
rect 9312 20204 9364 20256
rect 13176 20204 13228 20256
rect 13360 20204 13412 20256
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 18052 20204 18104 20256
rect 19524 20204 19576 20256
rect 22560 20204 22612 20256
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 27068 20204 27120 20256
rect 27988 20247 28040 20256
rect 27988 20213 27997 20247
rect 27997 20213 28031 20247
rect 28031 20213 28040 20247
rect 27988 20204 28040 20213
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 3792 20000 3844 20052
rect 4712 20000 4764 20052
rect 7748 20000 7800 20052
rect 7840 20000 7892 20052
rect 7932 20000 7984 20052
rect 8668 20000 8720 20052
rect 11060 20000 11112 20052
rect 12716 20000 12768 20052
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 16212 20000 16264 20052
rect 17868 20043 17920 20052
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 7288 19932 7340 19984
rect 3608 19864 3660 19916
rect 7748 19864 7800 19916
rect 3148 19796 3200 19848
rect 6552 19796 6604 19848
rect 7196 19796 7248 19848
rect 8116 19932 8168 19984
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 8116 19796 8168 19848
rect 10968 19932 11020 19984
rect 11980 19864 12032 19916
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 2228 19660 2280 19712
rect 4160 19728 4212 19780
rect 4896 19728 4948 19780
rect 5632 19728 5684 19780
rect 6828 19728 6880 19780
rect 7748 19771 7800 19780
rect 7748 19737 7765 19771
rect 7765 19737 7800 19771
rect 7748 19728 7800 19737
rect 8392 19728 8444 19780
rect 8484 19728 8536 19780
rect 11244 19771 11296 19780
rect 11244 19737 11253 19771
rect 11253 19737 11287 19771
rect 11287 19737 11296 19771
rect 11244 19728 11296 19737
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 12624 19839 12676 19848
rect 11796 19796 11848 19805
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 14188 19932 14240 19984
rect 14004 19864 14056 19916
rect 14648 19864 14700 19916
rect 14924 19907 14976 19916
rect 13636 19796 13688 19848
rect 13728 19796 13780 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14924 19873 14933 19907
rect 14933 19873 14967 19907
rect 14967 19873 14976 19907
rect 14924 19864 14976 19873
rect 14556 19796 14608 19805
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16028 19796 16080 19848
rect 17868 20009 17877 20043
rect 17877 20009 17911 20043
rect 17911 20009 17920 20043
rect 17868 20000 17920 20009
rect 19616 20000 19668 20052
rect 20076 20000 20128 20052
rect 23296 20000 23348 20052
rect 20812 19932 20864 19984
rect 21180 19932 21232 19984
rect 22008 19975 22060 19984
rect 22008 19941 22017 19975
rect 22017 19941 22051 19975
rect 22051 19941 22060 19975
rect 22008 19932 22060 19941
rect 7472 19660 7524 19712
rect 7564 19660 7616 19712
rect 10140 19660 10192 19712
rect 13636 19660 13688 19712
rect 14004 19660 14056 19712
rect 14832 19660 14884 19712
rect 20536 19864 20588 19916
rect 21640 19864 21692 19916
rect 23848 20000 23900 20052
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 25596 20000 25648 20052
rect 28080 20000 28132 20052
rect 18420 19796 18472 19848
rect 18512 19796 18564 19848
rect 19432 19796 19484 19848
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 20628 19796 20680 19848
rect 22192 19796 22244 19848
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 19064 19728 19116 19780
rect 20904 19728 20956 19780
rect 23664 19728 23716 19780
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24400 19796 24452 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 24308 19728 24360 19780
rect 24860 19728 24912 19780
rect 25596 19796 25648 19848
rect 27344 19864 27396 19916
rect 27160 19796 27212 19848
rect 26148 19728 26200 19780
rect 27896 19771 27948 19780
rect 18788 19703 18840 19712
rect 18788 19669 18797 19703
rect 18797 19669 18831 19703
rect 18831 19669 18840 19703
rect 19432 19703 19484 19712
rect 18788 19660 18840 19669
rect 19432 19669 19441 19703
rect 19441 19669 19475 19703
rect 19475 19669 19484 19703
rect 19432 19660 19484 19669
rect 21364 19660 21416 19712
rect 23388 19660 23440 19712
rect 23572 19660 23624 19712
rect 27160 19703 27212 19712
rect 27160 19669 27169 19703
rect 27169 19669 27203 19703
rect 27203 19669 27212 19703
rect 27160 19660 27212 19669
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27896 19737 27905 19771
rect 27905 19737 27939 19771
rect 27939 19737 27948 19771
rect 27896 19728 27948 19737
rect 27252 19660 27304 19669
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 3240 19456 3292 19508
rect 6000 19456 6052 19508
rect 8300 19456 8352 19508
rect 9588 19456 9640 19508
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 13176 19456 13228 19508
rect 2872 19388 2924 19440
rect 5356 19431 5408 19440
rect 5356 19397 5365 19431
rect 5365 19397 5399 19431
rect 5399 19397 5408 19431
rect 5356 19388 5408 19397
rect 5448 19431 5500 19440
rect 5448 19397 5457 19431
rect 5457 19397 5491 19431
rect 5491 19397 5500 19431
rect 5448 19388 5500 19397
rect 7012 19388 7064 19440
rect 7656 19388 7708 19440
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 4436 19363 4488 19372
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 4896 19320 4948 19372
rect 5080 19252 5132 19304
rect 5172 19184 5224 19236
rect 6736 19320 6788 19372
rect 7472 19320 7524 19372
rect 8760 19320 8812 19372
rect 9220 19363 9272 19372
rect 9220 19329 9230 19363
rect 9230 19329 9264 19363
rect 9264 19329 9272 19363
rect 10416 19388 10468 19440
rect 15476 19456 15528 19508
rect 19064 19456 19116 19508
rect 21180 19456 21232 19508
rect 24584 19456 24636 19508
rect 15384 19388 15436 19440
rect 9220 19320 9272 19329
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 13452 19320 13504 19372
rect 12532 19252 12584 19304
rect 14004 19320 14056 19372
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 15936 19320 15988 19372
rect 19432 19388 19484 19440
rect 21272 19388 21324 19440
rect 18420 19320 18472 19372
rect 18696 19320 18748 19372
rect 9680 19184 9732 19236
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 19616 19320 19668 19372
rect 21180 19363 21232 19372
rect 13452 19184 13504 19236
rect 4896 19116 4948 19168
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 10048 19116 10100 19168
rect 10508 19116 10560 19168
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 13544 19116 13596 19168
rect 19340 19252 19392 19304
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22560 19388 22612 19440
rect 26056 19456 26108 19508
rect 27528 19499 27580 19508
rect 24860 19388 24912 19440
rect 27528 19465 27537 19499
rect 27537 19465 27571 19499
rect 27571 19465 27580 19499
rect 27528 19456 27580 19465
rect 25044 19320 25096 19372
rect 25872 19363 25924 19372
rect 25872 19329 25881 19363
rect 25881 19329 25915 19363
rect 25915 19329 25924 19363
rect 25872 19320 25924 19329
rect 20812 19252 20864 19304
rect 23020 19252 23072 19304
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 21088 19184 21140 19236
rect 24308 19184 24360 19236
rect 24492 19252 24544 19304
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 27344 19431 27396 19440
rect 27344 19397 27369 19431
rect 27369 19397 27396 19431
rect 27344 19388 27396 19397
rect 26056 19320 26108 19329
rect 27896 19320 27948 19372
rect 26148 19252 26200 19304
rect 25964 19184 26016 19236
rect 14004 19116 14056 19168
rect 14280 19116 14332 19168
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 20536 19116 20588 19168
rect 23572 19116 23624 19168
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 27160 19116 27212 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 5356 18912 5408 18964
rect 7748 18912 7800 18964
rect 13360 18912 13412 18964
rect 13452 18912 13504 18964
rect 14648 18912 14700 18964
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 17960 18912 18012 18964
rect 18696 18912 18748 18964
rect 19892 18912 19944 18964
rect 14556 18844 14608 18896
rect 27344 18912 27396 18964
rect 15844 18776 15896 18828
rect 1584 18708 1636 18760
rect 4160 18708 4212 18760
rect 4804 18708 4856 18760
rect 4988 18751 5040 18760
rect 4988 18717 5022 18751
rect 5022 18717 5040 18751
rect 4988 18708 5040 18717
rect 8484 18708 8536 18760
rect 9496 18708 9548 18760
rect 12716 18708 12768 18760
rect 13636 18708 13688 18760
rect 16580 18708 16632 18760
rect 16856 18708 16908 18760
rect 17224 18708 17276 18760
rect 17960 18708 18012 18760
rect 25044 18844 25096 18896
rect 26332 18844 26384 18896
rect 26516 18844 26568 18896
rect 19800 18776 19852 18828
rect 20720 18819 20772 18828
rect 20720 18785 20729 18819
rect 20729 18785 20763 18819
rect 20763 18785 20772 18819
rect 20720 18776 20772 18785
rect 20904 18776 20956 18828
rect 18696 18708 18748 18760
rect 18880 18708 18932 18760
rect 19892 18751 19944 18760
rect 9864 18683 9916 18692
rect 9864 18649 9898 18683
rect 9898 18649 9916 18683
rect 9864 18640 9916 18649
rect 11980 18683 12032 18692
rect 11980 18649 12014 18683
rect 12014 18649 12032 18683
rect 11980 18640 12032 18649
rect 12992 18640 13044 18692
rect 14280 18683 14332 18692
rect 14280 18649 14289 18683
rect 14289 18649 14323 18683
rect 14323 18649 14332 18683
rect 14280 18640 14332 18649
rect 17500 18683 17552 18692
rect 17500 18649 17509 18683
rect 17509 18649 17543 18683
rect 17543 18649 17552 18683
rect 19892 18717 19901 18751
rect 19901 18717 19935 18751
rect 19935 18717 19944 18751
rect 19892 18708 19944 18717
rect 19984 18751 20036 18760
rect 19984 18717 19993 18751
rect 19993 18717 20027 18751
rect 20027 18717 20036 18751
rect 20812 18751 20864 18760
rect 19984 18708 20036 18717
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 22744 18708 22796 18760
rect 23020 18708 23072 18760
rect 23572 18776 23624 18828
rect 24860 18776 24912 18828
rect 25688 18776 25740 18828
rect 25044 18708 25096 18760
rect 25872 18751 25924 18760
rect 25872 18717 25881 18751
rect 25881 18717 25915 18751
rect 25915 18717 25924 18751
rect 25872 18708 25924 18717
rect 25964 18751 26016 18760
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 26424 18776 26476 18828
rect 25964 18708 26016 18717
rect 26516 18708 26568 18760
rect 17500 18640 17552 18649
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 4068 18615 4120 18624
rect 4068 18581 4077 18615
rect 4077 18581 4111 18615
rect 4111 18581 4120 18615
rect 4068 18572 4120 18581
rect 4712 18572 4764 18624
rect 5172 18572 5224 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 8484 18572 8536 18624
rect 10232 18572 10284 18624
rect 10324 18572 10376 18624
rect 13452 18572 13504 18624
rect 16580 18572 16632 18624
rect 19064 18572 19116 18624
rect 20812 18572 20864 18624
rect 23756 18640 23808 18692
rect 24492 18640 24544 18692
rect 25780 18640 25832 18692
rect 26056 18640 26108 18692
rect 21548 18572 21600 18624
rect 21640 18572 21692 18624
rect 23204 18572 23256 18624
rect 27160 18572 27212 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 5080 18368 5132 18420
rect 4344 18343 4396 18352
rect 4344 18309 4353 18343
rect 4353 18309 4387 18343
rect 4387 18309 4396 18343
rect 4344 18300 4396 18309
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 2228 18232 2280 18284
rect 3884 18232 3936 18284
rect 7104 18300 7156 18352
rect 7656 18368 7708 18420
rect 9220 18368 9272 18420
rect 11980 18368 12032 18420
rect 13360 18368 13412 18420
rect 19892 18368 19944 18420
rect 21548 18368 21600 18420
rect 23572 18411 23624 18420
rect 23572 18377 23581 18411
rect 23581 18377 23615 18411
rect 23615 18377 23624 18411
rect 23572 18368 23624 18377
rect 5080 18275 5132 18284
rect 3240 18164 3292 18216
rect 5080 18241 5089 18275
rect 5089 18241 5123 18275
rect 5123 18241 5132 18275
rect 5080 18232 5132 18241
rect 5356 18232 5408 18284
rect 7748 18232 7800 18284
rect 8484 18232 8536 18284
rect 10232 18300 10284 18352
rect 6736 18207 6788 18216
rect 2504 18096 2556 18148
rect 2228 18028 2280 18080
rect 3332 18096 3384 18148
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 11060 18232 11112 18284
rect 11244 18232 11296 18284
rect 11980 18232 12032 18284
rect 13452 18300 13504 18352
rect 14740 18343 14792 18352
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 15200 18232 15252 18284
rect 8944 18164 8996 18216
rect 9220 18164 9272 18216
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 10508 18164 10560 18216
rect 10876 18164 10928 18216
rect 7932 18096 7984 18148
rect 9036 18096 9088 18148
rect 14096 18164 14148 18216
rect 15844 18232 15896 18284
rect 15752 18164 15804 18216
rect 17868 18232 17920 18284
rect 18144 18232 18196 18284
rect 18880 18275 18932 18284
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 19524 18300 19576 18352
rect 14556 18096 14608 18148
rect 16028 18164 16080 18216
rect 18696 18207 18748 18216
rect 16764 18096 16816 18148
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19340 18164 19392 18216
rect 20168 18232 20220 18284
rect 20720 18164 20772 18216
rect 21088 18232 21140 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 21640 18164 21692 18216
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 23204 18275 23256 18284
rect 22376 18232 22428 18241
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 25044 18232 25096 18284
rect 25964 18232 26016 18284
rect 26332 18232 26384 18284
rect 23756 18207 23808 18216
rect 23756 18173 23765 18207
rect 23765 18173 23799 18207
rect 23799 18173 23808 18207
rect 23756 18164 23808 18173
rect 25596 18207 25648 18216
rect 25596 18173 25605 18207
rect 25605 18173 25639 18207
rect 25639 18173 25648 18207
rect 25596 18164 25648 18173
rect 26240 18207 26292 18216
rect 26240 18173 26249 18207
rect 26249 18173 26283 18207
rect 26283 18173 26292 18207
rect 26240 18164 26292 18173
rect 27252 18207 27304 18216
rect 27252 18173 27261 18207
rect 27261 18173 27295 18207
rect 27295 18173 27304 18207
rect 27252 18164 27304 18173
rect 9404 18028 9456 18080
rect 9772 18028 9824 18080
rect 17868 18028 17920 18080
rect 21180 18028 21232 18080
rect 22284 18096 22336 18148
rect 27896 18096 27948 18148
rect 24308 18071 24360 18080
rect 24308 18037 24317 18071
rect 24317 18037 24351 18071
rect 24351 18037 24360 18071
rect 24308 18028 24360 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 5908 17756 5960 17808
rect 8392 17824 8444 17876
rect 9128 17824 9180 17876
rect 10968 17824 11020 17876
rect 13084 17824 13136 17876
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 15200 17824 15252 17876
rect 18236 17824 18288 17876
rect 21272 17824 21324 17876
rect 2136 17620 2188 17672
rect 2320 17663 2372 17672
rect 2320 17629 2354 17663
rect 2354 17629 2372 17663
rect 2320 17620 2372 17629
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 4344 17663 4396 17672
rect 4344 17629 4353 17663
rect 4353 17629 4387 17663
rect 4387 17629 4396 17663
rect 4344 17620 4396 17629
rect 5356 17620 5408 17672
rect 8576 17756 8628 17808
rect 9864 17756 9916 17808
rect 13176 17756 13228 17808
rect 16672 17756 16724 17808
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 8392 17663 8444 17672
rect 7932 17620 7984 17629
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 5080 17552 5132 17604
rect 7012 17552 7064 17604
rect 7748 17552 7800 17604
rect 8852 17620 8904 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9772 17620 9824 17672
rect 9864 17620 9916 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 4344 17484 4396 17536
rect 6460 17484 6512 17536
rect 7196 17484 7248 17536
rect 8300 17484 8352 17536
rect 10324 17552 10376 17604
rect 16764 17688 16816 17740
rect 17592 17688 17644 17740
rect 17960 17688 18012 17740
rect 11888 17620 11940 17672
rect 13084 17620 13136 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 12164 17552 12216 17604
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 10232 17484 10284 17536
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 12348 17484 12400 17536
rect 13268 17484 13320 17536
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 18972 17688 19024 17740
rect 19524 17756 19576 17808
rect 20444 17756 20496 17808
rect 21364 17756 21416 17808
rect 20536 17688 20588 17740
rect 21272 17688 21324 17740
rect 21456 17688 21508 17740
rect 25688 17824 25740 17876
rect 25964 17867 26016 17876
rect 25964 17833 25973 17867
rect 25973 17833 26007 17867
rect 26007 17833 26016 17867
rect 25964 17824 26016 17833
rect 26424 17824 26476 17876
rect 27252 17824 27304 17876
rect 14556 17620 14608 17629
rect 13820 17552 13872 17604
rect 15292 17595 15344 17604
rect 14004 17484 14056 17536
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 15292 17561 15301 17595
rect 15301 17561 15335 17595
rect 15335 17561 15344 17595
rect 15292 17552 15344 17561
rect 17408 17484 17460 17536
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 18696 17620 18748 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 20076 17620 20128 17672
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 22192 17620 22244 17672
rect 22376 17620 22428 17672
rect 23848 17688 23900 17740
rect 25780 17688 25832 17740
rect 18788 17595 18840 17604
rect 18788 17561 18797 17595
rect 18797 17561 18831 17595
rect 18831 17561 18840 17595
rect 18788 17552 18840 17561
rect 18880 17595 18932 17604
rect 18880 17561 18889 17595
rect 18889 17561 18923 17595
rect 18923 17561 18932 17595
rect 18880 17552 18932 17561
rect 19156 17552 19208 17604
rect 20536 17552 20588 17604
rect 22284 17552 22336 17604
rect 23388 17663 23440 17672
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 24768 17663 24820 17672
rect 23756 17552 23808 17604
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 26240 17620 26292 17672
rect 27160 17663 27212 17672
rect 27160 17629 27169 17663
rect 27169 17629 27203 17663
rect 27203 17629 27212 17663
rect 27160 17620 27212 17629
rect 24860 17552 24912 17604
rect 19524 17484 19576 17536
rect 20352 17484 20404 17536
rect 21548 17484 21600 17536
rect 22468 17527 22520 17536
rect 22468 17493 22477 17527
rect 22477 17493 22511 17527
rect 22511 17493 22520 17527
rect 22468 17484 22520 17493
rect 22836 17527 22888 17536
rect 22836 17493 22845 17527
rect 22845 17493 22879 17527
rect 22879 17493 22888 17527
rect 22836 17484 22888 17493
rect 23572 17527 23624 17536
rect 23572 17493 23581 17527
rect 23581 17493 23615 17527
rect 23615 17493 23624 17527
rect 23572 17484 23624 17493
rect 23940 17484 23992 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 8392 17280 8444 17332
rect 2780 17212 2832 17264
rect 5632 17212 5684 17264
rect 6460 17212 6512 17264
rect 11704 17280 11756 17332
rect 4712 17144 4764 17196
rect 4896 17187 4948 17196
rect 4896 17153 4930 17187
rect 4930 17153 4948 17187
rect 4896 17144 4948 17153
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 6828 17187 6880 17196
rect 2136 17119 2188 17128
rect 2136 17085 2145 17119
rect 2145 17085 2179 17119
rect 2179 17085 2188 17119
rect 2136 17076 2188 17085
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7656 17144 7708 17196
rect 7748 17144 7800 17196
rect 9312 17144 9364 17196
rect 9956 17144 10008 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10784 17212 10836 17264
rect 12164 17255 12216 17264
rect 12164 17221 12173 17255
rect 12173 17221 12207 17255
rect 12207 17221 12216 17255
rect 12164 17212 12216 17221
rect 3516 17051 3568 17060
rect 3516 17017 3525 17051
rect 3525 17017 3559 17051
rect 3559 17017 3568 17051
rect 3516 17008 3568 17017
rect 6000 17051 6052 17060
rect 6000 17017 6009 17051
rect 6009 17017 6043 17051
rect 6043 17017 6052 17051
rect 6000 17008 6052 17017
rect 7288 17008 7340 17060
rect 9128 17051 9180 17060
rect 9128 17017 9137 17051
rect 9137 17017 9171 17051
rect 9171 17017 9180 17051
rect 9128 17008 9180 17017
rect 9680 17008 9732 17060
rect 10416 17008 10468 17060
rect 10784 17008 10836 17060
rect 5356 16940 5408 16992
rect 9404 16940 9456 16992
rect 10600 16940 10652 16992
rect 12256 17187 12308 17196
rect 13912 17280 13964 17332
rect 13176 17212 13228 17264
rect 12256 17153 12273 17187
rect 12273 17153 12307 17187
rect 12307 17153 12308 17187
rect 12256 17144 12308 17153
rect 13544 17144 13596 17196
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 19248 17280 19300 17332
rect 20352 17280 20404 17332
rect 19616 17212 19668 17264
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 16212 17144 16264 17196
rect 16764 17144 16816 17196
rect 19892 17144 19944 17196
rect 20076 17187 20128 17196
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 21272 17212 21324 17264
rect 21456 17212 21508 17264
rect 22192 17323 22244 17332
rect 22192 17289 22217 17323
rect 22217 17289 22244 17323
rect 22192 17280 22244 17289
rect 22836 17280 22888 17332
rect 22652 17212 22704 17264
rect 24768 17212 24820 17264
rect 21640 17144 21692 17196
rect 21732 17144 21784 17196
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 24860 17144 24912 17196
rect 27344 17144 27396 17196
rect 27896 17187 27948 17196
rect 27896 17153 27905 17187
rect 27905 17153 27939 17187
rect 27939 17153 27948 17187
rect 27896 17144 27948 17153
rect 16028 17076 16080 17128
rect 16672 17076 16724 17128
rect 19340 17076 19392 17128
rect 19800 17076 19852 17128
rect 21364 17076 21416 17128
rect 23388 17076 23440 17128
rect 15200 17008 15252 17060
rect 21456 17008 21508 17060
rect 12164 16940 12216 16992
rect 17224 16940 17276 16992
rect 18236 16983 18288 16992
rect 18236 16949 18245 16983
rect 18245 16949 18279 16983
rect 18279 16949 18288 16983
rect 18236 16940 18288 16949
rect 20812 16940 20864 16992
rect 21180 16983 21232 16992
rect 21180 16949 21189 16983
rect 21189 16949 21223 16983
rect 21223 16949 21232 16983
rect 21180 16940 21232 16949
rect 21732 16940 21784 16992
rect 22284 17008 22336 17060
rect 22744 17008 22796 17060
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 23756 17119 23808 17128
rect 23756 17085 23765 17119
rect 23765 17085 23799 17119
rect 23799 17085 23808 17119
rect 23756 17076 23808 17085
rect 24952 17008 25004 17060
rect 24768 16940 24820 16992
rect 25688 16983 25740 16992
rect 25688 16949 25697 16983
rect 25697 16949 25731 16983
rect 25731 16949 25740 16983
rect 25688 16940 25740 16949
rect 27068 16940 27120 16992
rect 27620 16940 27672 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 5724 16736 5776 16788
rect 8760 16736 8812 16788
rect 10232 16736 10284 16788
rect 5264 16668 5316 16720
rect 3516 16600 3568 16652
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 7472 16600 7524 16652
rect 2688 16464 2740 16516
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 4436 16464 4488 16516
rect 6736 16532 6788 16584
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 7748 16464 7800 16516
rect 8576 16532 8628 16584
rect 10140 16532 10192 16584
rect 12348 16736 12400 16788
rect 14004 16736 14056 16788
rect 16212 16736 16264 16788
rect 16948 16736 17000 16788
rect 13636 16668 13688 16720
rect 16396 16668 16448 16720
rect 18236 16736 18288 16788
rect 18696 16736 18748 16788
rect 21364 16779 21416 16788
rect 21364 16745 21373 16779
rect 21373 16745 21407 16779
rect 21407 16745 21416 16779
rect 21364 16736 21416 16745
rect 24308 16736 24360 16788
rect 27804 16779 27856 16788
rect 27804 16745 27813 16779
rect 27813 16745 27847 16779
rect 27847 16745 27856 16779
rect 27804 16736 27856 16745
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 15200 16600 15252 16652
rect 16672 16600 16724 16652
rect 21088 16668 21140 16720
rect 21272 16668 21324 16720
rect 12624 16532 12676 16584
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 8484 16464 8536 16516
rect 10048 16464 10100 16516
rect 4344 16396 4396 16448
rect 6552 16396 6604 16448
rect 8300 16396 8352 16448
rect 8944 16396 8996 16448
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 13360 16507 13412 16516
rect 13360 16473 13369 16507
rect 13369 16473 13403 16507
rect 13403 16473 13412 16507
rect 13544 16507 13596 16516
rect 13360 16464 13412 16473
rect 13544 16473 13553 16507
rect 13553 16473 13587 16507
rect 13587 16473 13596 16507
rect 13544 16464 13596 16473
rect 14740 16464 14792 16516
rect 16580 16532 16632 16584
rect 17224 16532 17276 16584
rect 20260 16600 20312 16652
rect 19800 16532 19852 16584
rect 21548 16600 21600 16652
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20720 16575 20772 16584
rect 20536 16532 20588 16541
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 20812 16532 20864 16584
rect 21640 16575 21692 16584
rect 18236 16464 18288 16516
rect 21180 16464 21232 16516
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 22468 16600 22520 16652
rect 25688 16668 25740 16720
rect 25596 16643 25648 16652
rect 25596 16609 25605 16643
rect 25605 16609 25639 16643
rect 25639 16609 25648 16643
rect 25596 16600 25648 16609
rect 22376 16575 22428 16584
rect 22376 16541 22385 16575
rect 22385 16541 22419 16575
rect 22419 16541 22428 16575
rect 22376 16532 22428 16541
rect 22560 16532 22612 16584
rect 23388 16532 23440 16584
rect 23480 16532 23532 16584
rect 23940 16532 23992 16584
rect 24768 16532 24820 16584
rect 25780 16532 25832 16584
rect 15292 16396 15344 16448
rect 17500 16396 17552 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 20076 16396 20128 16448
rect 20628 16439 20680 16448
rect 20628 16405 20637 16439
rect 20637 16405 20671 16439
rect 20671 16405 20680 16439
rect 20628 16396 20680 16405
rect 20996 16396 21048 16448
rect 22744 16396 22796 16448
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 23572 16396 23624 16448
rect 24952 16464 25004 16516
rect 27160 16532 27212 16584
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 27436 16532 27488 16584
rect 26700 16507 26752 16516
rect 26700 16473 26709 16507
rect 26709 16473 26743 16507
rect 26743 16473 26752 16507
rect 26700 16464 26752 16473
rect 26056 16396 26108 16448
rect 26976 16439 27028 16448
rect 26976 16405 26985 16439
rect 26985 16405 27019 16439
rect 27019 16405 27028 16439
rect 26976 16396 27028 16405
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 2136 16192 2188 16244
rect 6828 16192 6880 16244
rect 2964 16124 3016 16176
rect 7380 16124 7432 16176
rect 7748 16192 7800 16244
rect 12440 16192 12492 16244
rect 12716 16192 12768 16244
rect 16764 16192 16816 16244
rect 16948 16235 17000 16244
rect 16948 16201 16957 16235
rect 16957 16201 16991 16235
rect 16991 16201 17000 16235
rect 16948 16192 17000 16201
rect 21640 16192 21692 16244
rect 23112 16192 23164 16244
rect 9496 16124 9548 16176
rect 10416 16167 10468 16176
rect 10416 16133 10425 16167
rect 10425 16133 10459 16167
rect 10459 16133 10468 16167
rect 10416 16124 10468 16133
rect 11152 16124 11204 16176
rect 13360 16124 13412 16176
rect 13912 16124 13964 16176
rect 16396 16124 16448 16176
rect 17408 16124 17460 16176
rect 21548 16124 21600 16176
rect 22560 16124 22612 16176
rect 22744 16167 22796 16176
rect 22744 16133 22753 16167
rect 22753 16133 22787 16167
rect 22787 16133 22796 16167
rect 22744 16124 22796 16133
rect 3792 16056 3844 16108
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 7840 16099 7892 16108
rect 6552 15920 6604 15972
rect 6736 15920 6788 15972
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 10324 16099 10376 16108
rect 10324 16065 10331 16099
rect 10331 16065 10376 16099
rect 10324 16056 10376 16065
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 10784 16056 10836 16108
rect 11060 16056 11112 16108
rect 11796 16056 11848 16108
rect 15016 16056 15068 16108
rect 15844 16056 15896 16108
rect 16120 16056 16172 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 9956 15988 10008 16040
rect 14004 15988 14056 16040
rect 14832 15988 14884 16040
rect 15568 15988 15620 16040
rect 10140 15920 10192 15972
rect 10600 15920 10652 15972
rect 4896 15852 4948 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 11244 15852 11296 15904
rect 17040 15920 17092 15972
rect 17224 16056 17276 16108
rect 18696 16099 18748 16108
rect 17868 15988 17920 16040
rect 18144 15988 18196 16040
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 20260 16056 20312 16108
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 27436 16192 27488 16244
rect 27620 16192 27672 16244
rect 24768 16124 24820 16176
rect 19800 16031 19852 16040
rect 19800 15997 19809 16031
rect 19809 15997 19843 16031
rect 19843 15997 19852 16031
rect 19800 15988 19852 15997
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 20720 15988 20772 16040
rect 21548 15988 21600 16040
rect 22376 15988 22428 16040
rect 23664 16056 23716 16108
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 25596 16124 25648 16176
rect 25688 16056 25740 16108
rect 25964 16124 26016 16176
rect 26608 16124 26660 16176
rect 22836 15988 22888 16040
rect 23848 15988 23900 16040
rect 20904 15920 20956 15972
rect 21640 15920 21692 15972
rect 24860 16031 24912 16040
rect 24860 15997 24869 16031
rect 24869 15997 24903 16031
rect 24903 15997 24912 16031
rect 24860 15988 24912 15997
rect 25964 15988 26016 16040
rect 26700 16056 26752 16108
rect 27712 16031 27764 16040
rect 27712 15997 27721 16031
rect 27721 15997 27755 16031
rect 27755 15997 27764 16031
rect 27712 15988 27764 15997
rect 28080 15920 28132 15972
rect 13544 15852 13596 15904
rect 14096 15852 14148 15904
rect 15844 15852 15896 15904
rect 19340 15852 19392 15904
rect 19708 15852 19760 15904
rect 22560 15852 22612 15904
rect 22928 15852 22980 15904
rect 24952 15852 25004 15904
rect 25780 15852 25832 15904
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 2044 15691 2096 15700
rect 2044 15657 2053 15691
rect 2053 15657 2087 15691
rect 2087 15657 2096 15691
rect 2044 15648 2096 15657
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 12624 15648 12676 15700
rect 14832 15648 14884 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 7748 15580 7800 15632
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 4804 15512 4856 15564
rect 6644 15512 6696 15564
rect 9496 15580 9548 15632
rect 20628 15648 20680 15700
rect 21180 15648 21232 15700
rect 19708 15623 19760 15632
rect 4988 15444 5040 15496
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 7104 15444 7156 15496
rect 8024 15487 8076 15496
rect 8024 15453 8031 15487
rect 8031 15453 8076 15487
rect 8024 15444 8076 15453
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 10692 15512 10744 15564
rect 3332 15419 3384 15428
rect 3332 15385 3341 15419
rect 3341 15385 3375 15419
rect 3375 15385 3384 15419
rect 3332 15376 3384 15385
rect 5448 15376 5500 15428
rect 5264 15308 5316 15360
rect 8944 15376 8996 15428
rect 12808 15444 12860 15496
rect 9496 15419 9548 15428
rect 9496 15385 9505 15419
rect 9505 15385 9539 15419
rect 9539 15385 9548 15419
rect 9496 15376 9548 15385
rect 11060 15376 11112 15428
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 15016 15444 15068 15496
rect 13360 15376 13412 15428
rect 16304 15444 16356 15496
rect 18052 15444 18104 15496
rect 18512 15512 18564 15564
rect 19432 15555 19484 15564
rect 19432 15521 19441 15555
rect 19441 15521 19475 15555
rect 19475 15521 19484 15555
rect 19432 15512 19484 15521
rect 19708 15589 19717 15623
rect 19717 15589 19751 15623
rect 19751 15589 19760 15623
rect 19708 15580 19760 15589
rect 25136 15648 25188 15700
rect 25688 15648 25740 15700
rect 20076 15512 20128 15564
rect 22468 15580 22520 15632
rect 23388 15580 23440 15632
rect 21548 15512 21600 15564
rect 22744 15512 22796 15564
rect 23480 15555 23532 15564
rect 23480 15521 23489 15555
rect 23489 15521 23523 15555
rect 23523 15521 23532 15555
rect 23480 15512 23532 15521
rect 17684 15376 17736 15428
rect 18236 15376 18288 15428
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20352 15444 20404 15453
rect 20628 15444 20680 15496
rect 21272 15444 21324 15496
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 25596 15580 25648 15632
rect 23848 15444 23900 15496
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 25596 15444 25648 15496
rect 25780 15487 25832 15496
rect 25780 15453 25789 15487
rect 25789 15453 25823 15487
rect 25823 15453 25832 15487
rect 25780 15444 25832 15453
rect 26976 15648 27028 15700
rect 27712 15648 27764 15700
rect 28080 15691 28132 15700
rect 28080 15657 28089 15691
rect 28089 15657 28123 15691
rect 28123 15657 28132 15691
rect 28080 15648 28132 15657
rect 27344 15555 27396 15564
rect 27344 15521 27353 15555
rect 27353 15521 27387 15555
rect 27387 15521 27396 15555
rect 27344 15512 27396 15521
rect 27620 15512 27672 15564
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 18788 15376 18840 15428
rect 21548 15419 21600 15428
rect 21548 15385 21557 15419
rect 21557 15385 21591 15419
rect 21591 15385 21600 15419
rect 21548 15376 21600 15385
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 9680 15308 9732 15360
rect 12532 15308 12584 15360
rect 12992 15308 13044 15360
rect 13728 15308 13780 15360
rect 15568 15308 15620 15360
rect 18880 15308 18932 15360
rect 19524 15308 19576 15360
rect 20812 15308 20864 15360
rect 23572 15308 23624 15360
rect 23940 15308 23992 15360
rect 26056 15308 26108 15360
rect 27988 15444 28040 15496
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 5448 15104 5500 15156
rect 4068 15079 4120 15088
rect 4068 15045 4077 15079
rect 4077 15045 4111 15079
rect 4111 15045 4120 15079
rect 4068 15036 4120 15045
rect 5080 15036 5132 15088
rect 6736 15104 6788 15156
rect 4712 14968 4764 15020
rect 5264 14968 5316 15020
rect 5816 14968 5868 15020
rect 9036 15104 9088 15156
rect 9772 15104 9824 15156
rect 11980 15104 12032 15156
rect 12164 15104 12216 15156
rect 12624 15104 12676 15156
rect 10968 15079 11020 15088
rect 10968 15045 10977 15079
rect 10977 15045 11011 15079
rect 11011 15045 11020 15079
rect 10968 15036 11020 15045
rect 12348 15036 12400 15088
rect 14096 15036 14148 15088
rect 16120 15104 16172 15156
rect 20076 15147 20128 15156
rect 7104 14968 7156 15020
rect 8484 14968 8536 15020
rect 1768 14832 1820 14884
rect 3332 14764 3384 14816
rect 8576 14900 8628 14952
rect 11152 14968 11204 15020
rect 12532 14968 12584 15020
rect 12992 14968 13044 15020
rect 13544 14968 13596 15020
rect 14924 14968 14976 15020
rect 15568 15011 15620 15020
rect 11704 14943 11756 14952
rect 9128 14832 9180 14884
rect 10140 14832 10192 14884
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 13452 14900 13504 14952
rect 13820 14900 13872 14952
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 16948 14968 17000 15020
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 17132 14968 17184 15020
rect 18236 15036 18288 15088
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 20076 15113 20085 15147
rect 20085 15113 20119 15147
rect 20119 15113 20128 15147
rect 20076 15104 20128 15113
rect 20444 15104 20496 15156
rect 20628 15104 20680 15156
rect 20720 15104 20772 15156
rect 22376 15104 22428 15156
rect 22008 15036 22060 15088
rect 23664 15104 23716 15156
rect 25596 15147 25648 15156
rect 25596 15113 25605 15147
rect 25605 15113 25639 15147
rect 25639 15113 25648 15147
rect 25596 15104 25648 15113
rect 27344 15147 27396 15156
rect 27344 15113 27353 15147
rect 27353 15113 27387 15147
rect 27387 15113 27396 15147
rect 27344 15104 27396 15113
rect 23480 15036 23532 15088
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20076 14968 20128 15020
rect 20352 14968 20404 15020
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 21456 15011 21508 15020
rect 21456 14977 21465 15011
rect 21465 14977 21499 15011
rect 21499 14977 21508 15011
rect 21456 14968 21508 14977
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 22744 14968 22796 15020
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24768 15036 24820 15088
rect 25688 15079 25740 15088
rect 25688 15045 25697 15079
rect 25697 15045 25731 15079
rect 25731 15045 25740 15079
rect 25688 15036 25740 15045
rect 25964 15036 26016 15088
rect 26976 15036 27028 15088
rect 26608 14968 26660 15020
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 19248 14943 19300 14952
rect 14280 14832 14332 14884
rect 14372 14832 14424 14884
rect 14648 14832 14700 14884
rect 17868 14832 17920 14884
rect 18512 14875 18564 14884
rect 18512 14841 18521 14875
rect 18521 14841 18555 14875
rect 18555 14841 18564 14875
rect 18512 14832 18564 14841
rect 18788 14832 18840 14884
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 19340 14900 19392 14952
rect 20260 14900 20312 14952
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 21088 14832 21140 14884
rect 22836 14875 22888 14884
rect 22836 14841 22845 14875
rect 22845 14841 22879 14875
rect 22879 14841 22888 14875
rect 22836 14832 22888 14841
rect 13728 14764 13780 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 14556 14764 14608 14816
rect 14924 14764 14976 14816
rect 15476 14764 15528 14816
rect 15752 14764 15804 14816
rect 16764 14764 16816 14816
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 18236 14764 18288 14816
rect 20076 14764 20128 14816
rect 20904 14764 20956 14816
rect 22192 14764 22244 14816
rect 22928 14764 22980 14816
rect 23388 14764 23440 14816
rect 24584 14807 24636 14816
rect 24584 14773 24593 14807
rect 24593 14773 24627 14807
rect 24627 14773 24636 14807
rect 24584 14764 24636 14773
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1860 14560 1912 14612
rect 3240 14560 3292 14612
rect 11244 14560 11296 14612
rect 11980 14560 12032 14612
rect 16948 14560 17000 14612
rect 17776 14560 17828 14612
rect 18604 14560 18656 14612
rect 18788 14560 18840 14612
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 24308 14560 24360 14612
rect 24584 14560 24636 14612
rect 5264 14492 5316 14544
rect 2044 14467 2096 14476
rect 2044 14433 2053 14467
rect 2053 14433 2087 14467
rect 2087 14433 2096 14467
rect 2044 14424 2096 14433
rect 5448 14424 5500 14476
rect 7104 14424 7156 14476
rect 9404 14424 9456 14476
rect 2320 14399 2372 14408
rect 2320 14365 2354 14399
rect 2354 14365 2372 14399
rect 4252 14399 4304 14408
rect 2320 14356 2372 14365
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 5356 14356 5408 14408
rect 6368 14356 6420 14408
rect 8300 14356 8352 14408
rect 8484 14356 8536 14408
rect 8944 14356 8996 14408
rect 10876 14492 10928 14544
rect 12900 14492 12952 14544
rect 15752 14492 15804 14544
rect 18420 14492 18472 14544
rect 19064 14492 19116 14544
rect 20076 14492 20128 14544
rect 23664 14492 23716 14544
rect 13544 14424 13596 14476
rect 12348 14356 12400 14408
rect 13084 14356 13136 14408
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 14280 14399 14332 14408
rect 13268 14356 13320 14365
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 16856 14424 16908 14476
rect 14740 14356 14792 14408
rect 15568 14356 15620 14408
rect 15752 14356 15804 14408
rect 18144 14424 18196 14476
rect 22468 14424 22520 14476
rect 4896 14288 4948 14340
rect 5080 14288 5132 14340
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 18880 14356 18932 14408
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20720 14356 20772 14408
rect 21088 14399 21140 14408
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 8668 14220 8720 14272
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 9588 14288 9640 14340
rect 12900 14288 12952 14340
rect 13728 14288 13780 14340
rect 10324 14220 10376 14272
rect 10416 14220 10468 14272
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 16488 14288 16540 14340
rect 18052 14288 18104 14340
rect 18144 14288 18196 14340
rect 18328 14288 18380 14340
rect 18696 14288 18748 14340
rect 20444 14331 20496 14340
rect 17224 14220 17276 14272
rect 18236 14220 18288 14272
rect 18788 14263 18840 14272
rect 18788 14229 18797 14263
rect 18797 14229 18831 14263
rect 18831 14229 18840 14263
rect 18788 14220 18840 14229
rect 20444 14297 20453 14331
rect 20453 14297 20487 14331
rect 20487 14297 20496 14331
rect 20444 14288 20496 14297
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 21548 14356 21600 14408
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 21640 14220 21692 14272
rect 22008 14288 22060 14340
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 24952 14356 25004 14408
rect 24400 14288 24452 14340
rect 22928 14263 22980 14272
rect 22928 14229 22937 14263
rect 22937 14229 22971 14263
rect 22971 14229 22980 14263
rect 22928 14220 22980 14229
rect 24492 14220 24544 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 1768 14016 1820 14068
rect 5816 14016 5868 14068
rect 7288 14059 7340 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2228 13880 2280 13932
rect 5540 13948 5592 14000
rect 1860 13744 1912 13796
rect 3424 13812 3476 13864
rect 6460 13880 6512 13932
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10692 14016 10744 14068
rect 12440 14016 12492 14068
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13360 14016 13412 14068
rect 14648 14059 14700 14068
rect 11244 13948 11296 14000
rect 12808 13948 12860 14000
rect 14004 13948 14056 14000
rect 6184 13812 6236 13864
rect 3792 13787 3844 13796
rect 3792 13753 3801 13787
rect 3801 13753 3835 13787
rect 3835 13753 3844 13787
rect 3792 13744 3844 13753
rect 6460 13744 6512 13796
rect 7288 13880 7340 13932
rect 7748 13880 7800 13932
rect 8300 13880 8352 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 10692 13880 10744 13932
rect 10876 13880 10928 13932
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 8484 13812 8536 13864
rect 8944 13812 8996 13864
rect 10784 13812 10836 13864
rect 11704 13855 11756 13864
rect 9036 13744 9088 13796
rect 3056 13676 3108 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 8576 13676 8628 13728
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 15660 14016 15712 14068
rect 15936 14016 15988 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 17224 14016 17276 14068
rect 17132 13948 17184 14000
rect 17684 13991 17736 14000
rect 17684 13957 17693 13991
rect 17693 13957 17727 13991
rect 17727 13957 17736 13991
rect 17684 13948 17736 13957
rect 20720 14016 20772 14068
rect 20536 13948 20588 14000
rect 20628 13948 20680 14000
rect 13728 13880 13780 13889
rect 14096 13812 14148 13864
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 15292 13880 15344 13932
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16028 13923 16080 13932
rect 16028 13889 16042 13923
rect 16042 13889 16076 13923
rect 16076 13889 16080 13923
rect 16028 13880 16080 13889
rect 12808 13744 12860 13796
rect 13912 13744 13964 13796
rect 11980 13676 12032 13728
rect 14188 13676 14240 13728
rect 15936 13744 15988 13796
rect 16120 13812 16172 13864
rect 17316 13880 17368 13932
rect 18696 13923 18748 13932
rect 16304 13812 16356 13864
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 19892 13880 19944 13932
rect 22468 13923 22520 13932
rect 19708 13812 19760 13864
rect 20720 13812 20772 13864
rect 22468 13889 22477 13923
rect 22477 13889 22511 13923
rect 22511 13889 22520 13923
rect 22468 13880 22520 13889
rect 22928 13880 22980 13932
rect 16948 13744 17000 13796
rect 17224 13744 17276 13796
rect 20352 13744 20404 13796
rect 24584 13880 24636 13932
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25596 13880 25648 13932
rect 14648 13676 14700 13728
rect 15476 13676 15528 13728
rect 20168 13676 20220 13728
rect 21456 13676 21508 13728
rect 23112 13676 23164 13728
rect 24952 13676 25004 13728
rect 25136 13719 25188 13728
rect 25136 13685 25145 13719
rect 25145 13685 25179 13719
rect 25179 13685 25188 13719
rect 25136 13676 25188 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 2780 13472 2832 13524
rect 3976 13472 4028 13524
rect 6552 13472 6604 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12532 13472 12584 13524
rect 13820 13472 13872 13524
rect 14464 13472 14516 13524
rect 16580 13472 16632 13524
rect 20904 13472 20956 13524
rect 14740 13404 14792 13456
rect 19616 13404 19668 13456
rect 19984 13404 20036 13456
rect 20444 13404 20496 13456
rect 9036 13336 9088 13388
rect 1860 13268 1912 13320
rect 4528 13268 4580 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 4804 13268 4856 13320
rect 7196 13268 7248 13320
rect 8300 13268 8352 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 2136 13200 2188 13252
rect 5816 13200 5868 13252
rect 6276 13200 6328 13252
rect 9404 13336 9456 13388
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10968 13268 11020 13320
rect 13268 13268 13320 13320
rect 16580 13336 16632 13388
rect 19708 13379 19760 13388
rect 19708 13345 19717 13379
rect 19717 13345 19751 13379
rect 19751 13345 19760 13379
rect 19708 13336 19760 13345
rect 20720 13336 20772 13388
rect 3700 13132 3752 13184
rect 5356 13132 5408 13184
rect 5908 13132 5960 13184
rect 10232 13200 10284 13252
rect 12164 13200 12216 13252
rect 14464 13268 14516 13320
rect 13912 13200 13964 13252
rect 14280 13200 14332 13252
rect 11888 13132 11940 13184
rect 12624 13132 12676 13184
rect 13084 13132 13136 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 15752 13268 15804 13320
rect 18236 13268 18288 13320
rect 16304 13200 16356 13252
rect 20260 13268 20312 13320
rect 24400 13472 24452 13524
rect 25044 13404 25096 13456
rect 20352 13200 20404 13252
rect 19432 13132 19484 13184
rect 19984 13175 20036 13184
rect 19984 13141 19993 13175
rect 19993 13141 20027 13175
rect 20027 13141 20036 13175
rect 19984 13132 20036 13141
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 25872 13336 25924 13388
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 23112 13268 23164 13320
rect 23204 13200 23256 13252
rect 25320 13268 25372 13320
rect 25596 13311 25648 13320
rect 25596 13277 25605 13311
rect 25605 13277 25639 13311
rect 25639 13277 25648 13311
rect 25596 13268 25648 13277
rect 25964 13311 26016 13320
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 20812 13132 20864 13184
rect 21548 13132 21600 13184
rect 25136 13200 25188 13252
rect 25688 13132 25740 13184
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 4252 12928 4304 12980
rect 4712 12928 4764 12980
rect 4160 12792 4212 12844
rect 7380 12928 7432 12980
rect 9312 12928 9364 12980
rect 4712 12792 4764 12844
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 5080 12792 5132 12844
rect 5448 12792 5500 12844
rect 5724 12792 5776 12844
rect 6460 12860 6512 12912
rect 10416 12928 10468 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 19432 12971 19484 12980
rect 6092 12792 6144 12844
rect 5632 12699 5684 12708
rect 4436 12588 4488 12640
rect 5080 12588 5132 12640
rect 5632 12665 5641 12699
rect 5641 12665 5675 12699
rect 5675 12665 5684 12699
rect 5632 12656 5684 12665
rect 5724 12588 5776 12640
rect 6000 12588 6052 12640
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7288 12835 7340 12844
rect 7288 12801 7296 12835
rect 7296 12801 7330 12835
rect 7330 12801 7340 12835
rect 7288 12792 7340 12801
rect 7564 12792 7616 12844
rect 8668 12792 8720 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10416 12835 10468 12844
rect 10232 12792 10284 12801
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10692 12792 10744 12844
rect 11704 12860 11756 12912
rect 13176 12860 13228 12912
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 7656 12724 7708 12776
rect 14004 12792 14056 12844
rect 14096 12792 14148 12844
rect 15568 12860 15620 12912
rect 15292 12792 15344 12844
rect 16304 12903 16356 12912
rect 16304 12869 16313 12903
rect 16313 12869 16347 12903
rect 16347 12869 16356 12903
rect 16304 12860 16356 12869
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20720 12928 20772 12980
rect 23204 12971 23256 12980
rect 23204 12937 23213 12971
rect 23213 12937 23247 12971
rect 23247 12937 23256 12971
rect 23204 12928 23256 12937
rect 18052 12903 18104 12912
rect 18052 12869 18061 12903
rect 18061 12869 18095 12903
rect 18095 12869 18104 12903
rect 18052 12860 18104 12869
rect 18144 12860 18196 12912
rect 17684 12835 17736 12844
rect 7472 12656 7524 12708
rect 6828 12588 6880 12640
rect 8484 12588 8536 12640
rect 9036 12588 9088 12640
rect 12624 12724 12676 12776
rect 15476 12724 15528 12776
rect 14556 12656 14608 12708
rect 16764 12724 16816 12776
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 18236 12792 18288 12844
rect 22376 12860 22428 12912
rect 19248 12835 19300 12844
rect 19248 12801 19279 12835
rect 19279 12801 19300 12835
rect 19248 12792 19300 12801
rect 20536 12792 20588 12844
rect 20720 12792 20772 12844
rect 21272 12792 21324 12844
rect 21456 12792 21508 12844
rect 17960 12724 18012 12776
rect 22560 12792 22612 12844
rect 22744 12792 22796 12844
rect 25320 12928 25372 12980
rect 26056 12928 26108 12980
rect 25964 12860 26016 12912
rect 12808 12588 12860 12640
rect 16672 12656 16724 12708
rect 21456 12656 21508 12708
rect 22560 12656 22612 12708
rect 23664 12835 23716 12844
rect 23664 12801 23699 12835
rect 23699 12801 23716 12835
rect 24492 12835 24544 12844
rect 23664 12792 23716 12801
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 24768 12792 24820 12844
rect 25780 12792 25832 12844
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 24400 12767 24452 12776
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 25596 12724 25648 12776
rect 25688 12767 25740 12776
rect 25688 12733 25697 12767
rect 25697 12733 25731 12767
rect 25731 12733 25740 12767
rect 25688 12724 25740 12733
rect 25228 12656 25280 12708
rect 25964 12656 26016 12708
rect 16580 12588 16632 12640
rect 18052 12588 18104 12640
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 19340 12588 19392 12640
rect 20996 12588 21048 12640
rect 24952 12588 25004 12640
rect 25044 12588 25096 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 2412 12384 2464 12436
rect 6644 12384 6696 12436
rect 9128 12384 9180 12436
rect 11244 12384 11296 12436
rect 11888 12384 11940 12436
rect 12072 12384 12124 12436
rect 12716 12384 12768 12436
rect 14464 12384 14516 12436
rect 5540 12180 5592 12232
rect 3700 12112 3752 12164
rect 3976 12155 4028 12164
rect 3976 12121 3985 12155
rect 3985 12121 4019 12155
rect 4019 12121 4028 12155
rect 3976 12112 4028 12121
rect 4068 12112 4120 12164
rect 6828 12180 6880 12232
rect 8668 12316 8720 12368
rect 17592 12384 17644 12436
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 20720 12384 20772 12436
rect 22376 12427 22428 12436
rect 22376 12393 22385 12427
rect 22385 12393 22419 12427
rect 22419 12393 22428 12427
rect 22376 12384 22428 12393
rect 23848 12384 23900 12436
rect 20444 12316 20496 12368
rect 10416 12248 10468 12300
rect 15660 12291 15712 12300
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 8944 12180 8996 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9496 12180 9548 12232
rect 9680 12180 9732 12232
rect 10692 12180 10744 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 7564 12112 7616 12164
rect 6920 12044 6972 12096
rect 7196 12044 7248 12096
rect 8484 12112 8536 12164
rect 10416 12112 10468 12164
rect 9036 12044 9088 12096
rect 9496 12044 9548 12096
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16028 12248 16080 12300
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 14096 12180 14148 12232
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15292 12180 15344 12232
rect 14188 12112 14240 12164
rect 16764 12180 16816 12232
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 15752 12112 15804 12164
rect 14464 12044 14516 12096
rect 17224 12112 17276 12164
rect 18144 12112 18196 12164
rect 20260 12180 20312 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21272 12180 21324 12232
rect 21456 12180 21508 12232
rect 24124 12248 24176 12300
rect 23112 12223 23164 12232
rect 23112 12189 23121 12223
rect 23121 12189 23155 12223
rect 23155 12189 23164 12223
rect 23112 12180 23164 12189
rect 25044 12316 25096 12368
rect 25412 12316 25464 12368
rect 24768 12248 24820 12300
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25044 12223 25096 12232
rect 25044 12189 25053 12223
rect 25053 12189 25087 12223
rect 25087 12189 25096 12223
rect 25044 12180 25096 12189
rect 25412 12180 25464 12232
rect 25964 12223 26016 12232
rect 17776 12044 17828 12096
rect 18236 12044 18288 12096
rect 18972 12044 19024 12096
rect 23296 12112 23348 12164
rect 24584 12155 24636 12164
rect 24584 12121 24593 12155
rect 24593 12121 24627 12155
rect 24627 12121 24636 12155
rect 24584 12112 24636 12121
rect 24676 12155 24728 12164
rect 24676 12121 24685 12155
rect 24685 12121 24719 12155
rect 24719 12121 24728 12155
rect 24676 12112 24728 12121
rect 25136 12112 25188 12164
rect 25596 12112 25648 12164
rect 25964 12189 25973 12223
rect 25973 12189 26007 12223
rect 26007 12189 26016 12223
rect 25964 12180 26016 12189
rect 20536 12044 20588 12096
rect 22652 12044 22704 12096
rect 23388 12044 23440 12096
rect 25228 12087 25280 12096
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 25228 12044 25280 12053
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 2228 11840 2280 11892
rect 3516 11840 3568 11892
rect 6552 11840 6604 11892
rect 7012 11840 7064 11892
rect 8668 11840 8720 11892
rect 9220 11840 9272 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 3792 11772 3844 11824
rect 5356 11772 5408 11824
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2872 11747 2924 11756
rect 2872 11713 2906 11747
rect 2906 11713 2924 11747
rect 2872 11704 2924 11713
rect 5632 11704 5684 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 2044 11636 2096 11688
rect 4344 11636 4396 11688
rect 6368 11636 6420 11688
rect 8300 11704 8352 11756
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 6276 11500 6328 11552
rect 7564 11500 7616 11552
rect 9036 11636 9088 11688
rect 8668 11500 8720 11552
rect 9496 11772 9548 11824
rect 12164 11815 12216 11824
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 12164 11781 12173 11815
rect 12173 11781 12207 11815
rect 12207 11781 12216 11815
rect 12164 11772 12216 11781
rect 19432 11840 19484 11892
rect 22192 11840 22244 11892
rect 22836 11840 22888 11892
rect 14188 11772 14240 11824
rect 15568 11772 15620 11824
rect 16028 11772 16080 11824
rect 17408 11772 17460 11824
rect 18144 11772 18196 11824
rect 10048 11704 10100 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 12716 11636 12768 11688
rect 14648 11636 14700 11688
rect 15752 11636 15804 11688
rect 16856 11679 16908 11688
rect 16856 11645 16865 11679
rect 16865 11645 16899 11679
rect 16899 11645 16908 11679
rect 16856 11636 16908 11645
rect 18788 11772 18840 11824
rect 19800 11815 19852 11824
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 19800 11781 19809 11815
rect 19809 11781 19843 11815
rect 19843 11781 19852 11815
rect 19800 11772 19852 11781
rect 19984 11772 20036 11824
rect 19892 11704 19944 11756
rect 25228 11772 25280 11824
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22468 11704 22520 11756
rect 23480 11704 23532 11756
rect 25964 11840 26016 11892
rect 26056 11704 26108 11756
rect 21364 11636 21416 11688
rect 22100 11636 22152 11688
rect 24860 11636 24912 11688
rect 25872 11636 25924 11688
rect 10508 11500 10560 11552
rect 10784 11500 10836 11552
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 12072 11500 12124 11552
rect 17776 11500 17828 11552
rect 19984 11568 20036 11620
rect 20812 11611 20864 11620
rect 20812 11577 20821 11611
rect 20821 11577 20855 11611
rect 20855 11577 20864 11611
rect 20812 11568 20864 11577
rect 22744 11568 22796 11620
rect 24400 11568 24452 11620
rect 18696 11500 18748 11552
rect 20076 11500 20128 11552
rect 22192 11500 22244 11552
rect 23664 11500 23716 11552
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 6184 11296 6236 11348
rect 11336 11296 11388 11348
rect 10784 11228 10836 11280
rect 8576 11160 8628 11212
rect 14556 11296 14608 11348
rect 16856 11296 16908 11348
rect 14004 11228 14056 11280
rect 19616 11296 19668 11348
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 20260 11296 20312 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 24676 11296 24728 11348
rect 24860 11296 24912 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 13176 11160 13228 11212
rect 15292 11160 15344 11212
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 11060 11092 11112 11144
rect 17960 11160 18012 11212
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 18052 11092 18104 11144
rect 23112 11160 23164 11212
rect 4712 11024 4764 11076
rect 6736 11024 6788 11076
rect 5264 10956 5316 11008
rect 6552 10956 6604 11008
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 8208 10956 8260 11008
rect 8392 10956 8444 11008
rect 8668 11024 8720 11076
rect 9864 11024 9916 11076
rect 10784 11024 10836 11076
rect 10508 10956 10560 11008
rect 14648 11024 14700 11076
rect 17960 11024 18012 11076
rect 19156 11024 19208 11076
rect 19248 11024 19300 11076
rect 19800 11024 19852 11076
rect 20260 11092 20312 11144
rect 21272 11092 21324 11144
rect 21456 11092 21508 11144
rect 22100 11092 22152 11144
rect 23572 11160 23624 11212
rect 24308 11160 24360 11212
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 24400 11092 24452 11144
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 25136 11092 25188 11144
rect 25688 11092 25740 11144
rect 25872 11092 25924 11144
rect 19432 10956 19484 11008
rect 20168 10956 20220 11008
rect 20720 10956 20772 11008
rect 21456 10956 21508 11008
rect 22284 10999 22336 11008
rect 22284 10965 22293 10999
rect 22293 10965 22327 10999
rect 22327 10965 22336 10999
rect 22284 10956 22336 10965
rect 23756 10999 23808 11008
rect 23756 10965 23765 10999
rect 23765 10965 23799 10999
rect 23799 10965 23808 10999
rect 23756 10956 23808 10965
rect 24216 11024 24268 11076
rect 25136 10956 25188 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 4344 10752 4396 10804
rect 4712 10752 4764 10804
rect 4896 10752 4948 10804
rect 5448 10752 5500 10804
rect 5724 10752 5776 10804
rect 5908 10795 5960 10804
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 7288 10752 7340 10804
rect 7380 10752 7432 10804
rect 9772 10752 9824 10804
rect 12716 10752 12768 10804
rect 2780 10684 2832 10736
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 3608 10616 3660 10668
rect 5080 10659 5132 10668
rect 3884 10548 3936 10600
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 7472 10684 7524 10736
rect 10968 10684 11020 10736
rect 11244 10684 11296 10736
rect 11336 10684 11388 10736
rect 17408 10752 17460 10804
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 6828 10659 6880 10668
rect 5356 10548 5408 10600
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 8852 10616 8904 10668
rect 9036 10616 9088 10668
rect 10508 10616 10560 10668
rect 11888 10616 11940 10668
rect 12072 10616 12124 10668
rect 12164 10616 12216 10668
rect 18880 10616 18932 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19892 10752 19944 10804
rect 20904 10752 20956 10804
rect 21088 10752 21140 10804
rect 21548 10752 21600 10804
rect 21824 10752 21876 10804
rect 10048 10548 10100 10600
rect 15292 10548 15344 10600
rect 16672 10548 16724 10600
rect 11980 10480 12032 10532
rect 20536 10616 20588 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 22928 10684 22980 10736
rect 24124 10684 24176 10736
rect 24584 10752 24636 10804
rect 26148 10684 26200 10736
rect 21088 10616 21140 10625
rect 22376 10616 22428 10668
rect 23296 10616 23348 10668
rect 20996 10548 21048 10600
rect 23756 10548 23808 10600
rect 24676 10616 24728 10668
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 24584 10548 24636 10600
rect 22284 10480 22336 10532
rect 22652 10480 22704 10532
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 7380 10412 7432 10464
rect 10508 10412 10560 10464
rect 13912 10412 13964 10464
rect 17960 10412 18012 10464
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 19524 10412 19576 10464
rect 20260 10412 20312 10464
rect 21180 10412 21232 10464
rect 21548 10412 21600 10464
rect 23664 10480 23716 10532
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2688 10208 2740 10260
rect 5540 10208 5592 10260
rect 9588 10208 9640 10260
rect 9680 10208 9732 10260
rect 12072 10208 12124 10260
rect 12164 10208 12216 10260
rect 16672 10251 16724 10260
rect 8024 10140 8076 10192
rect 8300 10140 8352 10192
rect 10416 10140 10468 10192
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4160 10004 4212 10056
rect 6368 10072 6420 10124
rect 6552 10072 6604 10124
rect 5264 10047 5316 10056
rect 4252 9936 4304 9988
rect 1676 9868 1728 9920
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 10600 10072 10652 10124
rect 8024 10004 8076 10056
rect 8944 10004 8996 10056
rect 7104 9936 7156 9988
rect 7380 9936 7432 9988
rect 7564 9936 7616 9988
rect 9772 9979 9824 9988
rect 9772 9945 9781 9979
rect 9781 9945 9815 9979
rect 9815 9945 9824 9979
rect 9772 9936 9824 9945
rect 5080 9868 5132 9920
rect 6828 9868 6880 9920
rect 9588 9868 9640 9920
rect 13912 10004 13964 10056
rect 13820 9936 13872 9988
rect 12808 9868 12860 9920
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 21548 10208 21600 10260
rect 21732 10208 21784 10260
rect 22652 10208 22704 10260
rect 17408 10140 17460 10192
rect 15200 10072 15252 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 17040 10004 17092 10056
rect 23112 10140 23164 10192
rect 24676 10208 24728 10260
rect 25136 10208 25188 10260
rect 26148 10208 26200 10260
rect 25872 10140 25924 10192
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 23480 10072 23532 10124
rect 14740 9936 14792 9988
rect 18696 9936 18748 9988
rect 20168 9979 20220 9988
rect 20168 9945 20177 9979
rect 20177 9945 20211 9979
rect 20211 9945 20220 9979
rect 20168 9936 20220 9945
rect 16028 9868 16080 9920
rect 16672 9868 16724 9920
rect 19800 9868 19852 9920
rect 20260 9868 20312 9920
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 21180 10047 21232 10056
rect 20904 10004 20956 10013
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 20996 9936 21048 9988
rect 21640 9936 21692 9988
rect 22836 10004 22888 10056
rect 23388 10004 23440 10056
rect 24860 10004 24912 10056
rect 22468 9936 22520 9988
rect 23940 9936 23992 9988
rect 24768 9979 24820 9988
rect 22192 9868 22244 9920
rect 22376 9868 22428 9920
rect 23388 9868 23440 9920
rect 24768 9945 24795 9979
rect 24795 9945 24820 9979
rect 24768 9936 24820 9945
rect 25044 9936 25096 9988
rect 24124 9868 24176 9920
rect 25596 9911 25648 9920
rect 25596 9877 25605 9911
rect 25605 9877 25639 9911
rect 25639 9877 25648 9911
rect 25596 9868 25648 9877
rect 26240 9911 26292 9920
rect 26240 9877 26249 9911
rect 26249 9877 26283 9911
rect 26283 9877 26292 9911
rect 26240 9868 26292 9877
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 1952 9664 2004 9716
rect 6828 9664 6880 9716
rect 4712 9596 4764 9648
rect 5172 9596 5224 9648
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 3332 9528 3384 9580
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 6092 9596 6144 9648
rect 6368 9596 6420 9648
rect 13820 9664 13872 9716
rect 17224 9664 17276 9716
rect 17868 9664 17920 9716
rect 18052 9664 18104 9716
rect 6460 9528 6512 9580
rect 9404 9596 9456 9648
rect 11704 9596 11756 9648
rect 4068 9392 4120 9444
rect 5724 9392 5776 9444
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 6092 9460 6144 9512
rect 7656 9460 7708 9512
rect 10968 9528 11020 9580
rect 12164 9528 12216 9580
rect 14372 9596 14424 9648
rect 19800 9664 19852 9716
rect 21548 9664 21600 9716
rect 21640 9664 21692 9716
rect 13176 9528 13228 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13728 9528 13780 9580
rect 10232 9460 10284 9512
rect 11612 9460 11664 9512
rect 15844 9503 15896 9512
rect 7196 9324 7248 9376
rect 9404 9324 9456 9376
rect 11060 9324 11112 9376
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 11980 9324 12032 9333
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 17776 9528 17828 9580
rect 18604 9528 18656 9580
rect 19064 9596 19116 9648
rect 19156 9596 19208 9648
rect 22652 9596 22704 9648
rect 24676 9664 24728 9716
rect 25044 9664 25096 9716
rect 25872 9664 25924 9716
rect 24124 9596 24176 9648
rect 18972 9528 19024 9580
rect 22560 9528 22612 9580
rect 15016 9392 15068 9444
rect 21088 9460 21140 9512
rect 22284 9503 22336 9512
rect 13176 9324 13228 9376
rect 16396 9324 16448 9376
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18144 9324 18196 9376
rect 19892 9392 19944 9444
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 22928 9528 22980 9580
rect 23112 9571 23164 9580
rect 23112 9537 23121 9571
rect 23121 9537 23155 9571
rect 23155 9537 23164 9571
rect 23112 9528 23164 9537
rect 23480 9460 23532 9512
rect 22744 9392 22796 9444
rect 22836 9392 22888 9444
rect 23204 9392 23256 9444
rect 24032 9528 24084 9580
rect 24584 9571 24636 9580
rect 24584 9537 24593 9571
rect 24593 9537 24627 9571
rect 24627 9537 24636 9571
rect 24584 9528 24636 9537
rect 24676 9571 24728 9580
rect 24676 9537 24685 9571
rect 24685 9537 24719 9571
rect 24719 9537 24728 9571
rect 24676 9528 24728 9537
rect 25136 9528 25188 9580
rect 23940 9460 23992 9512
rect 24768 9460 24820 9512
rect 20076 9324 20128 9376
rect 21088 9324 21140 9376
rect 21824 9324 21876 9376
rect 22192 9324 22244 9376
rect 22652 9324 22704 9376
rect 24124 9392 24176 9444
rect 23480 9324 23532 9376
rect 23848 9324 23900 9376
rect 24952 9392 25004 9444
rect 26240 9460 26292 9512
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 2872 9120 2924 9172
rect 4896 9163 4948 9172
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 5264 9120 5316 9172
rect 7012 9120 7064 9172
rect 7288 9120 7340 9172
rect 7656 9120 7708 9172
rect 10324 9120 10376 9172
rect 12992 9120 13044 9172
rect 15844 9120 15896 9172
rect 18880 9120 18932 9172
rect 19156 9120 19208 9172
rect 20904 9120 20956 9172
rect 22284 9120 22336 9172
rect 22744 9120 22796 9172
rect 23204 9120 23256 9172
rect 24676 9120 24728 9172
rect 25596 9120 25648 9172
rect 3976 9052 4028 9104
rect 2964 8984 3016 9036
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 4252 8984 4304 9036
rect 5448 9052 5500 9104
rect 18144 9052 18196 9104
rect 18788 9052 18840 9104
rect 19248 9052 19300 9104
rect 1952 8848 2004 8900
rect 2688 8848 2740 8900
rect 3700 8916 3752 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4804 8984 4856 9036
rect 2412 8780 2464 8832
rect 3516 8780 3568 8832
rect 3608 8780 3660 8832
rect 5172 8916 5224 8968
rect 5816 8916 5868 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 7104 8984 7156 9036
rect 8576 8984 8628 9036
rect 6184 8848 6236 8900
rect 6644 8916 6696 8968
rect 7564 8916 7616 8968
rect 5724 8780 5776 8832
rect 6644 8780 6696 8832
rect 7472 8848 7524 8900
rect 8760 8916 8812 8968
rect 10692 8984 10744 9036
rect 11060 9027 11112 9036
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11060 8984 11112 8993
rect 13544 8984 13596 9036
rect 15752 8984 15804 9036
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17592 8984 17644 9036
rect 10876 8916 10928 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 20260 8916 20312 8968
rect 21732 9052 21784 9104
rect 21824 9052 21876 9104
rect 22560 9052 22612 9104
rect 23388 9052 23440 9104
rect 21456 8984 21508 9036
rect 11244 8848 11296 8900
rect 11980 8848 12032 8900
rect 13728 8891 13780 8900
rect 7656 8780 7708 8832
rect 7748 8780 7800 8832
rect 9128 8780 9180 8832
rect 10600 8780 10652 8832
rect 12900 8780 12952 8832
rect 13728 8857 13737 8891
rect 13737 8857 13771 8891
rect 13771 8857 13780 8891
rect 13728 8848 13780 8857
rect 15016 8848 15068 8900
rect 15936 8848 15988 8900
rect 15384 8780 15436 8832
rect 15476 8780 15528 8832
rect 17132 8848 17184 8900
rect 19340 8780 19392 8832
rect 19616 8780 19668 8832
rect 19984 8848 20036 8900
rect 22100 8959 22152 8968
rect 22100 8925 22109 8959
rect 22109 8925 22143 8959
rect 22143 8925 22152 8959
rect 23388 8959 23440 8968
rect 22100 8916 22152 8925
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 24768 9052 24820 9104
rect 23848 9027 23900 9036
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 24032 8984 24084 9036
rect 23480 8916 23532 8925
rect 21088 8848 21140 8900
rect 21364 8848 21416 8900
rect 24860 8848 24912 8900
rect 22652 8780 22704 8832
rect 23204 8823 23256 8832
rect 23204 8789 23213 8823
rect 23213 8789 23247 8823
rect 23247 8789 23256 8823
rect 23204 8780 23256 8789
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1676 8576 1728 8628
rect 5264 8576 5316 8628
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 5908 8619 5960 8628
rect 5908 8585 5917 8619
rect 5917 8585 5951 8619
rect 5951 8585 5960 8619
rect 5908 8576 5960 8585
rect 6000 8576 6052 8628
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 1952 8551 2004 8560
rect 1952 8517 1961 8551
rect 1961 8517 1995 8551
rect 1995 8517 2004 8551
rect 1952 8508 2004 8517
rect 3056 8551 3108 8560
rect 3056 8517 3065 8551
rect 3065 8517 3099 8551
rect 3099 8517 3108 8551
rect 3056 8508 3108 8517
rect 3424 8551 3476 8560
rect 3424 8517 3433 8551
rect 3433 8517 3467 8551
rect 3467 8517 3476 8551
rect 3424 8508 3476 8517
rect 5448 8508 5500 8560
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3608 8440 3660 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 5908 8440 5960 8492
rect 7104 8440 7156 8492
rect 7656 8440 7708 8492
rect 12900 8576 12952 8628
rect 9680 8508 9732 8560
rect 14648 8576 14700 8628
rect 15936 8576 15988 8628
rect 16028 8576 16080 8628
rect 17132 8576 17184 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17776 8619 17828 8628
rect 17408 8576 17460 8585
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 19892 8576 19944 8628
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 13912 8508 13964 8560
rect 15108 8508 15160 8560
rect 18972 8508 19024 8560
rect 19064 8508 19116 8560
rect 22192 8619 22244 8628
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 24124 8619 24176 8628
rect 24124 8585 24133 8619
rect 24133 8585 24167 8619
rect 24167 8585 24176 8619
rect 24124 8576 24176 8585
rect 7564 8415 7616 8424
rect 2504 8347 2556 8356
rect 2504 8313 2513 8347
rect 2513 8313 2547 8347
rect 2547 8313 2556 8347
rect 2504 8304 2556 8313
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8300 8372 8352 8424
rect 11152 8415 11204 8424
rect 11152 8381 11161 8415
rect 11161 8381 11195 8415
rect 11195 8381 11204 8415
rect 11152 8372 11204 8381
rect 15476 8440 15528 8492
rect 13268 8372 13320 8424
rect 15660 8415 15712 8424
rect 15660 8381 15669 8415
rect 15669 8381 15703 8415
rect 15703 8381 15712 8415
rect 15660 8372 15712 8381
rect 18052 8440 18104 8492
rect 16580 8372 16632 8424
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 9312 8304 9364 8356
rect 9404 8304 9456 8356
rect 10692 8304 10744 8356
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 18328 8440 18380 8492
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 23204 8508 23256 8560
rect 20628 8440 20680 8492
rect 21180 8440 21232 8492
rect 21640 8440 21692 8492
rect 22836 8440 22888 8492
rect 24768 8440 24820 8492
rect 20720 8372 20772 8424
rect 24584 8372 24636 8424
rect 25136 8415 25188 8424
rect 25136 8381 25145 8415
rect 25145 8381 25179 8415
rect 25179 8381 25188 8415
rect 25136 8372 25188 8381
rect 13452 8304 13504 8313
rect 19340 8304 19392 8356
rect 21180 8304 21232 8356
rect 4804 8236 4856 8288
rect 5540 8236 5592 8288
rect 7288 8236 7340 8288
rect 9864 8236 9916 8288
rect 16856 8236 16908 8288
rect 17132 8236 17184 8288
rect 19156 8236 19208 8288
rect 19892 8279 19944 8288
rect 19892 8245 19901 8279
rect 19901 8245 19935 8279
rect 19935 8245 19944 8279
rect 19892 8236 19944 8245
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 21456 8236 21508 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 2964 8032 3016 8084
rect 3332 8032 3384 8084
rect 6092 8032 6144 8084
rect 7380 8032 7432 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 4344 7964 4396 8016
rect 7196 7964 7248 8016
rect 10048 7964 10100 8016
rect 11244 8032 11296 8084
rect 12256 8032 12308 8084
rect 14648 8032 14700 8084
rect 12900 7964 12952 8016
rect 13636 7964 13688 8016
rect 17132 7964 17184 8016
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 5724 7896 5776 7948
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 4252 7828 4304 7880
rect 5356 7828 5408 7880
rect 7196 7828 7248 7880
rect 7472 7828 7524 7880
rect 4068 7760 4120 7812
rect 4896 7760 4948 7812
rect 10600 7896 10652 7948
rect 9128 7828 9180 7880
rect 9312 7803 9364 7812
rect 9312 7769 9321 7803
rect 9321 7769 9355 7803
rect 9355 7769 9364 7803
rect 9312 7760 9364 7769
rect 9864 7828 9916 7880
rect 11060 7828 11112 7880
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 9220 7692 9272 7744
rect 11980 7896 12032 7948
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12624 7896 12676 7948
rect 12992 7896 13044 7948
rect 14372 7896 14424 7948
rect 15108 7896 15160 7948
rect 12164 7828 12216 7837
rect 14648 7828 14700 7880
rect 17960 7964 18012 8016
rect 18236 8032 18288 8084
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 18144 7964 18196 8016
rect 19248 7964 19300 8016
rect 19340 7964 19392 8016
rect 19432 7896 19484 7948
rect 18696 7871 18748 7880
rect 12716 7692 12768 7744
rect 13452 7692 13504 7744
rect 16672 7760 16724 7812
rect 16764 7760 16816 7812
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18788 7828 18840 7880
rect 23388 8032 23440 8084
rect 24124 8032 24176 8084
rect 20720 7896 20772 7948
rect 21272 7964 21324 8016
rect 24216 7964 24268 8016
rect 18236 7760 18288 7812
rect 21180 7871 21232 7880
rect 19432 7803 19484 7812
rect 19432 7769 19441 7803
rect 19441 7769 19475 7803
rect 19475 7769 19484 7803
rect 19432 7760 19484 7769
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21088 7760 21140 7812
rect 21548 7828 21600 7880
rect 23296 7896 23348 7948
rect 20996 7692 21048 7744
rect 22284 7803 22336 7812
rect 22284 7769 22293 7803
rect 22293 7769 22327 7803
rect 22327 7769 22336 7803
rect 22284 7760 22336 7769
rect 22652 7760 22704 7812
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1768 7488 1820 7540
rect 4160 7488 4212 7540
rect 4988 7488 5040 7540
rect 6736 7488 6788 7540
rect 7104 7488 7156 7540
rect 7472 7488 7524 7540
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 9404 7488 9456 7540
rect 10968 7488 11020 7540
rect 12624 7488 12676 7540
rect 4344 7420 4396 7472
rect 7380 7463 7432 7472
rect 7380 7429 7389 7463
rect 7389 7429 7423 7463
rect 7423 7429 7432 7463
rect 7380 7420 7432 7429
rect 4896 7352 4948 7404
rect 5632 7352 5684 7404
rect 7104 7352 7156 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7748 7352 7800 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9864 7352 9916 7404
rect 10048 7395 10100 7404
rect 10048 7361 10082 7395
rect 10082 7361 10100 7395
rect 10048 7352 10100 7361
rect 11796 7420 11848 7472
rect 10968 7352 11020 7404
rect 16488 7488 16540 7540
rect 16856 7488 16908 7540
rect 17408 7488 17460 7540
rect 14004 7420 14056 7472
rect 19432 7488 19484 7540
rect 23572 7488 23624 7540
rect 19064 7420 19116 7472
rect 22284 7420 22336 7472
rect 9588 7284 9640 7336
rect 12164 7284 12216 7336
rect 12440 7284 12492 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 8484 7148 8536 7200
rect 9680 7216 9732 7268
rect 12900 7259 12952 7268
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 19892 7352 19944 7404
rect 22560 7352 22612 7404
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 13728 7216 13780 7268
rect 15292 7284 15344 7336
rect 17132 7327 17184 7336
rect 16672 7216 16724 7268
rect 14096 7148 14148 7200
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 17500 7284 17552 7336
rect 17132 7148 17184 7200
rect 18696 7148 18748 7200
rect 21548 7216 21600 7268
rect 22744 7148 22796 7200
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 7104 6944 7156 6996
rect 7472 6944 7524 6996
rect 7748 6944 7800 6996
rect 9680 6944 9732 6996
rect 4804 6876 4856 6928
rect 8300 6876 8352 6928
rect 2504 6808 2556 6860
rect 3884 6808 3936 6860
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5816 6808 5868 6860
rect 11888 6944 11940 6996
rect 12624 6944 12676 6996
rect 16580 6919 16632 6928
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 6644 6740 6696 6792
rect 7564 6740 7616 6792
rect 8484 6740 8536 6792
rect 9588 6740 9640 6792
rect 9772 6740 9824 6792
rect 2688 6672 2740 6724
rect 7380 6672 7432 6724
rect 3332 6604 3384 6656
rect 7196 6604 7248 6656
rect 8668 6672 8720 6724
rect 10692 6740 10744 6792
rect 13268 6740 13320 6792
rect 14096 6808 14148 6860
rect 16580 6885 16589 6919
rect 16589 6885 16623 6919
rect 16623 6885 16632 6919
rect 16580 6876 16632 6885
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 15936 6740 15988 6792
rect 16856 6740 16908 6792
rect 10048 6672 10100 6724
rect 11428 6672 11480 6724
rect 14556 6715 14608 6724
rect 14556 6681 14565 6715
rect 14565 6681 14599 6715
rect 14599 6681 14608 6715
rect 14556 6672 14608 6681
rect 16764 6672 16816 6724
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 19340 6672 19392 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 20812 6672 20864 6724
rect 20720 6604 20772 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 5448 6443 5500 6452
rect 3332 6400 3384 6409
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 7748 6400 7800 6452
rect 8300 6400 8352 6452
rect 12440 6400 12492 6452
rect 4344 6375 4396 6384
rect 4344 6341 4353 6375
rect 4353 6341 4387 6375
rect 4387 6341 4396 6375
rect 4344 6332 4396 6341
rect 8392 6332 8444 6384
rect 2688 6264 2740 6316
rect 3608 6264 3660 6316
rect 7472 6264 7524 6316
rect 8668 6264 8720 6316
rect 9312 6264 9364 6316
rect 9588 6264 9640 6316
rect 11428 6332 11480 6384
rect 11704 6375 11756 6384
rect 11704 6341 11713 6375
rect 11713 6341 11747 6375
rect 11747 6341 11756 6375
rect 11704 6332 11756 6341
rect 14648 6400 14700 6452
rect 15016 6400 15068 6452
rect 18144 6400 18196 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 20904 6400 20956 6452
rect 6644 6196 6696 6248
rect 11060 6264 11112 6316
rect 13820 6332 13872 6384
rect 12716 6264 12768 6316
rect 14832 6264 14884 6316
rect 4160 6128 4212 6180
rect 7288 6128 7340 6180
rect 14280 6196 14332 6248
rect 16764 6332 16816 6384
rect 16948 6332 17000 6384
rect 15936 6307 15988 6316
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 16028 6264 16080 6316
rect 18236 6264 18288 6316
rect 18880 6332 18932 6384
rect 19064 6332 19116 6384
rect 20444 6332 20496 6384
rect 20812 6375 20864 6384
rect 20812 6341 20821 6375
rect 20821 6341 20855 6375
rect 20855 6341 20864 6375
rect 20812 6332 20864 6341
rect 18696 6264 18748 6316
rect 2872 6060 2924 6112
rect 3608 6060 3660 6112
rect 5172 6060 5224 6112
rect 5816 6060 5868 6112
rect 13636 6128 13688 6180
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16672 6196 16724 6248
rect 17224 6196 17276 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19248 6196 19300 6248
rect 19432 6196 19484 6248
rect 21088 6264 21140 6316
rect 20996 6196 21048 6248
rect 16028 6060 16080 6112
rect 22192 6128 22244 6180
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 20 5856 72 5908
rect 13360 5856 13412 5908
rect 14464 5856 14516 5908
rect 14740 5856 14792 5908
rect 15936 5856 15988 5908
rect 17960 5856 18012 5908
rect 19064 5856 19116 5908
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 20444 5856 20496 5908
rect 2688 5788 2740 5840
rect 4160 5788 4212 5840
rect 4528 5831 4580 5840
rect 4528 5797 4537 5831
rect 4537 5797 4571 5831
rect 4571 5797 4580 5831
rect 4528 5788 4580 5797
rect 5080 5831 5132 5840
rect 5080 5797 5089 5831
rect 5089 5797 5123 5831
rect 5123 5797 5132 5831
rect 5080 5788 5132 5797
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 2872 5720 2924 5772
rect 4252 5720 4304 5772
rect 7748 5720 7800 5772
rect 8760 5720 8812 5772
rect 8576 5652 8628 5704
rect 15844 5788 15896 5840
rect 19524 5788 19576 5840
rect 20076 5788 20128 5840
rect 12900 5720 12952 5772
rect 9588 5652 9640 5704
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12440 5695 12492 5704
rect 12256 5652 12308 5661
rect 12440 5661 12458 5695
rect 12458 5661 12492 5695
rect 12440 5652 12492 5661
rect 13360 5652 13412 5704
rect 14832 5695 14884 5704
rect 8300 5584 8352 5636
rect 9864 5584 9916 5636
rect 11152 5584 11204 5636
rect 10968 5516 11020 5568
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 15660 5720 15712 5772
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 19616 5720 19668 5772
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 20168 5720 20220 5772
rect 17960 5652 18012 5704
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 18880 5652 18932 5704
rect 20628 5652 20680 5704
rect 16488 5584 16540 5636
rect 15476 5516 15528 5568
rect 20996 5584 21048 5636
rect 19892 5559 19944 5568
rect 19892 5525 19901 5559
rect 19901 5525 19935 5559
rect 19935 5525 19944 5559
rect 19892 5516 19944 5525
rect 22284 5516 22336 5568
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 2320 5312 2372 5364
rect 4252 5312 4304 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 5448 5312 5500 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 12348 5312 12400 5364
rect 12440 5312 12492 5364
rect 5816 5244 5868 5296
rect 5724 5176 5776 5228
rect 6644 5176 6696 5228
rect 10968 5244 11020 5296
rect 15292 5244 15344 5296
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9864 5176 9916 5228
rect 10416 5176 10468 5228
rect 13176 5176 13228 5228
rect 12164 5108 12216 5160
rect 12440 5108 12492 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12900 5151 12952 5160
rect 12624 5108 12676 5117
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 14188 5151 14240 5160
rect 7932 5040 7984 5092
rect 8484 4972 8536 5024
rect 10784 4972 10836 5024
rect 12808 4972 12860 5024
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 19892 5312 19944 5364
rect 16672 5244 16724 5296
rect 17592 5244 17644 5296
rect 18420 5244 18472 5296
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 18696 5176 18748 5228
rect 20996 5176 21048 5228
rect 21640 5176 21692 5228
rect 22284 5312 22336 5364
rect 22468 5244 22520 5296
rect 19432 5108 19484 5160
rect 20628 5108 20680 5160
rect 19340 5040 19392 5092
rect 14188 4972 14240 5024
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 17224 4972 17276 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20628 4972 20680 5024
rect 22284 4972 22336 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 4804 4768 4856 4820
rect 4896 4768 4948 4820
rect 6644 4811 6696 4820
rect 6644 4777 6653 4811
rect 6653 4777 6687 4811
rect 6687 4777 6696 4811
rect 6644 4768 6696 4777
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 12624 4768 12676 4820
rect 10416 4700 10468 4752
rect 12992 4743 13044 4752
rect 12992 4709 13001 4743
rect 13001 4709 13035 4743
rect 13035 4709 13044 4743
rect 12992 4700 13044 4709
rect 10508 4632 10560 4684
rect 14648 4632 14700 4684
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 9496 4564 9548 4616
rect 8300 4496 8352 4548
rect 12992 4564 13044 4616
rect 14740 4564 14792 4616
rect 16212 4632 16264 4684
rect 19984 4632 20036 4684
rect 17040 4564 17092 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 22192 4564 22244 4616
rect 22928 4564 22980 4616
rect 9864 4496 9916 4548
rect 10232 4496 10284 4548
rect 11152 4496 11204 4548
rect 10416 4428 10468 4480
rect 11336 4428 11388 4480
rect 11888 4428 11940 4480
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 13360 4471 13412 4480
rect 12256 4428 12308 4437
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 20536 4496 20588 4548
rect 24492 4496 24544 4548
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 16580 4428 16632 4480
rect 20904 4471 20956 4480
rect 20904 4437 20913 4471
rect 20913 4437 20947 4471
rect 20947 4437 20956 4471
rect 20904 4428 20956 4437
rect 21456 4471 21508 4480
rect 21456 4437 21465 4471
rect 21465 4437 21499 4471
rect 21499 4437 21508 4471
rect 21456 4428 21508 4437
rect 22744 4428 22796 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 5724 4224 5776 4276
rect 17224 4267 17276 4276
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 10784 4156 10836 4208
rect 17224 4233 17233 4267
rect 17233 4233 17267 4267
rect 17267 4233 17276 4267
rect 17224 4224 17276 4233
rect 9864 4088 9916 4140
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 11980 4088 12032 4140
rect 14188 4088 14240 4140
rect 14556 4131 14608 4140
rect 14556 4097 14590 4131
rect 14590 4097 14608 4131
rect 14556 4088 14608 4097
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16396 4088 16448 4140
rect 19432 4156 19484 4208
rect 19984 4156 20036 4208
rect 20628 4224 20680 4276
rect 20720 4156 20772 4208
rect 21640 4156 21692 4208
rect 22284 4199 22336 4208
rect 22284 4165 22318 4199
rect 22318 4165 22336 4199
rect 22284 4156 22336 4165
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 10416 4020 10468 4072
rect 16764 4020 16816 4072
rect 20076 4088 20128 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 20904 4020 20956 4072
rect 12348 3952 12400 4004
rect 15292 3952 15344 4004
rect 21364 3995 21416 4004
rect 21364 3961 21373 3995
rect 21373 3961 21407 3995
rect 21407 3961 21416 3995
rect 21364 3952 21416 3961
rect 23204 3952 23256 4004
rect 23388 3995 23440 4004
rect 23388 3961 23397 3995
rect 23397 3961 23431 3995
rect 23431 3961 23440 3995
rect 23388 3952 23440 3961
rect 9312 3884 9364 3936
rect 11980 3927 12032 3936
rect 11980 3893 11989 3927
rect 11989 3893 12023 3927
rect 12023 3893 12032 3927
rect 11980 3884 12032 3893
rect 15568 3884 15620 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 16120 3927 16172 3936
rect 15660 3884 15712 3893
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 19616 3884 19668 3936
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 22928 3884 22980 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 9588 3680 9640 3732
rect 11704 3680 11756 3732
rect 12256 3680 12308 3732
rect 11520 3612 11572 3664
rect 13360 3680 13412 3732
rect 16304 3680 16356 3732
rect 20352 3680 20404 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 22192 3680 22244 3732
rect 23112 3723 23164 3732
rect 20168 3655 20220 3664
rect 20168 3621 20177 3655
rect 20177 3621 20211 3655
rect 20211 3621 20220 3655
rect 20168 3612 20220 3621
rect 8300 3544 8352 3596
rect 13820 3544 13872 3596
rect 14648 3544 14700 3596
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 11704 3476 11756 3528
rect 9680 3408 9732 3460
rect 9128 3340 9180 3392
rect 12164 3408 12216 3460
rect 11888 3340 11940 3392
rect 15292 3476 15344 3528
rect 15936 3519 15988 3528
rect 15936 3485 15945 3519
rect 15945 3485 15979 3519
rect 15979 3485 15988 3519
rect 15936 3476 15988 3485
rect 16580 3476 16632 3528
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 19708 3476 19760 3528
rect 22744 3476 22796 3528
rect 23388 3587 23440 3596
rect 23388 3553 23397 3587
rect 23397 3553 23431 3587
rect 23431 3553 23440 3587
rect 23388 3544 23440 3553
rect 23572 3544 23624 3596
rect 23480 3476 23532 3528
rect 21456 3408 21508 3460
rect 23204 3408 23256 3460
rect 12992 3340 13044 3392
rect 16304 3340 16356 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 19616 3340 19668 3392
rect 20996 3340 21048 3392
rect 22376 3340 22428 3392
rect 23296 3340 23348 3392
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 9128 3136 9180 3188
rect 11152 3179 11204 3188
rect 8392 3068 8444 3120
rect 9864 3068 9916 3120
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 11796 3136 11848 3188
rect 15568 3136 15620 3188
rect 16028 3136 16080 3188
rect 19524 3136 19576 3188
rect 19984 3136 20036 3188
rect 11060 3068 11112 3120
rect 11888 3068 11940 3120
rect 16488 3068 16540 3120
rect 9220 3000 9272 3052
rect 9404 3000 9456 3052
rect 12072 3000 12124 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 17316 3043 17368 3052
rect 10968 2932 11020 2984
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 18880 3043 18932 3052
rect 18880 3009 18898 3043
rect 18898 3009 18932 3043
rect 18880 3000 18932 3009
rect 19340 3000 19392 3052
rect 22468 3136 22520 3188
rect 23572 3136 23624 3188
rect 23848 3136 23900 3188
rect 23940 3136 23992 3188
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 24584 3068 24636 3120
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 22100 3000 22152 3052
rect 23204 3000 23256 3052
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 572 2796 624 2848
rect 6092 2796 6144 2848
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 8300 2796 8352 2848
rect 11520 2796 11572 2848
rect 12716 2796 12768 2848
rect 14648 2796 14700 2848
rect 29276 2932 29328 2984
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 18144 2796 18196 2848
rect 21364 2839 21416 2848
rect 21364 2805 21373 2839
rect 21373 2805 21407 2839
rect 21407 2805 21416 2839
rect 21364 2796 21416 2805
rect 22652 2796 22704 2848
rect 24492 2864 24544 2916
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 8484 2592 8536 2644
rect 9680 2592 9732 2644
rect 11704 2592 11756 2644
rect 10508 2524 10560 2576
rect 4988 2388 5040 2440
rect 9404 2456 9456 2508
rect 15936 2592 15988 2644
rect 16304 2635 16356 2644
rect 16304 2601 16313 2635
rect 16313 2601 16347 2635
rect 16347 2601 16356 2635
rect 16304 2592 16356 2601
rect 18880 2592 18932 2644
rect 21548 2592 21600 2644
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 12532 2456 12584 2508
rect 12992 2499 13044 2508
rect 12992 2465 13001 2499
rect 13001 2465 13035 2499
rect 13035 2465 13044 2499
rect 12992 2456 13044 2465
rect 13820 2456 13872 2508
rect 16028 2524 16080 2576
rect 9864 2388 9916 2440
rect 10784 2388 10836 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 15476 2388 15528 2440
rect 16304 2388 16356 2440
rect 19340 2524 19392 2576
rect 21456 2524 21508 2576
rect 22376 2567 22428 2576
rect 22376 2533 22385 2567
rect 22385 2533 22419 2567
rect 22419 2533 22428 2567
rect 22376 2524 22428 2533
rect 22928 2524 22980 2576
rect 20260 2456 20312 2508
rect 20444 2456 20496 2508
rect 23756 2524 23808 2576
rect 23112 2456 23164 2508
rect 19156 2388 19208 2440
rect 19248 2388 19300 2440
rect 19616 2388 19668 2440
rect 20720 2388 20772 2440
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 23388 2388 23440 2440
rect 23848 2388 23900 2440
rect 24860 2388 24912 2440
rect 25964 2388 26016 2440
rect 27068 2388 27120 2440
rect 28172 2431 28224 2440
rect 28172 2397 28181 2431
rect 28181 2397 28215 2431
rect 28215 2397 28224 2431
rect 28172 2388 28224 2397
rect 1676 2252 1728 2304
rect 2780 2252 2832 2304
rect 3884 2252 3936 2304
rect 9312 2320 9364 2372
rect 9588 2252 9640 2304
rect 11060 2320 11112 2372
rect 11612 2252 11664 2304
rect 13820 2320 13872 2372
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 15292 2320 15344 2372
rect 16120 2252 16172 2304
rect 16396 2252 16448 2304
rect 18236 2320 18288 2372
rect 18144 2252 18196 2304
rect 19248 2252 19300 2304
rect 23296 2320 23348 2372
rect 24768 2252 24820 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 8392 2048 8444 2100
rect 11244 2048 11296 2100
rect 8484 1980 8536 2032
rect 12900 1980 12952 2032
<< metal2 >>
rect 1306 29322 1362 30000
rect 32 29294 1362 29322
rect 32 5914 60 29294
rect 1306 29200 1362 29294
rect 3790 29200 3846 30000
rect 6274 29322 6330 30000
rect 8758 29322 8814 30000
rect 6274 29294 6592 29322
rect 6274 29200 6330 29294
rect 3804 27606 3832 29200
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 3792 27600 3844 27606
rect 3792 27542 3844 27548
rect 6564 27470 6592 29294
rect 8588 29294 8814 29322
rect 8588 27606 8616 29294
rect 8758 29200 8814 29294
rect 11242 29200 11298 30000
rect 13726 29200 13782 30000
rect 16210 29200 16266 30000
rect 18694 29200 18750 30000
rect 21178 29200 21234 30000
rect 23662 29200 23718 30000
rect 26146 29200 26202 30000
rect 28630 29322 28686 30000
rect 28368 29294 28686 29322
rect 8576 27600 8628 27606
rect 8576 27542 8628 27548
rect 11256 27470 11284 29200
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 13740 27554 13768 29200
rect 13740 27526 13860 27554
rect 13832 27470 13860 27526
rect 16224 27470 16252 29200
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 17868 27600 17920 27606
rect 17868 27542 17920 27548
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 6552 27464 6604 27470
rect 6552 27406 6604 27412
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 4172 26353 4200 27270
rect 6748 26858 6776 27270
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 6736 26852 6788 26858
rect 6736 26794 6788 26800
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 8404 26382 8432 26930
rect 8392 26376 8444 26382
rect 4158 26344 4214 26353
rect 4068 26308 4120 26314
rect 8392 26318 8444 26324
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 4158 26279 4214 26288
rect 4068 26250 4120 26256
rect 2136 26240 2188 26246
rect 2136 26182 2188 26188
rect 2596 26240 2648 26246
rect 2596 26182 2648 26188
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 2148 24954 2176 26182
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 2240 25158 2268 25842
rect 2608 25838 2636 26182
rect 2596 25832 2648 25838
rect 2596 25774 2648 25780
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2136 24948 2188 24954
rect 2136 24890 2188 24896
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 22506 1808 24006
rect 1860 23792 1912 23798
rect 1860 23734 1912 23740
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 18766 1624 20198
rect 1872 19689 1900 23734
rect 2148 23526 2176 24890
rect 2240 24070 2268 25094
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2136 23520 2188 23526
rect 2136 23462 2188 23468
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 2056 22710 2084 22918
rect 2044 22704 2096 22710
rect 2044 22646 2096 22652
rect 2148 21554 2176 23054
rect 2240 22982 2268 24006
rect 2228 22976 2280 22982
rect 2228 22918 2280 22924
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2240 22642 2268 22918
rect 2424 22778 2452 22918
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2136 21548 2188 21554
rect 2136 21490 2188 21496
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 2056 19922 2084 20742
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1858 19680 1914 19689
rect 1858 19615 1914 19624
rect 1872 19334 1900 19615
rect 2056 19378 2084 19858
rect 2240 19718 2268 22578
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2424 21962 2452 22374
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 1780 19306 1900 19334
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1688 15162 1716 18226
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1688 11762 1716 15098
rect 1780 14890 1808 19306
rect 2240 18290 2268 19654
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2148 17134 2176 17614
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 15706 2084 16526
rect 2148 16250 2176 17070
rect 2240 16574 2268 18022
rect 2332 17678 2360 21286
rect 2516 20262 2544 24550
rect 2608 23186 2636 25774
rect 2688 25764 2740 25770
rect 2688 25706 2740 25712
rect 2700 24614 2728 25706
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 23866 2728 24550
rect 3160 24206 3188 26182
rect 4080 26042 4108 26250
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 3712 25158 3740 25638
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2700 20534 2728 23802
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2792 21894 2820 22510
rect 2884 21962 2912 23462
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2872 21956 2924 21962
rect 2872 21898 2924 21904
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2688 20528 2740 20534
rect 2688 20470 2740 20476
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2516 18154 2544 20198
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2792 17270 2820 21286
rect 2976 21026 3004 22918
rect 3068 22642 3096 23122
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3160 22522 3188 24142
rect 3712 23118 3740 25094
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3068 22506 3188 22522
rect 3056 22500 3188 22506
rect 3108 22494 3188 22500
rect 3056 22442 3108 22448
rect 3068 21554 3096 22442
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2884 20998 3004 21026
rect 2884 19446 2912 20998
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2976 18630 3004 20810
rect 3068 20806 3096 21490
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2240 16546 2360 16574
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1780 14074 1808 14826
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1768 13932 1820 13938
rect 1872 13920 1900 14554
rect 2056 14482 2084 15642
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2332 14414 2360 16546
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 1820 13892 1900 13920
rect 1952 13932 2004 13938
rect 1768 13874 1820 13880
rect 1952 13874 2004 13880
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1688 10674 1716 11698
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 9926 1716 10610
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1688 8634 1716 8910
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 7546 1808 13874
rect 1964 13841 1992 13874
rect 1950 13832 2006 13841
rect 1860 13796 1912 13802
rect 1950 13767 2006 13776
rect 1860 13738 1912 13744
rect 1872 13326 1900 13738
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 10266 1900 13262
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1964 9722 1992 11698
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2056 11354 2084 11630
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1964 8906 1992 9658
rect 2056 9586 2084 11290
rect 2148 10810 2176 13194
rect 2240 11898 2268 13874
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8566 1992 8842
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 20 5908 72 5914
rect 20 5850 72 5856
rect 2332 5370 2360 8910
rect 2424 8838 2452 12378
rect 2700 10266 2728 16458
rect 2976 16182 3004 18566
rect 3068 18426 3096 20334
rect 3160 19854 3188 22374
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3252 19514 3280 22918
rect 3712 22642 3740 23054
rect 3516 22636 3568 22642
rect 3700 22636 3752 22642
rect 3568 22596 3648 22624
rect 3516 22578 3568 22584
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3332 20528 3384 20534
rect 3330 20496 3332 20505
rect 3384 20496 3386 20505
rect 3330 20431 3386 20440
rect 3240 19508 3292 19514
rect 3292 19468 3372 19496
rect 3240 19450 3292 19456
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 3252 14618 3280 18158
rect 3344 18154 3372 19468
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3436 17882 3464 21626
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3528 17066 3556 21558
rect 3620 19922 3648 22596
rect 3700 22578 3752 22584
rect 3712 21554 3740 22578
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3528 16658 3556 17002
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3344 14822 3372 15370
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2792 10742 2820 13466
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2502 9480 2558 9489
rect 2502 9415 2558 9424
rect 2516 9178 2544 9415
rect 2884 9178 2912 11698
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 6866 2544 8298
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2700 6730 2728 8842
rect 2976 8498 3004 8978
rect 3068 8566 3096 13670
rect 3344 10062 3372 14758
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 8090 3004 8434
rect 3344 8090 3372 9522
rect 3436 8566 3464 13806
rect 3712 13190 3740 21490
rect 3804 20262 3832 24890
rect 3988 24614 4016 25230
rect 4712 25152 4764 25158
rect 4710 25120 4712 25129
rect 5080 25152 5132 25158
rect 4764 25120 4766 25129
rect 5080 25094 5132 25100
rect 4710 25055 4766 25064
rect 5092 24954 5120 25094
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24070 4016 24550
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 5000 24342 5028 24686
rect 5736 24682 5764 25298
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5736 24410 5764 24618
rect 5724 24404 5776 24410
rect 5644 24364 5724 24392
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 23594 4016 24006
rect 3976 23588 4028 23594
rect 3976 23530 4028 23536
rect 3792 20256 3844 20262
rect 3988 20244 4016 23530
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4080 22642 4108 23462
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 20398 4108 21966
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4068 20256 4120 20262
rect 3988 20216 4068 20244
rect 3792 20198 3844 20204
rect 4068 20198 4120 20204
rect 3804 20058 3832 20198
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 4080 19292 4108 20198
rect 4172 19786 4200 20470
rect 4264 20262 4292 24074
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 4356 21350 4384 23666
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4816 22030 4844 24006
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 4172 19417 4200 19722
rect 4158 19408 4214 19417
rect 4158 19343 4214 19352
rect 4080 19264 4292 19292
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3804 13802 3832 16050
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 8838 3556 11834
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 8838 3648 10610
rect 3712 8974 3740 12106
rect 3804 11830 3832 13738
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3896 10713 3924 18226
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3988 13530 4016 17614
rect 4080 15094 4108 18566
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4172 12850 4200 18702
rect 4264 17660 4292 19264
rect 4356 18358 4384 21286
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4724 20777 4752 20810
rect 4804 20800 4856 20806
rect 4710 20768 4766 20777
rect 4804 20742 4856 20748
rect 4710 20703 4766 20712
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4434 19544 4490 19553
rect 4434 19479 4490 19488
rect 4448 19378 4476 19479
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4724 19258 4752 19994
rect 4816 19553 4844 20742
rect 4908 20466 4936 24278
rect 5000 24206 5028 24278
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5368 23730 5396 24142
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 4988 22976 5040 22982
rect 4988 22918 5040 22924
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4802 19544 4858 19553
rect 4802 19479 4858 19488
rect 4908 19378 4936 19722
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4724 19230 4844 19258
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4816 18850 4844 19230
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4724 18822 4844 18850
rect 4724 18630 4752 18822
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4344 17672 4396 17678
rect 4264 17632 4344 17660
rect 4264 16574 4292 17632
rect 4344 17614 4396 17620
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 16674 4384 17478
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 17082 4752 17138
rect 4816 17082 4844 18702
rect 4908 17202 4936 19110
rect 5000 18766 5028 22918
rect 5092 21622 5120 23122
rect 5276 23118 5304 23530
rect 5368 23186 5396 23666
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 5092 19310 5120 21558
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5184 19242 5212 21830
rect 5276 20942 5304 23054
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5092 18426 5120 19110
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4986 17640 5042 17649
rect 5092 17610 5120 18226
rect 4986 17575 5042 17584
rect 5080 17604 5132 17610
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4724 17054 4844 17082
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4356 16646 4476 16674
rect 4344 16584 4396 16590
rect 4264 16546 4344 16574
rect 4344 16526 4396 16532
rect 4448 16522 4476 16646
rect 4436 16516 4488 16522
rect 4436 16458 4488 16464
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4264 12986 4292 14350
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4356 12434 4384 16390
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4816 15570 4844 17054
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4620 15496 4672 15502
rect 4618 15464 4620 15473
rect 4672 15464 4674 15473
rect 4618 15399 4674 15408
rect 4712 15020 4764 15026
rect 4908 15008 4936 15846
rect 5000 15502 5028 17575
rect 5080 17546 5132 17552
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4764 14980 4936 15008
rect 4712 14962 4764 14968
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4816 13326 4844 14980
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4434 12744 4490 12753
rect 4540 12730 4568 13262
rect 4724 12986 4752 13262
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4710 12880 4766 12889
rect 4710 12815 4712 12824
rect 4764 12815 4766 12824
rect 4804 12844 4856 12850
rect 4712 12786 4764 12792
rect 4804 12786 4856 12792
rect 4816 12730 4844 12786
rect 4540 12702 4844 12730
rect 4434 12679 4490 12688
rect 4448 12646 4476 12679
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4264 12406 4384 12434
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3882 10704 3938 10713
rect 3882 10639 3938 10648
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3620 8498 3648 8774
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3422 7984 3478 7993
rect 3422 7919 3424 7928
rect 3476 7919 3478 7928
rect 3424 7890 3476 7896
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2700 6322 2728 6666
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6458 3372 6598
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3620 6322 3648 8434
rect 3896 6866 3924 10542
rect 3988 9110 4016 12106
rect 4080 9450 4108 12106
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4080 7818 4108 9386
rect 4172 8974 4200 9998
rect 4264 9994 4292 12406
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4356 11150 4384 11630
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4816 11234 4844 12702
rect 4448 11206 4844 11234
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10810 4384 11086
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4448 10452 4476 11206
rect 4908 11098 4936 14282
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4816 11070 4936 11098
rect 4724 10810 4752 11018
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4356 10424 4476 10452
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4172 7546 4200 8910
rect 4264 7886 4292 8978
rect 4356 8022 4384 10424
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4816 9738 4844 11070
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4724 9710 4844 9738
rect 4724 9654 4752 9710
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4816 9042 4844 9522
rect 4908 9178 4936 10746
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 2700 5846 2728 6258
rect 3620 6118 3648 6258
rect 4172 6186 4200 7482
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2884 5778 2912 6054
rect 4172 5846 4200 6122
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4264 5778 4292 7822
rect 4356 7478 4384 7958
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4356 6866 4384 7414
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4816 6934 4844 8230
rect 4908 7818 4936 8434
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 7410 4936 7754
rect 5000 7546 5028 15438
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5092 14346 5120 15030
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 12850 5120 14282
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5184 12753 5212 18566
rect 5276 16726 5304 20742
rect 5368 19446 5396 22986
rect 5460 21894 5488 24006
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 20806 5488 21830
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5446 20360 5502 20369
rect 5446 20295 5502 20304
rect 5460 19689 5488 20295
rect 5446 19680 5502 19689
rect 5446 19615 5502 19624
rect 5460 19446 5488 19615
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5368 18970 5396 19382
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5368 17678 5396 18226
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5276 15026 5304 15302
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5170 12744 5226 12753
rect 5170 12679 5226 12688
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12481 5120 12582
rect 5078 12472 5134 12481
rect 5276 12434 5304 14486
rect 5368 14414 5396 16934
rect 5552 16794 5580 20470
rect 5644 19786 5672 24364
rect 5724 24346 5776 24352
rect 5828 23730 5856 25638
rect 6472 25265 6500 26182
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6458 25256 6514 25265
rect 6458 25191 6514 25200
rect 6472 25158 6500 25191
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6472 24342 6500 25094
rect 6460 24336 6512 24342
rect 6460 24278 6512 24284
rect 6472 24206 6500 24278
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 6288 22778 6316 24074
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 5736 22438 5764 22714
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5736 20534 5764 22374
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5460 15162 5488 15370
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5078 12407 5134 12416
rect 5184 12406 5304 12434
rect 5078 10976 5134 10985
rect 5078 10911 5134 10920
rect 5092 10674 5120 10911
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9586 5120 9862
rect 5184 9654 5212 12406
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5276 11014 5304 12038
rect 5368 11830 5396 13126
rect 5460 12850 5488 14418
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10062 5304 10950
rect 5368 10690 5396 11766
rect 5460 10810 5488 12786
rect 5552 12238 5580 13942
rect 5644 12714 5672 17206
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5736 12850 5764 16730
rect 5828 15026 5856 20198
rect 5920 17814 5948 22374
rect 6380 20262 6408 23666
rect 6472 22642 6500 24142
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 22710 6684 24006
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6472 20466 6500 22578
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6564 22030 6592 22510
rect 6748 22030 6776 23462
rect 6932 22094 6960 25774
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7668 25265 7696 25638
rect 7654 25256 7710 25265
rect 7654 25191 7710 25200
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7024 24206 7052 24686
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7024 23186 7052 24142
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 6932 22066 7052 22094
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6564 21146 6592 21966
rect 7024 21486 7052 22066
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6380 19553 6408 20198
rect 6564 19854 6592 20198
rect 6552 19848 6604 19854
rect 6550 19816 6552 19825
rect 6604 19816 6606 19825
rect 6550 19751 6606 19760
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6366 19544 6422 19553
rect 6000 19508 6052 19514
rect 6366 19479 6422 19488
rect 6000 19450 6052 19456
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 6012 17066 6040 19450
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 6380 14414 6408 19479
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6748 18222 6776 19314
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 17882 6776 18158
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6642 17504 6698 17513
rect 6472 17270 6500 17478
rect 6642 17439 6698 17448
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6564 16454 6592 17138
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6552 15972 6604 15978
rect 6656 15960 6684 17439
rect 6840 17202 6868 19722
rect 7024 19446 7052 21286
rect 7116 21146 7144 21490
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 17610 7052 18566
rect 7116 18358 7144 20198
rect 7208 19854 7236 21014
rect 7300 20942 7328 23598
rect 7484 23322 7512 23666
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 8312 23118 8340 26182
rect 8404 25514 8432 26318
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8496 25906 8524 26250
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8404 25498 8524 25514
rect 8404 25492 8536 25498
rect 8404 25486 8484 25492
rect 8484 25434 8536 25440
rect 8588 24682 8616 26318
rect 8956 25906 8984 26998
rect 9404 26920 9456 26926
rect 9324 26868 9404 26874
rect 9324 26862 9456 26868
rect 9324 26846 9444 26862
rect 9324 26382 9352 26846
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9324 25974 9352 26318
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 8944 25900 8996 25906
rect 8944 25842 8996 25848
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 8956 25430 8984 25842
rect 8944 25424 8996 25430
rect 8944 25366 8996 25372
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8496 23798 8524 24006
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 7656 23112 7708 23118
rect 8300 23112 8352 23118
rect 7656 23054 7708 23060
rect 8298 23080 8300 23089
rect 8484 23112 8536 23118
rect 8352 23080 8354 23089
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 20936 7340 20942
rect 7392 20913 7420 21490
rect 7288 20878 7340 20884
rect 7378 20904 7434 20913
rect 7378 20839 7434 20848
rect 7484 20262 7512 22714
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7576 20466 7604 21490
rect 7668 20602 7696 23054
rect 8484 23054 8536 23060
rect 8298 23015 8354 23024
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 21570 7788 22918
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 8312 22438 8340 23015
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7760 21554 8064 21570
rect 7760 21548 8076 21554
rect 7760 21542 8024 21548
rect 8024 21490 8076 21496
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 16130 6776 16526
rect 6840 16250 6868 17138
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6748 16114 6868 16130
rect 6736 16108 6868 16114
rect 6788 16102 6868 16108
rect 6736 16050 6788 16056
rect 6604 15932 6684 15960
rect 6736 15972 6788 15978
rect 6552 15914 6604 15920
rect 6736 15914 6788 15920
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5828 13734 5856 14010
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5736 12646 5764 12786
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5368 10662 5488 10690
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8956 5120 9522
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5172 8968 5224 8974
rect 5092 8928 5172 8956
rect 5172 8910 5224 8916
rect 5276 8634 5304 9114
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8129 5120 8434
rect 5078 8120 5134 8129
rect 5078 8055 5134 8064
rect 5078 7984 5134 7993
rect 5078 7919 5134 7928
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6390 4384 6802
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4264 5370 4292 5714
rect 4540 5370 4568 5782
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4816 4826 4844 6870
rect 4908 4826 4936 7346
rect 4986 6896 5042 6905
rect 4986 6831 4988 6840
rect 5040 6831 5042 6840
rect 4988 6802 5040 6808
rect 5092 5846 5120 7919
rect 5368 7886 5396 10542
rect 5460 9110 5488 10662
rect 5552 10266 5580 12174
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10010 5672 11698
rect 5724 10804 5776 10810
rect 5828 10792 5856 13194
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 10810 5948 13126
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5998 12744 6054 12753
rect 5998 12679 6054 12688
rect 6012 12646 6040 12679
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5776 10764 5856 10792
rect 5908 10804 5960 10810
rect 5724 10746 5776 10752
rect 5908 10746 5960 10752
rect 5722 10704 5778 10713
rect 6012 10690 6040 11494
rect 5722 10639 5724 10648
rect 5776 10639 5778 10648
rect 5920 10662 6040 10690
rect 5724 10610 5776 10616
rect 5552 9982 5672 10010
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5552 8634 5580 9982
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5460 6458 5488 8502
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5552 8294 5580 8327
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5644 7410 5672 9318
rect 5736 8838 5764 9386
rect 5828 9382 5856 9551
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5722 8528 5778 8537
rect 5722 8463 5724 8472
rect 5776 8463 5778 8472
rect 5828 8480 5856 8910
rect 5920 8634 5948 10662
rect 6104 9654 6132 12786
rect 6196 11354 6224 13806
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6288 11558 6316 13194
rect 6380 11694 6408 14350
rect 6458 13968 6514 13977
rect 6458 13903 6460 13912
rect 6512 13903 6514 13912
rect 6460 13874 6512 13880
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6472 12918 6500 13738
rect 6564 13530 6592 15914
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6196 9674 6224 11290
rect 6380 10130 6408 11630
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6092 9648 6144 9654
rect 6012 9596 6092 9602
rect 6196 9646 6316 9674
rect 6380 9654 6408 10066
rect 6012 9590 6144 9596
rect 6012 9574 6132 9590
rect 6012 8634 6040 9574
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 8974 6132 9454
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5908 8492 5960 8498
rect 5828 8452 5908 8480
rect 5724 8434 5776 8440
rect 5908 8434 5960 8440
rect 5736 7954 5764 8434
rect 6104 8090 6132 8910
rect 6184 8900 6236 8906
rect 6288 8888 6316 9646
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6472 9586 6500 12854
rect 6656 12832 6684 15506
rect 6748 15162 6776 15914
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6840 12889 6868 16102
rect 6564 12804 6684 12832
rect 6826 12880 6882 12889
rect 6826 12815 6882 12824
rect 6564 11898 6592 12804
rect 6932 12764 6960 17138
rect 7024 15502 7052 17546
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15502 7144 15846
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14482 7144 14962
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7208 13326 7236 17478
rect 7300 17066 7328 19926
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7484 19378 7512 19654
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7286 14376 7342 14385
rect 7286 14311 7342 14320
rect 7300 14074 7328 14311
rect 7392 14278 7420 16118
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7300 13172 7328 13874
rect 7208 13144 7328 13172
rect 7102 12880 7158 12889
rect 7012 12844 7064 12850
rect 7102 12815 7158 12824
rect 7012 12786 7064 12792
rect 6656 12736 6960 12764
rect 6656 12442 6684 12736
rect 6828 12640 6880 12646
rect 7024 12617 7052 12786
rect 6828 12582 6880 12588
rect 7010 12608 7066 12617
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6840 12238 6868 12582
rect 7010 12543 7066 12552
rect 7116 12458 7144 12815
rect 7024 12430 7144 12458
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6564 11014 6592 11698
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6550 10704 6606 10713
rect 6550 10639 6606 10648
rect 6564 10130 6592 10639
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6236 8860 6316 8888
rect 6184 8842 6236 8848
rect 6564 8537 6592 10066
rect 6656 8974 6684 10406
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8634 6684 8774
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6550 8528 6606 8537
rect 6550 8463 6606 8472
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5184 5370 5212 6054
rect 5460 5370 5488 6394
rect 5736 5846 5764 7890
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5828 6118 5856 6802
rect 6656 6798 6684 8570
rect 6748 7546 6776 11018
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6840 9926 6868 10610
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9722 6868 9862
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6932 9160 6960 12038
rect 7024 11898 7052 12430
rect 7208 12102 7236 13144
rect 7392 12986 7420 14214
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7300 10810 7328 12786
rect 7484 12714 7512 16594
rect 7576 12850 7604 19654
rect 7668 19446 7696 20334
rect 7760 20058 7788 21422
rect 8298 20904 8354 20913
rect 8298 20839 8354 20848
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7852 20369 7880 20538
rect 8114 20496 8170 20505
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8024 20460 8076 20466
rect 8114 20431 8170 20440
rect 8024 20402 8076 20408
rect 7838 20360 7894 20369
rect 7838 20295 7894 20304
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 20058 7880 20198
rect 7944 20058 7972 20402
rect 8036 20369 8064 20402
rect 8022 20360 8078 20369
rect 8022 20295 8078 20304
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8128 19990 8156 20431
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7748 19916 7800 19922
rect 7800 19876 7880 19904
rect 7748 19858 7800 19864
rect 7852 19836 7880 19876
rect 8116 19848 8168 19854
rect 7852 19808 8116 19836
rect 8116 19790 8168 19796
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 7668 18426 7696 19382
rect 7760 18970 7788 19722
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 8312 19514 8340 20839
rect 8404 20806 8432 22034
rect 8496 21010 8524 23054
rect 8588 22710 8616 24346
rect 8576 22704 8628 22710
rect 8680 22681 8708 25230
rect 8956 24954 8984 25366
rect 9140 25276 9168 25842
rect 9220 25288 9272 25294
rect 9140 25248 9220 25276
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8944 24948 8996 24954
rect 8944 24890 8996 24896
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 24342 8800 24686
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8772 23866 8800 24278
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 8772 22692 8800 23802
rect 8864 23322 8892 24754
rect 9048 24274 9076 25162
rect 9140 24886 9168 25248
rect 9220 25230 9272 25236
rect 9220 25152 9272 25158
rect 9220 25094 9272 25100
rect 9128 24880 9180 24886
rect 9128 24822 9180 24828
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 9048 23866 9076 24074
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9048 22778 9076 23054
rect 9140 22982 9168 24822
rect 9232 24818 9260 25094
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9232 24206 9260 24754
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 8576 22646 8628 22652
rect 8666 22672 8722 22681
rect 8588 22030 8616 22646
rect 8772 22664 8984 22692
rect 8956 22658 8984 22664
rect 9140 22658 9168 22714
rect 8956 22630 9168 22658
rect 9232 22642 9260 24142
rect 9324 24138 9352 25910
rect 9784 25702 9812 26182
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9416 25265 9444 25298
rect 9680 25288 9732 25294
rect 9402 25256 9458 25265
rect 9680 25230 9732 25236
rect 9402 25191 9458 25200
rect 9588 25220 9640 25226
rect 9588 25162 9640 25168
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 9416 24954 9444 25094
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9416 24018 9444 24890
rect 9600 24818 9628 25162
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9692 24750 9720 25230
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9324 23990 9444 24018
rect 9324 23066 9352 23990
rect 9496 23724 9548 23730
rect 9416 23684 9496 23712
rect 9416 23186 9444 23684
rect 9496 23666 9548 23672
rect 9600 23594 9628 24142
rect 9692 23798 9720 24686
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9784 24206 9812 24550
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 9876 23662 9904 27066
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9968 26382 9996 26726
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9968 25906 9996 26318
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 10060 25498 10088 26726
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10152 25378 10180 27270
rect 10888 27130 10916 27270
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11796 26988 11848 26994
rect 11796 26930 11848 26936
rect 10704 26586 10732 26930
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10612 26042 10640 26318
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10060 25350 10180 25378
rect 10704 25362 10732 26522
rect 10980 26382 11008 26930
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 26586 11192 26726
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 11808 26382 11836 26930
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12268 26518 12296 26862
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12360 26382 12388 26794
rect 12636 26450 12664 27406
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10692 25356 10744 25362
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9324 23038 9444 23066
rect 9416 22982 9444 23038
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9324 22642 9352 22918
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9220 22636 9272 22642
rect 8666 22607 8722 22616
rect 8680 22094 8708 22607
rect 9220 22578 9272 22584
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9232 22098 9260 22578
rect 8680 22066 8984 22094
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8680 20942 8708 21014
rect 8668 20936 8720 20942
rect 8482 20904 8538 20913
rect 8668 20878 8720 20884
rect 8482 20839 8538 20848
rect 8576 20868 8628 20874
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 20262 8432 20742
rect 8496 20602 8524 20839
rect 8576 20810 8628 20816
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8404 19786 8432 20198
rect 8482 19816 8538 19825
rect 8392 19780 8444 19786
rect 8482 19751 8484 19760
rect 8392 19722 8444 19728
rect 8536 19751 8538 19760
rect 8484 19722 8536 19728
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18290 7788 18906
rect 8496 18766 8524 19110
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8496 18290 8524 18566
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7944 17678 7972 18090
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8404 17678 8432 17818
rect 8588 17814 8616 20810
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 7932 17672 7984 17678
rect 7930 17640 7932 17649
rect 8392 17672 8444 17678
rect 7984 17640 7986 17649
rect 7748 17604 7800 17610
rect 7930 17575 7986 17584
rect 8390 17640 8392 17649
rect 8444 17640 8446 17649
rect 8390 17575 8446 17584
rect 7748 17546 7800 17552
rect 7760 17513 7788 17546
rect 8300 17536 8352 17542
rect 7746 17504 7802 17513
rect 8300 17478 8352 17484
rect 7746 17439 7802 17448
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7668 15620 7696 17138
rect 7760 16522 7788 17138
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 16250 7788 16458
rect 8312 16454 8340 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 15632 7800 15638
rect 7668 15592 7748 15620
rect 7748 15574 7800 15580
rect 7760 13938 7788 15574
rect 7852 15473 7880 16050
rect 8024 15496 8076 15502
rect 7838 15464 7894 15473
rect 7838 15399 7894 15408
rect 8022 15464 8024 15473
rect 8076 15464 8078 15473
rect 8022 15399 8078 15408
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8312 13938 8340 14350
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 7654 13832 7710 13841
rect 7654 13767 7710 13776
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7668 12782 7696 13767
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7378 12608 7434 12617
rect 7378 12543 7434 12552
rect 7392 10810 7420 12543
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11558 7604 12106
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 8312 11880 8340 13262
rect 8220 11852 8340 11880
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7116 9994 7144 10610
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7012 9172 7064 9178
rect 6932 9132 7012 9160
rect 7012 9114 7064 9120
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8498 7144 8978
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 7546 7144 8434
rect 7208 8022 7236 9318
rect 7300 9178 7328 10746
rect 7392 10470 7420 10746
rect 7484 10742 7512 10950
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7576 9994 7604 11494
rect 8220 11014 8248 11852
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 8312 10198 8340 11698
rect 8404 11150 8432 17274
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8496 15706 8524 16458
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 14414 8524 14962
rect 8588 14958 8616 16526
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8680 14278 8708 19994
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8772 16794 8800 19314
rect 8864 17678 8892 21830
rect 8956 21162 8984 22066
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 9324 22030 9352 22578
rect 9416 22574 9444 22714
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9324 21690 9352 21966
rect 9416 21962 9444 22510
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 8956 21134 9076 21162
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20398 8984 20742
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8956 18222 8984 20334
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8864 16674 8892 17614
rect 8772 16646 8892 16674
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 12646 8524 13806
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8588 12238 8616 13670
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12481 8708 12786
rect 8666 12472 8722 12481
rect 8666 12407 8722 12416
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8036 10062 8064 10134
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7392 9674 7420 9930
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 7392 9646 7696 9674
rect 7668 9518 7696 9646
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7116 7002 7144 7346
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6254 6684 6734
rect 7208 6662 7236 7822
rect 7300 7410 7328 8230
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7478 7420 8026
rect 7484 7886 7512 8842
rect 7576 8430 7604 8910
rect 7668 8838 7696 9114
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7392 6730 7420 7414
rect 7484 7002 7512 7482
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7484 6322 7512 6938
rect 7576 6798 7604 7686
rect 7668 6984 7696 8434
rect 7760 7954 7788 8774
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 8300 8424 8352 8430
rect 8220 8384 8300 8412
rect 8220 8129 8248 8384
rect 8300 8366 8352 8372
rect 8206 8120 8262 8129
rect 8206 8055 8262 8064
rect 8220 7954 8248 8055
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7760 7410 7788 7890
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7748 6996 7800 7002
rect 7668 6956 7748 6984
rect 7748 6938 7800 6944
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7760 6458 7788 6938
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8312 6458 8340 6870
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6390 8432 10950
rect 8496 7546 8524 12106
rect 8588 11218 8616 12174
rect 8680 11898 8708 12310
rect 8772 12220 8800 16646
rect 8956 16574 8984 18158
rect 9048 18154 9076 21134
rect 9310 20360 9366 20369
rect 9310 20295 9366 20304
rect 9324 20262 9352 20295
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9508 19922 9536 23462
rect 9600 22778 9628 23530
rect 9876 23118 9904 23598
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 10060 23050 10088 25350
rect 10692 25298 10744 25304
rect 10796 25294 10824 25842
rect 10888 25430 10916 25978
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 10416 25288 10468 25294
rect 10784 25288 10836 25294
rect 10468 25248 10548 25276
rect 10416 25230 10468 25236
rect 10520 25242 10548 25248
rect 10520 25236 10784 25242
rect 10836 25236 10916 25242
rect 10520 25214 10916 25236
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10612 24274 10640 24754
rect 10888 24750 10916 25214
rect 11072 25158 11100 25978
rect 11152 25764 11204 25770
rect 11152 25706 11204 25712
rect 11164 25226 11192 25706
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11808 25498 11836 26318
rect 12728 25838 12756 26998
rect 12820 26994 12848 27406
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12912 26586 12940 26998
rect 13004 26994 13032 27270
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14004 27056 14056 27062
rect 14004 26998 14056 27004
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13820 26988 13872 26994
rect 13872 26948 13952 26976
rect 13820 26930 13872 26936
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 13096 26518 13124 26726
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 13188 26382 13216 26862
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11072 24886 11100 25094
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 10692 24608 10744 24614
rect 10980 24596 11008 24754
rect 10692 24550 10744 24556
rect 10888 24568 11008 24596
rect 10600 24268 10652 24274
rect 10600 24210 10652 24216
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 10152 22642 10180 23802
rect 10612 23730 10640 24006
rect 10704 23866 10732 24550
rect 10888 24342 10916 24568
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 11072 24188 11100 24822
rect 11808 24818 11836 25162
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11152 24200 11204 24206
rect 11072 24160 11152 24188
rect 11152 24142 11204 24148
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10980 23730 11008 24006
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10244 22642 10272 23598
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9600 19514 9628 20470
rect 9692 19922 9720 21830
rect 10336 21622 10364 22918
rect 10428 21962 10456 23054
rect 10612 22710 10640 23666
rect 10876 23044 10928 23050
rect 10876 22986 10928 22992
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10796 22642 10824 22918
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10888 22545 10916 22986
rect 11164 22982 11192 24142
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 11256 23118 11284 23462
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11716 23304 11744 23666
rect 11624 23276 11744 23304
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10874 22536 10930 22545
rect 10874 22471 10930 22480
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9126 19408 9182 19417
rect 9126 19343 9182 19352
rect 9220 19372 9272 19378
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9140 17882 9168 19343
rect 9220 19314 9272 19320
rect 9232 18426 9260 19314
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9508 18222 9536 18702
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9140 17066 9168 17818
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9232 16946 9260 18158
rect 9404 18080 9456 18086
rect 9600 18034 9628 19450
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9404 18022 9456 18028
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9324 17202 9352 17614
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9416 16998 9444 18022
rect 9508 18006 9628 18034
rect 8864 16546 8984 16574
rect 9048 16918 9260 16946
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 8864 12345 8892 16546
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 15434 8984 16390
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 8956 15042 8984 15370
rect 9048 15162 9076 16918
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9218 15464 9274 15473
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8956 15014 9076 15042
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8956 13870 8984 14350
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9048 13802 9076 15014
rect 9140 14890 9168 15438
rect 9218 15399 9274 15408
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13977 9168 14214
rect 9126 13968 9182 13977
rect 9126 13903 9182 13912
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 13394 9076 13738
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8942 12472 8998 12481
rect 8942 12407 8998 12416
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8956 12238 8984 12407
rect 8944 12232 8996 12238
rect 8772 12192 8892 12220
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8680 11082 8708 11494
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8864 10674 8892 12192
rect 8944 12174 8996 12180
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8956 10062 8984 12174
rect 9048 12102 9076 12582
rect 9140 12442 9168 13262
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9232 12238 9260 15399
rect 9324 12986 9352 16594
rect 9508 16182 9536 18006
rect 9692 17066 9720 19178
rect 10060 19174 10088 21286
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10244 20534 10272 20946
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9784 18086 9812 19110
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9876 17814 9904 18634
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9508 15638 9536 16118
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9416 13394 9444 14418
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9232 11898 9260 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11762 9352 12922
rect 9508 12434 9536 15370
rect 9680 15360 9732 15366
rect 9784 15348 9812 17614
rect 9876 17105 9904 17614
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9862 17096 9918 17105
rect 9862 17031 9918 17040
rect 9968 16046 9996 17138
rect 10046 17096 10102 17105
rect 10046 17031 10102 17040
rect 10060 16674 10088 17031
rect 10152 16776 10180 19654
rect 10428 19446 10456 21898
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10520 20466 10548 20742
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10888 19854 10916 22471
rect 10980 22098 11008 22646
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10980 20806 11008 21422
rect 11072 20942 11100 21830
rect 11164 21690 11192 22918
rect 11348 22642 11376 23122
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11624 22574 11652 23276
rect 11808 22642 11836 24754
rect 12084 24206 12112 25638
rect 12728 25294 12756 25774
rect 12820 25362 12848 25842
rect 12912 25498 12940 26318
rect 13188 26042 13216 26318
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 13280 25906 13308 26522
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12728 24954 12756 25230
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12820 24614 12848 25298
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24342 12848 24550
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12084 23712 12112 24142
rect 12268 23730 12296 24142
rect 12820 23730 12848 24278
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12256 23724 12308 23730
rect 12084 23684 12204 23712
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23118 12112 23462
rect 12176 23186 12204 23684
rect 12256 23666 12308 23672
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12912 23186 12940 24006
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11256 22234 11284 22442
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 11716 22166 11744 22578
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 11808 22098 11836 22578
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11808 21690 11836 22034
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 11900 20466 11928 22986
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11992 22545 12020 22578
rect 11978 22536 12034 22545
rect 11978 22471 12034 22480
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12084 20466 12112 22170
rect 12176 21622 12204 22374
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12728 22137 12756 22170
rect 12714 22128 12770 22137
rect 12440 22092 12492 22098
rect 12714 22063 12770 22072
rect 12808 22092 12860 22098
rect 12440 22034 12492 22040
rect 12808 22034 12860 22040
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 10980 19990 11008 20402
rect 11980 20392 12032 20398
rect 11978 20360 11980 20369
rect 12032 20360 12034 20369
rect 12452 20330 12480 22034
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 11978 20295 12034 20304
rect 12440 20324 12492 20330
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10244 18358 10272 18566
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10244 17678 10272 18294
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10336 17610 10364 18566
rect 10520 18222 10548 19110
rect 11072 18290 11100 19994
rect 11992 19922 12020 20295
rect 12440 20266 12492 20272
rect 12544 19922 12572 21898
rect 12636 20602 12664 21966
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 20058 12756 20402
rect 12820 20330 12848 22034
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21350 13032 21830
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13004 20380 13032 21082
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 12912 20352 13032 20380
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11256 18290 11284 19722
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17202 10272 17478
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 17105 10272 17138
rect 10230 17096 10286 17105
rect 10230 17031 10286 17040
rect 10232 16788 10284 16794
rect 10152 16748 10232 16776
rect 10232 16730 10284 16736
rect 10060 16646 10272 16674
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9732 15320 9812 15348
rect 9680 15302 9732 15308
rect 9784 15162 9812 15320
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9416 12406 9536 12434
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 10674 9076 11630
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9416 9654 9444 12406
rect 9494 12336 9550 12345
rect 9494 12271 9550 12280
rect 9508 12238 9536 12271
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11830 9536 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9600 10266 9628 14282
rect 10060 14074 10088 16458
rect 10152 16114 10180 16526
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 14890 10180 15914
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10152 13841 10180 14826
rect 10244 13938 10272 16646
rect 10336 16114 10364 17546
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 10796 17066 10824 17206
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10428 16182 10456 17002
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 10266 9720 12174
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10962 9904 11018
rect 9784 10934 9904 10962
rect 9784 10810 9812 10934
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9692 10146 9720 10202
rect 9600 10118 9720 10146
rect 9600 9926 9628 10118
rect 9784 9994 9812 10746
rect 10060 10606 10088 11698
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 8574 9072 8630 9081
rect 8574 9007 8576 9016
rect 8628 9007 8630 9016
rect 8576 8978 8628 8984
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 6798 8524 7142
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5736 5234 5764 5782
rect 5828 5302 5856 6054
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5736 4282 5764 5170
rect 6656 4826 6684 5170
rect 7300 4826 7328 6122
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 7760 4146 7788 5714
rect 8404 5658 8432 6326
rect 8588 5710 8616 6598
rect 8680 6322 8708 6666
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8772 5778 8800 8910
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 7886 9168 8774
rect 9416 8498 9444 9318
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8362 9444 8434
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7410 9168 7822
rect 9324 7818 9352 8298
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8312 5642 8432 5658
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8300 5636 8432 5642
rect 8352 5630 8432 5636
rect 8300 5578 8352 5584
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8208 5364 8260 5370
rect 8312 5352 8340 5578
rect 8260 5324 8340 5352
rect 8208 5306 8260 5312
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7944 4826 7972 5034
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 8312 3602 8340 4490
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8404 3534 8432 4558
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 8404 3126 8432 3470
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 584 800 612 2790
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 1688 800 1716 2246
rect 2792 800 2820 2246
rect 3896 800 3924 2246
rect 5000 800 5028 2382
rect 6104 800 6132 2790
rect 7208 800 7236 2790
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 8312 800 8340 2790
rect 8496 2650 8524 4966
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3194 9168 3334
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9232 3058 9260 7686
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9324 5234 9352 6258
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4078 9352 5170
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3074 9352 3878
rect 9416 3534 9444 7482
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9600 7154 9628 7278
rect 9692 7274 9720 8502
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9600 7126 9720 7154
rect 9692 7002 9720 7126
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6322 9628 6734
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9588 5704 9640 5710
rect 9508 5664 9588 5692
rect 9508 4622 9536 5664
rect 9692 5692 9720 6938
rect 9784 6798 9812 9930
rect 9864 8288 9916 8294
rect 9916 8236 9996 8242
rect 9864 8230 9996 8236
rect 9876 8214 9996 8230
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7410 9904 7822
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9968 7290 9996 8214
rect 10152 8090 10180 13767
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10244 12850 10272 13194
rect 10336 12866 10364 14214
rect 10428 13326 10456 14214
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10336 12850 10456 12866
rect 10232 12844 10284 12850
rect 10336 12844 10468 12850
rect 10336 12838 10416 12844
rect 10232 12786 10284 12792
rect 10416 12786 10468 12792
rect 10244 12434 10272 12786
rect 10244 12406 10364 12434
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7410 10088 7958
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9876 7262 9996 7290
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9640 5664 9720 5692
rect 9588 5646 9640 5652
rect 9876 5642 9904 7262
rect 10060 6730 10088 7346
rect 10244 6769 10272 9454
rect 10336 9178 10364 12406
rect 10428 12306 10456 12786
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 10198 10456 12106
rect 10520 11558 10548 16050
rect 10612 15978 10640 16934
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10704 15570 10732 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10674 10548 10950
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10506 10568 10562 10577
rect 10506 10503 10562 10512
rect 10520 10470 10548 10503
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10612 10130 10640 14758
rect 10704 14074 10732 15506
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10690 13968 10746 13977
rect 10690 13903 10692 13912
rect 10744 13903 10746 13912
rect 10692 13874 10744 13880
rect 10704 12850 10732 13874
rect 10796 13870 10824 16050
rect 10888 14634 10916 18158
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10980 15094 11008 17818
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 16182 11192 17478
rect 11716 17338 11744 19314
rect 11808 17354 11836 19790
rect 11992 19334 12020 19858
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 11992 19306 12112 19334
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 17678 11928 19110
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11992 18426 12020 18634
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11704 17332 11756 17338
rect 11808 17326 11928 17354
rect 11704 17274 11756 17280
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15434 11100 16050
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10888 14606 11008 14634
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10888 13938 10916 14486
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11121 10732 12174
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11286 10824 11494
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10690 11112 10746 11121
rect 10690 11047 10746 11056
rect 10784 11076 10836 11082
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10324 9172 10376 9178
rect 10376 9132 10548 9160
rect 10324 9114 10376 9120
rect 10230 6760 10286 6769
rect 10048 6724 10100 6730
rect 10230 6695 10286 6704
rect 10048 6666 10100 6672
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9876 5234 9904 5578
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 10244 4554 10272 6695
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10428 4758 10456 5170
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10520 4690 10548 9132
rect 10704 9042 10732 11047
rect 10784 11018 10836 11024
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 7954 10640 8774
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10704 6798 10732 8298
rect 10796 8090 10824 11018
rect 10888 8974 10916 13874
rect 10980 13326 11008 14606
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11072 12866 11100 15370
rect 11164 15026 11192 16118
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11256 14618 11284 15846
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11164 12986 11192 13874
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11072 12850 11192 12866
rect 11072 12844 11204 12850
rect 11072 12838 11152 12844
rect 11152 12786 11204 12792
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10968 10736 11020 10742
rect 10966 10704 10968 10713
rect 11020 10704 11022 10713
rect 10966 10639 11022 10648
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10980 8922 11008 9522
rect 11072 9382 11100 11086
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 9042 11100 9318
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10980 8894 11100 8922
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 11072 7886 11100 8894
rect 11164 8430 11192 12786
rect 11256 12442 11284 13942
rect 11716 13870 11744 14894
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11716 13530 11744 13806
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 13410 11836 16050
rect 11716 13382 11836 13410
rect 11716 12918 11744 13382
rect 11900 13190 11928 17326
rect 11992 15162 12020 18226
rect 12084 17082 12112 19306
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17270 12204 17546
rect 12360 17542 12388 18226
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12256 17196 12308 17202
rect 12308 17156 12388 17184
rect 12256 17138 12308 17144
rect 12084 17054 12296 17082
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 15162 12204 16934
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 13734 12020 14554
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11256 10742 11284 12378
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11348 10742 11376 11290
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11716 9738 11744 12854
rect 11886 12744 11942 12753
rect 11886 12679 11942 12688
rect 11900 12442 11928 12679
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11992 11898 12020 13670
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12084 11558 12112 12378
rect 12176 11830 12204 13194
rect 12268 12986 12296 17054
rect 12360 16794 12388 17156
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 16250 12480 19110
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12544 15366 12572 19246
rect 12636 16590 12664 19790
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12728 19417 12756 19450
rect 12714 19408 12770 19417
rect 12714 19343 12770 19352
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 16658 12756 18702
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 15706 12664 16526
rect 12728 16250 12756 16594
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12912 16130 12940 20352
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12728 16102 12940 16130
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12360 14414 12388 15030
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12438 14920 12494 14929
rect 12438 14855 12494 14864
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12452 14074 12480 14855
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13530 12572 14962
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12636 13190 12664 15098
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11624 9710 11744 9738
rect 11624 9518 11652 9710
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10980 7410 11008 7482
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 11072 6322 11100 7822
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11164 5642 11192 8366
rect 11256 8090 11284 8842
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11440 6390 11468 6666
rect 11716 6390 11744 9590
rect 11808 7478 11836 11494
rect 11978 10704 12034 10713
rect 11888 10668 11940 10674
rect 12176 10674 12204 11766
rect 12636 11762 12664 12718
rect 12728 12442 12756 16102
rect 12808 15496 12860 15502
rect 13004 15484 13032 18634
rect 13096 17882 13124 20810
rect 13188 20602 13216 25706
rect 13280 25362 13308 25842
rect 13360 25696 13412 25702
rect 13360 25638 13412 25644
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13280 24818 13308 25298
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 22642 13308 23122
rect 13372 23118 13400 25638
rect 13464 24818 13492 25978
rect 13648 25294 13676 26726
rect 13924 26450 13952 26948
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 13924 25838 13952 26386
rect 14016 25906 14044 26998
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13636 25288 13688 25294
rect 13636 25230 13688 25236
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13372 22574 13400 23054
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13464 22094 13492 22918
rect 13556 22778 13584 25230
rect 14108 24818 14136 25842
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13648 22642 13676 24006
rect 13740 22982 13768 24142
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13372 22066 13492 22094
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13372 20534 13400 22066
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13464 21146 13492 21966
rect 13648 21622 13676 22578
rect 13740 22030 13768 22918
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13176 20392 13228 20398
rect 13174 20360 13176 20369
rect 13228 20360 13230 20369
rect 13174 20295 13230 20304
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13188 19514 13216 20198
rect 13372 20058 13400 20198
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13464 19378 13492 20742
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13556 19258 13584 21422
rect 13832 21078 13860 24006
rect 13924 22710 13952 24210
rect 14016 23526 14044 24550
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13912 22704 13964 22710
rect 14016 22681 14044 23462
rect 13912 22646 13964 22652
rect 14002 22672 14058 22681
rect 13924 22438 13952 22646
rect 14002 22607 14004 22616
rect 14056 22607 14058 22616
rect 14004 22578 14056 22584
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13832 20330 13860 20810
rect 14016 20346 14044 22102
rect 14096 21956 14148 21962
rect 14096 21898 14148 21904
rect 14108 21690 14136 21898
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14200 20942 14228 21490
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14200 20398 14228 20878
rect 14292 20466 14320 26726
rect 15212 26450 15240 27270
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 15304 26382 15332 27270
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 17052 26586 17080 26726
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 17696 26382 17724 27270
rect 17788 26450 17816 27474
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 14372 26240 14424 26246
rect 14372 26182 14424 26188
rect 14384 25974 14412 26182
rect 14476 26042 14504 26318
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 15672 25294 15700 26182
rect 16224 25906 16252 26182
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16856 25764 16908 25770
rect 16856 25706 16908 25712
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14476 22094 14504 25094
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24206 15240 24550
rect 15764 24290 15792 25638
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 15672 24262 15792 24290
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14568 22234 14596 22986
rect 14660 22982 14688 24074
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 15212 23798 15240 24142
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14660 22098 14688 22918
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14476 22066 14596 22094
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14476 20777 14504 21830
rect 14568 20942 14596 22066
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14936 22030 14964 22510
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14188 20392 14240 20398
rect 13820 20324 13872 20330
rect 14016 20318 14136 20346
rect 14188 20334 14240 20340
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 13820 20266 13872 20272
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13648 19910 13860 19938
rect 14016 19922 14044 20198
rect 13648 19854 13676 19910
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 19417 13676 19654
rect 13634 19408 13690 19417
rect 13634 19343 13690 19352
rect 13452 19236 13504 19242
rect 13556 19230 13676 19258
rect 13452 19178 13504 19184
rect 13464 18970 13492 19178
rect 13544 19168 13596 19174
rect 13542 19136 13544 19145
rect 13596 19136 13598 19145
rect 13542 19071 13598 19080
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13372 18426 13400 18906
rect 13648 18766 13676 19230
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13464 18358 13492 18566
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12860 15456 13032 15484
rect 12808 15438 12860 15444
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 15026 13032 15302
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12912 14346 12940 14486
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 14006 12848 14214
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 12646 12848 13738
rect 13004 13172 13032 14962
rect 13096 14414 13124 17614
rect 13188 17270 13216 17750
rect 13464 17610 13492 18294
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13084 13184 13136 13190
rect 13004 13144 13084 13172
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 12238 12848 12582
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 10810 12756 11630
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 11978 10639 12034 10648
rect 12072 10668 12124 10674
rect 11888 10610 11940 10616
rect 11900 10577 11928 10610
rect 11886 10568 11942 10577
rect 11992 10538 12020 10639
rect 12072 10610 12124 10616
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11886 10503 11942 10512
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 12084 10266 12112 10610
rect 12176 10266 12204 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 8906 12020 9318
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11888 6996 11940 7002
rect 11992 6984 12020 7890
rect 11940 6956 12020 6984
rect 11888 6938 11940 6944
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10980 5302 11008 5510
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 9876 4146 9904 4490
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10428 4078 10456 4422
rect 10796 4214 10824 4966
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9324 3058 9444 3074
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9324 3052 9456 3058
rect 9324 3046 9404 3052
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8404 2106 8432 2382
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8496 2038 8524 2586
rect 9324 2378 9352 3046
rect 9404 2994 9456 3000
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 9416 800 9444 2450
rect 9600 2310 9628 3674
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9692 2650 9720 3402
rect 9876 3126 9904 3470
rect 11164 3194 11192 4490
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11348 4026 11376 4422
rect 11900 4298 11928 4422
rect 11256 3998 11376 4026
rect 11716 4270 11928 4298
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9876 2446 9904 3062
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10980 2774 11008 2926
rect 10796 2746 11008 2774
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 10520 800 10548 2518
rect 10796 2446 10824 2746
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11072 2378 11100 3062
rect 11164 2446 11192 3130
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11256 2106 11284 3998
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11716 3738 11744 4270
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 2854 11560 3606
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 11716 2650 11744 3470
rect 11808 3194 11836 4082
rect 11992 3942 12020 4082
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11900 3126 11928 3334
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 12084 3058 12112 10202
rect 12176 9586 12204 10202
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 7970 12296 8026
rect 12268 7942 12388 7970
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7342 12204 7822
rect 12360 7426 12388 7942
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12636 7546 12664 7890
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12438 7440 12494 7449
rect 12360 7398 12438 7426
rect 12438 7375 12494 7384
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12176 5692 12204 7278
rect 12452 6458 12480 7278
rect 12636 7002 12664 7278
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12728 6322 12756 7686
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12256 5704 12308 5710
rect 12176 5664 12256 5692
rect 12176 5250 12204 5664
rect 12440 5704 12492 5710
rect 12256 5646 12308 5652
rect 12360 5652 12440 5658
rect 12360 5646 12492 5652
rect 12360 5630 12480 5646
rect 12360 5370 12388 5630
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 5250 12480 5306
rect 12176 5222 12480 5250
rect 12176 5166 12204 5222
rect 12164 5160 12216 5166
rect 12440 5160 12492 5166
rect 12164 5102 12216 5108
rect 12360 5108 12440 5114
rect 12360 5102 12492 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12360 5086 12480 5102
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 3738 12296 4422
rect 12360 4010 12388 5086
rect 12636 4826 12664 5102
rect 12820 5030 12848 9862
rect 13004 9178 13032 13144
rect 13084 13126 13136 13132
rect 13188 12918 13216 17206
rect 13280 14414 13308 17478
rect 13556 17202 13584 17614
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13450 17096 13506 17105
rect 13450 17031 13506 17040
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13372 16182 13400 16458
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13464 16028 13492 17031
rect 13648 16726 13676 18702
rect 13740 17882 13768 19790
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13832 17610 13860 19910
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14016 19378 14044 19654
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14004 19168 14056 19174
rect 13924 19128 14004 19156
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13924 17338 13952 19128
rect 14004 19110 14056 19116
rect 14108 18222 14136 20318
rect 14200 19990 14228 20334
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 16794 14044 17478
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13372 16000 13492 16028
rect 13372 15434 13400 16000
rect 13556 15910 13584 16458
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 13977 13308 14350
rect 13372 14074 13400 15370
rect 13464 14958 13492 15438
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13556 14482 13584 14962
rect 13740 14822 13768 15302
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13266 13968 13322 13977
rect 13740 13938 13768 14282
rect 13266 13903 13322 13912
rect 13728 13932 13780 13938
rect 13280 13326 13308 13903
rect 13728 13874 13780 13880
rect 13832 13530 13860 14894
rect 13924 14822 13952 16118
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 13802 13952 14758
rect 14016 14006 14044 15982
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15094 14136 15846
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13924 12434 13952 13194
rect 14016 12850 14044 13942
rect 14108 13870 14136 15030
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14200 13734 14228 19926
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18698 14320 19110
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14384 14890 14412 20334
rect 14660 19922 14688 20946
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14292 14414 14320 14826
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14292 13258 14320 14350
rect 14476 13530 14504 19314
rect 14568 18902 14596 19790
rect 14660 18970 14688 19858
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14752 18358 14780 21966
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14936 19922 14964 20334
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 14830 19816 14886 19825
rect 14830 19751 14886 19760
rect 14844 19718 14872 19751
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 15212 18290 15240 23598
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22030 15332 22374
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15580 21690 15608 22578
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15396 19446 15424 20402
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15488 20058 15516 20266
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15488 19514 15516 19994
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14568 17678 14596 18090
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 14822 14596 16526
rect 14752 16522 14780 17478
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 15212 17202 15240 17818
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15212 16658 15240 17002
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 15304 16454 15332 17546
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 15706 14872 15982
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 15028 15502 15056 16050
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14660 14074 14688 14826
rect 14936 14822 14964 14962
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13734 14688 13874
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14752 13462 14780 14350
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 13841 15332 13874
rect 15290 13832 15346 13841
rect 15290 13767 15346 13776
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13924 12406 14044 12434
rect 14016 11286 14044 12406
rect 14108 12238 14136 12786
rect 14476 12442 14504 13262
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 15396 12986 15424 19382
rect 15580 18970 15608 21490
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15580 15366 15608 15982
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 15026 15608 15302
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 13734 15516 14758
rect 15580 14414 15608 14962
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13190 15516 13670
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14568 12238 14596 12650
rect 15304 12238 15332 12786
rect 15488 12782 15516 13126
rect 15580 12918 15608 14350
rect 15672 14074 15700 24262
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 15764 23866 15792 24074
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15948 23730 15976 25094
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15856 23322 15884 23666
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15948 22545 15976 23666
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 15934 22536 15990 22545
rect 15934 22471 15990 22480
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15764 21078 15792 21490
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15752 20460 15804 20466
rect 15856 20448 15884 21490
rect 15804 20420 15884 20448
rect 15752 20402 15804 20408
rect 15948 20380 15976 22471
rect 16040 21554 16068 23530
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16408 22778 16436 23462
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16132 22234 16160 22646
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16132 20466 16160 22170
rect 16316 21690 16344 22374
rect 16408 22166 16436 22714
rect 16396 22160 16448 22166
rect 16396 22102 16448 22108
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 21078 16344 21626
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 15856 20352 15976 20380
rect 15856 19334 15884 20352
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19854 16068 20198
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15948 19378 15976 19790
rect 15764 19306 15884 19334
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15764 18222 15792 19306
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15856 18290 15884 18770
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15856 17202 15884 18226
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15856 16114 15884 17138
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15856 15910 15884 16050
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15948 15706 15976 19314
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 17134 16068 18158
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16132 16114 16160 20402
rect 16224 20058 16252 21014
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16224 17202 16252 19994
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16224 16794 16252 17138
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16408 16182 16436 16662
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16132 15162 16160 16050
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14550 15792 14758
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 14096 12232 14148 12238
rect 14556 12232 14608 12238
rect 14096 12174 14148 12180
rect 14384 12192 14556 12220
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11830 14228 12106
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13188 9586 13216 11154
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13924 10062 13952 10406
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9722 13860 9930
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8634 12940 8774
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12912 7274 12940 7958
rect 13004 7954 13032 9114
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 5778 12940 7210
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5166 12940 5714
rect 13188 5234 13216 9318
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 6798 13308 8366
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13372 5914 13400 9522
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13464 7750 13492 8298
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13556 6866 13584 8978
rect 13740 8906 13768 9522
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13648 6186 13676 7958
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13740 7274 13768 7375
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13832 6390 13860 9658
rect 13924 8566 13952 9998
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14016 7478 14044 11222
rect 14384 9654 14412 12192
rect 14556 12174 14608 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14004 7336 14056 7342
rect 14056 7296 14136 7324
rect 14004 7278 14056 7284
rect 14108 7206 14136 7296
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6866 14136 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 14292 6254 14320 8910
rect 14384 7954 14412 9590
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13360 5704 13412 5710
rect 13648 5692 13676 6122
rect 14476 5914 14504 12038
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 6730 14596 11290
rect 14660 11082 14688 11630
rect 15304 11218 15332 12174
rect 15580 11830 15608 12854
rect 15672 12306 15700 14010
rect 15764 13326 15792 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15842 13968 15898 13977
rect 15842 13903 15844 13912
rect 15896 13903 15898 13912
rect 15948 13920 15976 14010
rect 16028 13932 16080 13938
rect 15948 13892 16028 13920
rect 15844 13874 15896 13880
rect 16028 13874 16080 13880
rect 16316 13870 16344 15438
rect 16500 15065 16528 25094
rect 16868 24614 16896 25706
rect 17144 25294 17172 26182
rect 17880 25974 17908 27542
rect 18708 27470 18736 29200
rect 21192 27606 21220 29200
rect 23676 27606 23704 29200
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 26160 27606 26188 29200
rect 21180 27600 21232 27606
rect 21180 27542 21232 27548
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 28368 27470 28396 29294
rect 28630 29200 28686 29294
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17972 26042 18000 27338
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 23768 26518 23796 27270
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 18064 25838 18092 26386
rect 26252 26382 26280 27270
rect 28184 26450 28212 27270
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 26240 26376 26292 26382
rect 19522 26344 19578 26353
rect 26240 26318 26292 26324
rect 19522 26279 19524 26288
rect 19576 26279 19578 26288
rect 24952 26308 25004 26314
rect 19524 26250 19576 26256
rect 24952 26250 25004 26256
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 18708 25838 18736 26182
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18708 25702 18736 25774
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17592 25696 17644 25702
rect 18696 25696 18748 25702
rect 17592 25638 17644 25644
rect 18694 25664 18696 25673
rect 18748 25664 18750 25673
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24993 16988 25094
rect 16946 24984 17002 24993
rect 16946 24919 17002 24928
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16592 23866 16620 24346
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16868 23730 16896 24550
rect 17052 23866 17080 24754
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 17236 23730 17264 25638
rect 17604 25294 17632 25638
rect 18315 25596 18623 25605
rect 18694 25599 18750 25608
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 17420 23866 17448 24618
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16868 23322 16896 23666
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 20534 16712 21422
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16592 18766 16620 20470
rect 16776 19145 16804 22374
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16868 21486 16896 21966
rect 16948 21616 17000 21622
rect 17000 21576 17080 21604
rect 16948 21558 17000 21564
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16868 21146 16896 21422
rect 17052 21146 17080 21576
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17236 21010 17264 23666
rect 17420 22574 17448 23802
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17420 21554 17448 22510
rect 17604 21894 17632 24346
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17696 22574 17724 22918
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17236 20330 17264 20946
rect 17696 20806 17724 22510
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 16762 19136 16818 19145
rect 16762 19071 16818 19080
rect 17236 18766 17264 20266
rect 16580 18760 16632 18766
rect 16856 18760 16908 18766
rect 16632 18708 16712 18714
rect 16580 18702 16712 18708
rect 16856 18702 16908 18708
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 16592 18686 16712 18702
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 16590 16620 18566
rect 16684 17814 16712 18686
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16776 17746 16804 18090
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16658 16712 17070
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16578 15328 16634 15337
rect 16578 15263 16634 15272
rect 16486 15056 16542 15065
rect 16486 14991 16542 15000
rect 16500 14346 16528 14991
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16120 13864 16172 13870
rect 15948 13812 16120 13818
rect 15948 13806 16172 13812
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 15948 13802 16160 13806
rect 15936 13796 16160 13802
rect 15988 13790 16160 13796
rect 15936 13738 15988 13744
rect 16592 13530 16620 15263
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15764 12170 15792 13262
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12918 16344 13194
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16592 12646 16620 13330
rect 16684 12714 16712 16594
rect 16776 16250 16804 17138
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16868 15042 16896 18702
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16960 16250 16988 16730
rect 17236 16590 17264 16934
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17420 16182 17448 17478
rect 17512 16454 17540 18634
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 16948 16108 17000 16114
rect 17224 16108 17276 16114
rect 17000 16068 17224 16096
rect 16948 16050 17000 16056
rect 17224 16050 17276 16056
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 17052 15144 17080 15914
rect 17052 15116 17356 15144
rect 16776 15014 16896 15042
rect 16948 15020 17000 15026
rect 16776 14822 16804 15014
rect 17132 15020 17184 15026
rect 16948 14962 17000 14968
rect 17052 14980 17132 15008
rect 16856 14952 16908 14958
rect 16960 14929 16988 14962
rect 16856 14894 16908 14900
rect 16946 14920 17002 14929
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16868 14482 16896 14894
rect 16946 14855 17002 14864
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 13841 16896 14418
rect 16960 14074 16988 14554
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16854 13832 16910 13841
rect 16854 13767 16910 13776
rect 16948 13796 17000 13802
rect 17052 13784 17080 14980
rect 17132 14962 17184 14968
rect 17328 14929 17356 15116
rect 17314 14920 17370 14929
rect 17314 14855 17370 14864
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 14074 17264 14214
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17000 13756 17080 13784
rect 16948 13738 17000 13744
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15764 11694 15792 12106
rect 16040 11830 16068 12242
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14660 8634 14688 11018
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14660 7886 14688 8026
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 13412 5664 13676 5692
rect 13360 5646 13412 5652
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 5030 14228 5102
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13004 4622 13032 4694
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 13372 3738 13400 4422
rect 14200 4146 14228 4966
rect 14568 4146 14596 6666
rect 14660 6458 14688 7822
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 5914 14780 9930
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 8906 15056 9386
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 15108 8560 15160 8566
rect 15212 8514 15240 10066
rect 15160 8508 15240 8514
rect 15108 8502 15240 8508
rect 15120 8486 15240 8502
rect 15106 7984 15162 7993
rect 15106 7919 15108 7928
rect 15160 7919 15162 7928
rect 15108 7890 15160 7896
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 15304 7342 15332 10542
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15856 9178 15884 9454
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15384 8832 15436 8838
rect 15382 8800 15384 8809
rect 15476 8832 15528 8838
rect 15436 8800 15438 8809
rect 15476 8774 15528 8780
rect 15382 8735 15438 8744
rect 15488 8498 15516 8774
rect 15764 8514 15792 8978
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15948 8634 15976 8842
rect 16040 8634 16068 9862
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15672 8486 15792 8514
rect 15672 8430 15700 8486
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14844 5710 14872 6258
rect 15028 5710 15056 6394
rect 14832 5704 14884 5710
rect 14752 5664 14832 5692
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 12176 2530 12204 3402
rect 12268 3058 12296 3674
rect 14660 3602 14688 4626
rect 14752 4622 14780 5664
rect 14832 5646 14884 5652
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 15304 5302 15332 7278
rect 15948 6798 15976 8570
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 6322 16068 6598
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 5846 15884 6190
rect 15948 5914 15976 6258
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12176 2514 12572 2530
rect 12176 2508 12584 2514
rect 12176 2502 12532 2508
rect 12532 2450 12584 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 11624 800 11652 2246
rect 12728 800 12756 2790
rect 13004 2514 13032 3334
rect 13832 2514 13860 3538
rect 14660 2854 14688 3538
rect 15304 3534 15332 3946
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 15488 2446 15516 5510
rect 15672 3942 15700 5714
rect 16040 5234 16068 6054
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4690 16252 4966
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16408 4146 16436 9318
rect 16592 8616 16620 12582
rect 16776 12238 16804 12718
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16868 11354 16896 11630
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16684 10266 16712 10542
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16500 8588 16620 8616
rect 16500 7546 16528 8588
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16592 6934 16620 8366
rect 16684 7818 16712 9862
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16684 6254 16712 7210
rect 16776 6730 16804 7754
rect 16868 7546 16896 8230
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16868 6798 16896 7482
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16960 6390 16988 13738
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 7324 17080 9998
rect 17144 8906 17172 13942
rect 17328 13938 17356 14855
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 12170 17264 13738
rect 17604 12442 17632 17682
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 14006 17724 15370
rect 17788 14618 17816 25094
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 19444 24818 19564 24834
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19432 24812 19564 24818
rect 19484 24806 19564 24812
rect 19432 24754 19484 24760
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23118 17908 24006
rect 17972 23798 18000 24754
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18064 24206 18092 24686
rect 18236 24676 18288 24682
rect 18236 24618 18288 24624
rect 18052 24200 18104 24206
rect 18104 24160 18184 24188
rect 18052 24142 18104 24148
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17972 23322 18000 23734
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17880 22642 17908 23054
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 18064 22438 18092 23598
rect 18156 23322 18184 24160
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 22094 18092 22374
rect 18156 22234 18184 23122
rect 18248 22778 18276 24618
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18708 24206 18736 24754
rect 18880 24676 18932 24682
rect 18880 24618 18932 24624
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23866 18552 24006
rect 18708 23866 18736 24142
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 18248 22506 18276 22714
rect 18708 22574 18736 22986
rect 18800 22778 18828 24550
rect 18892 24206 18920 24618
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18984 23594 19012 24550
rect 19260 24206 19288 24754
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19260 23662 19288 24142
rect 19444 24070 19472 24618
rect 19536 24138 19564 24806
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 19628 24410 19656 24754
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 21284 24274 21312 24754
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19524 24132 19576 24138
rect 19576 24092 19656 24120
rect 19524 24074 19576 24080
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 19444 23322 19472 24006
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19248 23248 19300 23254
rect 19248 23190 19300 23196
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18144 22228 18196 22234
rect 18196 22188 18276 22216
rect 18144 22170 18196 22176
rect 18064 22066 18184 22094
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17880 20058 17908 21898
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17972 18970 18000 21558
rect 18156 20942 18184 22066
rect 18248 21690 18276 22188
rect 19168 22166 19196 22578
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19260 21706 19288 23190
rect 19536 23186 19564 23462
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19340 23112 19392 23118
rect 19628 23100 19656 24092
rect 20088 23730 20116 24142
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 19708 23112 19760 23118
rect 19628 23072 19708 23100
rect 19340 23054 19392 23060
rect 19708 23054 19760 23060
rect 19352 22438 19380 23054
rect 19720 22710 19748 23054
rect 20272 22982 20300 23666
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 22098 19380 22374
rect 19444 22234 19472 22646
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 19168 21678 19288 21706
rect 18248 20942 18276 21626
rect 19168 21350 19196 21678
rect 19352 21604 19380 21898
rect 19260 21576 19380 21604
rect 19260 21486 19288 21576
rect 19444 21554 19472 22170
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19536 21622 19564 22102
rect 19524 21616 19576 21622
rect 19524 21558 19576 21564
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 19260 20874 19288 21422
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 18052 20868 18104 20874
rect 19248 20868 19300 20874
rect 18052 20810 18104 20816
rect 19168 20828 19248 20856
rect 18064 20262 18092 20810
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17880 18086 17908 18226
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17972 17746 18000 18702
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 14890 17908 15982
rect 18064 15502 18092 20198
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18156 16046 18184 18226
rect 18248 17882 18276 20742
rect 19168 20534 19196 20828
rect 19248 20810 19300 20816
rect 19156 20528 19208 20534
rect 19156 20470 19208 20476
rect 19352 20466 19380 21354
rect 19628 20466 19656 22102
rect 20180 22098 20208 22510
rect 20272 22166 20300 22918
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19812 21690 19840 21966
rect 19904 21690 19932 21966
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 20180 21622 20208 22034
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19340 20460 19392 20466
rect 19260 20420 19340 20448
rect 19260 20380 19288 20420
rect 19340 20402 19392 20408
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19076 20352 19288 20380
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18420 19848 18472 19854
rect 18512 19848 18564 19854
rect 18420 19790 18472 19796
rect 18510 19816 18512 19825
rect 18564 19816 18566 19825
rect 18432 19378 18460 19790
rect 19076 19786 19104 20352
rect 19444 19854 19472 20402
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 18510 19751 18566 19760
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18708 18970 18736 19314
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18708 18766 18736 18906
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18326 17776 18382 17785
rect 18326 17711 18382 17720
rect 18340 17678 18368 17711
rect 18708 17678 18736 18158
rect 18800 17728 18828 19654
rect 19076 19514 19104 19722
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19444 19446 19472 19654
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18290 18920 18702
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18984 17746 19012 19110
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18972 17740 19024 17746
rect 18800 17700 18920 17728
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18892 17610 18920 17700
rect 18972 17682 19024 17688
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16794 18276 16934
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18708 16794 18736 17206
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18248 16522 18276 16730
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18694 16144 18750 16153
rect 18694 16079 18696 16088
rect 18748 16079 18750 16088
rect 18696 16050 18748 16056
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18512 15564 18564 15570
rect 18800 15552 18828 17546
rect 18512 15506 18564 15512
rect 18708 15524 18828 15552
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18248 15094 18276 15370
rect 18326 15192 18382 15201
rect 18326 15127 18382 15136
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 18248 14822 18276 15030
rect 18340 15026 18368 15127
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18524 14890 18552 15506
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 18156 14482 18184 14758
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18248 14362 18276 14758
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18432 14414 18460 14486
rect 18616 14414 18644 14554
rect 18420 14408 18472 14414
rect 18248 14346 18368 14362
rect 18420 14350 18472 14356
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18144 14340 18196 14346
rect 18248 14340 18380 14346
rect 18248 14334 18328 14340
rect 18144 14282 18196 14288
rect 18328 14282 18380 14288
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 18064 12918 18092 14282
rect 18156 12918 18184 14282
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13326 18276 14214
rect 18616 13818 18644 14350
rect 18708 14346 18736 15524
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18800 15026 18828 15370
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 14618 18828 14826
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18892 14414 18920 15302
rect 19076 14550 19104 18566
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19168 14940 19196 17546
rect 19260 17338 19288 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 18222 19380 19246
rect 19536 18358 19564 20198
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19628 19854 19656 19994
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19352 17134 19380 18158
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19536 17542 19564 17750
rect 19628 17678 19656 19314
rect 19812 18834 19840 20742
rect 19904 20466 19932 21082
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19904 18970 19932 19790
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19996 18766 20024 21286
rect 20088 21010 20116 21354
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20088 20058 20116 20946
rect 20364 20806 20392 21898
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20456 20466 20484 23666
rect 21284 23526 21312 24006
rect 21468 23798 21496 24550
rect 21560 24206 21588 24686
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22112 24342 22140 24550
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 21456 23792 21508 23798
rect 21456 23734 21508 23740
rect 22204 23730 22232 24074
rect 22296 24018 22324 24686
rect 22480 24682 22508 24754
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22468 24676 22520 24682
rect 22468 24618 22520 24624
rect 22480 24206 22508 24618
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 24274 22784 24550
rect 23124 24410 23152 24686
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22296 23990 22508 24018
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22296 23769 22324 23802
rect 22282 23760 22338 23769
rect 22192 23724 22244 23730
rect 22388 23730 22416 23802
rect 22282 23695 22338 23704
rect 22376 23724 22428 23730
rect 22192 23666 22244 23672
rect 22376 23666 22428 23672
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21088 23248 21140 23254
rect 21088 23190 21140 23196
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20548 22710 20576 23122
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 22778 21036 23054
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20548 22094 20576 22646
rect 20640 22234 20668 22646
rect 21100 22574 21128 23190
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22710 21220 22918
rect 21284 22778 21312 23462
rect 21916 23112 21968 23118
rect 22204 23066 22232 23666
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22296 23118 22324 23598
rect 21968 23060 22232 23066
rect 21916 23054 22232 23060
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22388 23066 22416 23666
rect 22480 23594 22508 23990
rect 22664 23662 22692 24142
rect 22756 23730 22784 24210
rect 23216 23866 23244 24210
rect 23308 23866 23336 24754
rect 24492 24676 24544 24682
rect 24492 24618 24544 24624
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23388 24132 23440 24138
rect 23388 24074 23440 24080
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22468 23588 22520 23594
rect 22468 23530 22520 23536
rect 22480 23338 22508 23530
rect 22480 23310 22600 23338
rect 22756 23322 22784 23666
rect 23216 23526 23244 23802
rect 23204 23520 23256 23526
rect 23204 23462 23256 23468
rect 21928 23038 22232 23054
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20548 22066 20668 22094
rect 20640 22030 20668 22066
rect 21100 22030 21128 22510
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21546 21992 21602 22001
rect 20548 20942 20576 21966
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20640 21554 20668 21830
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 20466 20576 20742
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 20330 20576 20402
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20548 19922 20576 20266
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 19854 20668 21286
rect 20732 20466 20760 21558
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20824 19990 20852 21966
rect 21376 21622 21404 21966
rect 21546 21927 21602 21936
rect 21364 21616 21416 21622
rect 21364 21558 21416 21564
rect 21376 20874 21404 21558
rect 21560 21078 21588 21927
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21560 20466 21588 21014
rect 21652 20942 21680 22918
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 22296 22760 22324 23054
rect 22388 23050 22508 23066
rect 22388 23044 22520 23050
rect 22388 23038 22468 23044
rect 22468 22986 22520 22992
rect 22572 22778 22600 23310
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 23216 23118 23244 23462
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23400 22778 23428 24074
rect 23492 23662 23520 24142
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23730 23612 24006
rect 23662 23760 23718 23769
rect 23572 23724 23624 23730
rect 23768 23730 23796 24074
rect 24504 23730 24532 24618
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24688 24274 24716 24550
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 23662 23695 23718 23704
rect 23756 23724 23808 23730
rect 23572 23666 23624 23672
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23676 23050 23704 23695
rect 23756 23666 23808 23672
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23860 23118 23888 23462
rect 23848 23112 23900 23118
rect 23768 23072 23848 23100
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 21928 22732 22324 22760
rect 22560 22772 22612 22778
rect 21928 22234 21956 22732
rect 22560 22714 22612 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22204 22234 22232 22578
rect 23676 22574 23704 22986
rect 23768 22642 23796 23072
rect 23848 23054 23900 23060
rect 24504 22642 24532 23666
rect 24596 23186 24624 23666
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 24872 23118 24900 24006
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 21914 21992 21970 22001
rect 21914 21927 21916 21936
rect 21968 21927 21970 21936
rect 21916 21898 21968 21904
rect 22112 21876 22140 22102
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 22468 21888 22520 21894
rect 22112 21848 22232 21876
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20916 19786 20944 20334
rect 21652 20330 21680 20878
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 21192 19514 21220 19926
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21192 19378 21220 19450
rect 21272 19440 21324 19446
rect 21272 19382 21324 19388
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19904 18426 19932 18702
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19628 17270 19656 17614
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19890 17232 19946 17241
rect 20088 17202 20116 17614
rect 19890 17167 19892 17176
rect 19944 17167 19946 17176
rect 20076 17196 20128 17202
rect 19892 17138 19944 17144
rect 20076 17138 20128 17144
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19812 16590 19840 17070
rect 19800 16584 19852 16590
rect 20088 16538 20116 17138
rect 19800 16526 19852 16532
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 14958 19380 15846
rect 19444 15570 19472 16390
rect 19812 16046 19840 16526
rect 19904 16510 20116 16538
rect 19904 16454 19932 16510
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19904 16114 19932 16390
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 20088 16046 20116 16390
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19720 15638 19748 15846
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 15026 19564 15302
rect 20088 15162 20116 15506
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19982 15056 20038 15065
rect 19524 15020 19576 15026
rect 19982 14991 19984 15000
rect 19524 14962 19576 14968
rect 20036 14991 20038 15000
rect 20076 15020 20128 15026
rect 19984 14962 20036 14968
rect 20076 14962 20128 14968
rect 19248 14952 19300 14958
rect 19168 14912 19248 14940
rect 19248 14894 19300 14900
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18708 13938 18736 14282
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18800 13841 18828 14214
rect 18892 13938 18920 14350
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18786 13832 18842 13841
rect 18616 13790 18736 13818
rect 18708 13682 18736 13790
rect 18786 13767 18842 13776
rect 19062 13832 19118 13841
rect 19062 13767 19118 13776
rect 18708 13654 18828 13682
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18248 12850 18276 13262
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17696 12238 17724 12786
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17972 12238 18000 12718
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18064 12345 18092 12582
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18708 12442 18736 12582
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18050 12336 18106 12345
rect 18050 12271 18106 12280
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17420 10810 17448 11766
rect 17788 11558 17816 12038
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9722 17264 10066
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17144 8634 17172 8842
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17236 8430 17264 9658
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9042 17356 9318
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17420 8634 17448 10134
rect 17788 9586 17816 11494
rect 17880 11218 18000 11234
rect 17880 11212 18012 11218
rect 17880 11206 17960 11212
rect 17880 9722 17908 11206
rect 17960 11154 18012 11160
rect 18064 11150 18092 12271
rect 18144 12164 18196 12170
rect 18144 12106 18196 12112
rect 18156 11830 18184 12106
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17972 10470 18000 11018
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17224 8424 17276 8430
rect 17420 8401 17448 8570
rect 17224 8366 17276 8372
rect 17406 8392 17462 8401
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 8022 17172 8230
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17132 7336 17184 7342
rect 17052 7296 17132 7324
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16500 4486 16528 5578
rect 16684 5302 16712 6190
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15580 3194 15608 3878
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15948 2650 15976 3470
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16040 2582 16068 3130
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 2038 12940 2246
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 13832 800 13860 2314
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 15304 1442 15332 2314
rect 16132 2310 16160 3878
rect 16316 3738 16344 4082
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 2650 16344 3334
rect 16500 3126 16528 4422
rect 16592 3534 16620 4422
rect 16776 4078 16804 6326
rect 17052 4622 17080 7296
rect 17132 7278 17184 7284
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 6866 17172 7142
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17236 6254 17264 8366
rect 17406 8327 17462 8336
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17420 7324 17448 7482
rect 17500 7336 17552 7342
rect 17420 7296 17500 7324
rect 17500 7278 17552 7284
rect 17406 6760 17462 6769
rect 17604 6746 17632 8978
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17788 8634 17816 8910
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17972 8022 18000 10406
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9722 18092 9998
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9110 18184 9318
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18052 8492 18104 8498
rect 18248 8480 18276 12038
rect 18800 11830 18828 13654
rect 18972 12096 19024 12102
rect 18892 12056 18972 12084
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18708 9994 18736 11494
rect 18892 10674 18920 12056
rect 18972 12038 19024 12044
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 18604 9580 18656 9586
rect 18656 9540 18736 9568
rect 18604 9522 18656 9528
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18104 8452 18276 8480
rect 18328 8492 18380 8498
rect 18052 8434 18104 8440
rect 18328 8434 18380 8440
rect 18340 8378 18368 8434
rect 18248 8350 18368 8378
rect 18248 8090 18276 8350
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 17960 8016 18012 8022
rect 18144 8016 18196 8022
rect 17960 7958 18012 7964
rect 18142 7984 18144 7993
rect 18196 7984 18198 7993
rect 18142 7919 18198 7928
rect 18248 7818 18276 8026
rect 18708 7886 18736 9540
rect 18892 9178 18920 10610
rect 19076 9654 19104 13767
rect 19260 12850 19288 14894
rect 20088 14822 20116 14962
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 13938 19932 14350
rect 19892 13932 19944 13938
rect 19944 13892 20024 13920
rect 19892 13874 19944 13880
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12986 19472 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19168 11082 19196 11698
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18800 7886 18828 9046
rect 18892 8090 18920 9114
rect 18984 8566 19012 9522
rect 19168 9178 19196 9590
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19062 8800 19118 8809
rect 19062 8735 19118 8744
rect 19076 8566 19104 8735
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 19076 7478 19104 8366
rect 19168 8294 19196 9114
rect 19260 9110 19288 11018
rect 19352 10470 19380 12582
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11898 19472 12242
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19628 11354 19656 13398
rect 19720 13394 19748 13806
rect 19996 13462 20024 13892
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19708 13388 19760 13394
rect 19760 13348 19932 13376
rect 19708 13330 19760 13336
rect 19800 11824 19852 11830
rect 19798 11792 19800 11801
rect 19852 11792 19854 11801
rect 19904 11762 19932 13348
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12238 20024 13126
rect 20088 12306 20116 14486
rect 20180 13734 20208 18226
rect 20456 17814 20484 19110
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17338 20392 17478
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20364 17202 20392 17274
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 16114 20300 16594
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20272 14958 20300 16050
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15026 20392 15438
rect 20456 15162 20484 17750
rect 20548 17746 20576 19110
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 18306 20760 18770
rect 20824 18766 20852 19246
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20812 18624 20864 18630
rect 20916 18612 20944 18770
rect 20864 18584 20944 18612
rect 20812 18566 20864 18572
rect 20732 18278 20944 18306
rect 21100 18290 21128 19178
rect 21284 18408 21312 19382
rect 21192 18380 21312 18408
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20548 17610 20576 17682
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20732 16590 20760 18158
rect 20812 16992 20864 16998
rect 20916 16980 20944 18278
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20994 17232 21050 17241
rect 20994 17167 21050 17176
rect 20864 16952 20944 16980
rect 20812 16934 20864 16940
rect 20824 16590 20852 16934
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 13802 20392 14214
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20272 12238 20300 13262
rect 20364 13258 20392 13738
rect 20456 13462 20484 14282
rect 20548 14006 20576 16526
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20640 15706 20668 16390
rect 20732 16130 20760 16526
rect 21008 16454 21036 17167
rect 21100 16726 21128 18226
rect 21192 18086 21220 18380
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21284 17882 21312 18226
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21376 17814 21404 19654
rect 21468 18714 21496 20266
rect 21652 19922 21680 20266
rect 22020 19990 22048 20402
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 22204 19854 22232 21848
rect 22468 21830 22520 21836
rect 22480 21418 22508 21830
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 23032 20942 23060 21422
rect 23124 20942 23152 21490
rect 23492 21026 23520 21626
rect 23400 21010 23520 21026
rect 23584 21010 23612 22034
rect 23676 22030 23704 22510
rect 23768 22234 23796 22578
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23952 22098 23980 22578
rect 24872 22574 24900 23054
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 24596 22030 24624 22374
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24688 21570 24716 22374
rect 24872 22234 24900 22510
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24780 21690 24808 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24412 21554 24716 21570
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 24400 21548 24716 21554
rect 24452 21542 24716 21548
rect 24400 21490 24452 21496
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23676 21146 23704 21354
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23388 21004 23520 21010
rect 23440 20998 23520 21004
rect 23572 21004 23624 21010
rect 23388 20946 23440 20952
rect 23572 20946 23624 20952
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23032 20262 23060 20878
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22204 19378 22232 19790
rect 22572 19446 22600 20198
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 21468 18686 21680 18714
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21284 17270 21312 17682
rect 21272 17264 21324 17270
rect 21270 17232 21272 17241
rect 21376 17252 21404 17750
rect 21468 17746 21496 18686
rect 21652 18630 21680 18686
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21560 18426 21588 18566
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21560 17678 21588 18362
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21548 17536 21600 17542
rect 21652 17524 21680 18158
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 21600 17496 21680 17524
rect 21548 17478 21600 17484
rect 21456 17264 21508 17270
rect 21324 17232 21326 17241
rect 21376 17224 21456 17252
rect 21456 17206 21508 17212
rect 21270 17167 21326 17176
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21192 16522 21220 16934
rect 21376 16794 21404 17070
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20732 16102 20852 16130
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 15337 20668 15438
rect 20626 15328 20682 15337
rect 20626 15263 20682 15272
rect 20732 15162 20760 15982
rect 20824 15366 20852 16102
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20824 15201 20852 15302
rect 20810 15192 20866 15201
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20720 15156 20772 15162
rect 20810 15127 20866 15136
rect 20720 15098 20772 15104
rect 20640 14006 20668 15098
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 14074 20760 14350
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20456 12374 20484 13398
rect 20732 13394 20760 13806
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20824 13274 20852 14962
rect 20916 14822 20944 15914
rect 21192 15706 21220 16050
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21284 15502 21312 16662
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21272 15020 21324 15026
rect 21376 15008 21404 16730
rect 21468 15026 21496 17002
rect 21560 16658 21588 17478
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22204 17338 22232 17614
rect 22296 17610 22324 18090
rect 22388 17678 22416 18226
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21560 16182 21588 16594
rect 21652 16590 21680 17138
rect 21744 16998 21772 17138
rect 22296 17066 22324 17546
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16590 22416 16934
rect 22480 16658 22508 17478
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22572 16590 22600 19382
rect 22756 18766 22784 19790
rect 23032 19310 23060 20198
rect 23308 20058 23336 20878
rect 23400 20874 23428 20946
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23400 20482 23428 20810
rect 23492 20602 23520 20878
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23400 20454 23520 20482
rect 23584 20466 23612 20946
rect 23860 20806 23888 21490
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23492 19854 23520 20454
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23480 19848 23532 19854
rect 23532 19796 23612 19802
rect 23480 19790 23612 19796
rect 23492 19774 23612 19790
rect 23676 19786 23704 20538
rect 23860 20398 23888 20742
rect 24596 20466 24624 21542
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24688 21146 24716 21422
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24780 20602 24808 21626
rect 24872 20942 24900 21898
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 24044 20058 24072 20402
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 23860 19854 23888 19994
rect 24596 19938 24624 20402
rect 24412 19910 24624 19938
rect 24412 19854 24440 19910
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 23584 19718 23612 19774
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 23388 19712 23440 19718
rect 23572 19712 23624 19718
rect 23440 19660 23520 19666
rect 23388 19654 23520 19660
rect 23572 19654 23624 19660
rect 23400 19638 23520 19654
rect 23492 19310 23520 19638
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 24320 19242 24348 19722
rect 24596 19514 24624 19790
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24872 19446 24900 19722
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23584 18834 23612 19110
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22848 17338 22876 17478
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 21652 16250 21680 16526
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 21560 15570 21588 15982
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21560 15434 21588 15506
rect 21652 15502 21680 15914
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 22388 15162 22416 15982
rect 22480 15638 22508 16050
rect 22572 15910 22600 16118
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 21324 14980 21404 15008
rect 21456 15020 21508 15026
rect 21272 14962 21324 14968
rect 21456 14962 21508 14968
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 13530 20944 14758
rect 21100 14414 21128 14826
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20732 13246 20852 13274
rect 20732 12986 20760 13246
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20720 12980 20772 12986
rect 20640 12940 20720 12968
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19798 11727 19854 11736
rect 19892 11756 19944 11762
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19812 11082 19840 11727
rect 19892 11698 19944 11704
rect 19996 11626 20024 11766
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10674 19472 10950
rect 19904 10810 19932 11290
rect 19996 11218 20024 11562
rect 20076 11552 20128 11558
rect 20074 11520 20076 11529
rect 20128 11520 20130 11529
rect 20074 11455 20130 11464
rect 20272 11354 20300 12174
rect 20548 12102 20576 12786
rect 20640 12322 20668 12940
rect 20720 12922 20772 12928
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20732 12442 20760 12786
rect 20824 12594 20852 13126
rect 21468 12850 21496 13670
rect 21560 13326 21588 14350
rect 22020 14346 22048 15030
rect 22572 15026 22600 15846
rect 22664 15450 22692 17206
rect 22848 17082 22876 17274
rect 23032 17202 23060 18702
rect 24504 18698 24532 19246
rect 24872 18834 24900 19382
rect 24860 18828 24912 18834
rect 24860 18770 24912 18776
rect 23756 18692 23808 18698
rect 23756 18634 23808 18640
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23216 18290 23244 18566
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23400 17134 23428 17614
rect 23584 17542 23612 18362
rect 23768 18222 23796 18634
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 24308 18080 24360 18086
rect 24308 18022 24360 18028
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23768 17134 23796 17546
rect 23860 17202 23888 17682
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17202 23980 17478
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 22756 17066 22876 17082
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 22744 17060 22876 17066
rect 22796 17054 22876 17060
rect 22744 17002 22796 17008
rect 23952 16590 23980 17138
rect 24320 16794 24348 18022
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24780 17270 24808 17614
rect 24872 17610 24900 18770
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24872 17202 24900 17546
rect 24860 17196 24912 17202
rect 24964 17184 24992 26250
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25148 23050 25176 23462
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25412 22976 25464 22982
rect 25608 22964 25636 23666
rect 25464 22936 25636 22964
rect 25780 22976 25832 22982
rect 25412 22918 25464 22924
rect 25780 22918 25832 22924
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 25056 22522 25084 22918
rect 25424 22710 25452 22918
rect 25412 22704 25464 22710
rect 25412 22646 25464 22652
rect 25792 22642 25820 22918
rect 26056 22704 26108 22710
rect 26056 22646 26108 22652
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25596 22568 25648 22574
rect 25056 22494 25176 22522
rect 25596 22510 25648 22516
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25056 22030 25084 22170
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25148 21690 25176 22494
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25608 21962 25636 22510
rect 25792 22030 25820 22578
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25148 21554 25176 21626
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25608 21350 25636 21898
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25608 21078 25636 21286
rect 25596 21072 25648 21078
rect 25596 21014 25648 21020
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25608 20058 25636 20878
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25608 19854 25636 19994
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 26068 19514 26096 22646
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26252 21418 26280 22510
rect 26344 22030 26372 22918
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26436 22166 26464 22374
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27172 21554 27200 21830
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 20942 26372 21286
rect 27172 21146 27200 21490
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 27264 20942 27292 21490
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 26332 20936 26384 20942
rect 26608 20936 26660 20942
rect 26384 20896 26608 20924
rect 26332 20878 26384 20884
rect 26608 20878 26660 20884
rect 27252 20936 27304 20942
rect 27436 20936 27488 20942
rect 27304 20896 27384 20924
rect 27252 20878 27304 20884
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 25056 18902 25084 19314
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 25056 18766 25084 18838
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25056 18290 25084 18702
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 24964 17156 25176 17184
rect 24860 17138 24912 17144
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24768 16992 24820 16998
rect 24820 16952 24900 16980
rect 24768 16934 24820 16940
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 22756 16182 22784 16390
rect 23124 16250 23152 16390
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22756 15570 22784 16118
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22664 15422 22784 15450
rect 22756 15026 22784 15422
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22848 14890 22876 15982
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22940 14822 22968 15846
rect 23400 15638 23428 16526
rect 23388 15632 23440 15638
rect 23388 15574 23440 15580
rect 23492 15570 23520 16526
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23492 15094 23520 15506
rect 23584 15502 23612 16390
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 13546 21680 14214
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 21652 13518 21772 13546
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 20996 12640 21048 12646
rect 20824 12588 20996 12594
rect 20824 12582 21048 12588
rect 20824 12566 21036 12582
rect 20720 12436 20772 12442
rect 20824 12434 20852 12566
rect 20824 12406 21128 12434
rect 20720 12378 20772 12384
rect 20640 12294 20760 12322
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19706 10568 19762 10577
rect 19706 10503 19762 10512
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19260 8022 19288 8434
rect 19352 8362 19380 8774
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 17462 6718 17632 6746
rect 17406 6695 17408 6704
rect 17460 6695 17462 6704
rect 17408 6666 17460 6672
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17604 5302 17632 6718
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17972 5710 18000 5850
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17236 4282 17264 4966
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 18156 3534 18184 6394
rect 18708 6322 18736 7142
rect 19352 6730 19380 7958
rect 19444 7954 19472 8434
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19444 7546 19472 7754
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6390 18920 6598
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18248 5710 18276 6258
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18432 5302 18460 5714
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18708 5234 18736 6258
rect 18892 5710 18920 6326
rect 19076 6254 19104 6326
rect 19260 6254 19288 6394
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19076 5914 19104 6190
rect 19444 5914 19472 6190
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19536 5846 19564 10406
rect 19720 10266 19748 10503
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19812 9722 19840 9862
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19904 9450 19932 9998
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19628 5778 19656 8774
rect 19904 8634 19932 9386
rect 19996 8906 20024 11154
rect 20272 11150 20300 11290
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 9994 20208 10950
rect 20272 10470 20300 11086
rect 20548 10674 20576 12038
rect 20732 11014 20760 12294
rect 21100 12238 21128 12406
rect 21284 12238 21312 12786
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21468 12238 21496 12650
rect 21560 12345 21588 13126
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20824 11529 20852 11562
rect 20810 11520 20866 11529
rect 20810 11455 20866 11464
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 21100 10810 21128 12174
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20916 10554 20944 10746
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 10600 21048 10606
rect 20916 10548 20996 10554
rect 20916 10542 21048 10548
rect 20916 10526 21036 10542
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20916 10062 20944 10526
rect 20904 10056 20956 10062
rect 20640 10004 20904 10010
rect 20640 9998 20956 10004
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20640 9982 20944 9998
rect 20996 9988 21048 9994
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 20088 8294 20116 9318
rect 20272 8974 20300 9862
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20640 8498 20668 9982
rect 20996 9930 21048 9936
rect 20902 9208 20958 9217
rect 20902 9143 20904 9152
rect 20956 9143 20958 9152
rect 20904 9114 20956 9120
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20902 8392 20958 8401
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19904 7410 19932 8230
rect 20732 7954 20760 8366
rect 21008 8378 21036 9930
rect 21100 9518 21128 10610
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21192 10062 21220 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8906 21128 9318
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20958 8350 21036 8378
rect 21100 8378 21128 8842
rect 21192 8498 21220 9998
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21100 8362 21220 8378
rect 21100 8356 21232 8362
rect 21100 8350 21180 8356
rect 20902 8327 20958 8336
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20456 6390 20484 6734
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20720 6656 20772 6662
rect 20640 6604 20720 6610
rect 20640 6598 20772 6604
rect 20640 6582 20760 6598
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 17328 3058 17356 3334
rect 19352 3058 19380 5034
rect 19444 4622 19472 5102
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4214 19472 4558
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19536 3194 19564 3538
rect 19628 3398 19656 3878
rect 19720 3534 19748 6054
rect 20456 5914 20484 6326
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19904 5370 19932 5510
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19996 5030 20024 5714
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4690 20024 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16316 2446 16344 2586
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 14936 1414 15332 1442
rect 14936 800 14964 1414
rect 16040 870 16160 898
rect 16040 800 16068 870
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3882 0 3938 800
rect 4986 0 5042 800
rect 6090 0 6146 800
rect 7194 0 7250 800
rect 8298 0 8354 800
rect 9402 0 9458 800
rect 10506 0 10562 800
rect 11610 0 11666 800
rect 12714 0 12770 800
rect 13818 0 13874 800
rect 14922 0 14978 800
rect 16026 0 16082 800
rect 16132 762 16160 870
rect 16408 762 16436 2246
rect 17144 800 17172 2790
rect 18156 2310 18184 2790
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18892 2650 18920 2994
rect 19536 2666 19564 3130
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 19260 2638 19564 2666
rect 19260 2530 19288 2638
rect 19168 2502 19288 2530
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19168 2446 19196 2502
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18248 800 18276 2314
rect 19260 2310 19288 2382
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19352 800 19380 2518
rect 19628 2446 19656 3334
rect 19996 3194 20024 4150
rect 20088 4146 20116 5782
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20180 3670 20208 5714
rect 20640 5710 20668 6582
rect 20824 6390 20852 6666
rect 20916 6458 20944 8327
rect 21180 8298 21232 8304
rect 21192 7886 21220 8298
rect 21284 8022 21312 11086
rect 21376 8906 21404 11630
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 11014 21496 11086
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21468 10146 21496 10950
rect 21560 10810 21588 12271
rect 21652 11354 21680 13518
rect 21744 13326 21772 13518
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 22204 11898 22232 14758
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 13938 22508 14418
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 13938 22968 14214
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22466 13832 22522 13841
rect 22466 13767 22522 13776
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22388 12442 22416 12854
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22190 11792 22246 11801
rect 22480 11762 22508 13767
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23124 13326 23152 13670
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 22572 12850 22600 13262
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22190 11727 22192 11736
rect 22244 11727 22246 11736
rect 22468 11756 22520 11762
rect 22192 11698 22244 11704
rect 22468 11698 22520 11704
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 22112 11150 22140 11630
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 10266 21588 10406
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21744 10146 21772 10202
rect 21468 10118 21772 10146
rect 21560 9722 21588 10118
rect 21836 10062 21864 10746
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21652 9722 21680 9930
rect 22204 9926 22232 11494
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10538 22324 10950
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22388 9926 22416 10610
rect 22572 10577 22600 12650
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22558 10568 22614 10577
rect 22664 10538 22692 12038
rect 22756 11626 22784 12786
rect 23124 12238 23152 13262
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23216 12986 23244 13194
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23400 12434 23428 14758
rect 23584 14618 23612 15302
rect 23676 15162 23704 16050
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23860 15502 23888 15982
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23952 15026 23980 15302
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 24320 14618 24348 16730
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24780 16182 24808 16526
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24872 16046 24900 16952
rect 24964 16522 24992 17002
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 16114 24992 16458
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24964 15502 24992 15846
rect 25148 15706 25176 17156
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25608 16658 25636 18158
rect 25700 17882 25728 18770
rect 25884 18766 25912 19314
rect 25964 19236 26016 19242
rect 25964 19178 26016 19184
rect 25976 18766 26004 19178
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25700 17082 25728 17818
rect 25792 17746 25820 18634
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25884 17678 25912 18702
rect 25976 18290 26004 18702
rect 26068 18698 26096 19314
rect 26160 19310 26188 19722
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25976 17882 26004 18226
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25872 17672 25924 17678
rect 26160 17660 26188 19246
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26252 18222 26280 19110
rect 26344 18902 26372 20334
rect 26528 18902 26556 20402
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 19666 27108 20198
rect 27172 19854 27200 20742
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27264 19718 27292 20742
rect 27356 20534 27384 20896
rect 27436 20878 27488 20884
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27160 19712 27212 19718
rect 27080 19660 27160 19666
rect 27080 19654 27212 19660
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27080 19638 27200 19654
rect 27172 19174 27200 19638
rect 27356 19446 27384 19858
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 27356 18970 27384 19382
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 26332 18896 26384 18902
rect 26332 18838 26384 18844
rect 26516 18896 26568 18902
rect 26516 18838 26568 18844
rect 26344 18290 26372 18838
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26436 17882 26464 18770
rect 26528 18766 26556 18838
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 27172 17678 27200 18566
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27264 17882 27292 18158
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 26240 17672 26292 17678
rect 26160 17632 26240 17660
rect 25872 17614 25924 17620
rect 26240 17614 26292 17620
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27344 17196 27396 17202
rect 27448 17184 27476 20878
rect 27540 19514 27568 20878
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 20330 27660 20742
rect 27724 20602 27752 21286
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 27896 19780 27948 19786
rect 27896 19722 27948 19728
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27908 19378 27936 19722
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27896 18148 27948 18154
rect 27896 18090 27948 18096
rect 27908 17202 27936 18090
rect 27396 17156 27476 17184
rect 27344 17138 27396 17144
rect 25700 17054 25820 17082
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25700 16726 25728 16934
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25608 16182 25636 16594
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25608 15994 25636 16118
rect 25700 16114 25728 16662
rect 25792 16590 25820 17054
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25792 16164 25820 16526
rect 26700 16516 26752 16522
rect 26700 16458 26752 16464
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 25964 16176 26016 16182
rect 25792 16136 25964 16164
rect 25964 16118 26016 16124
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25964 16040 26016 16046
rect 25608 15966 25728 15994
rect 25964 15982 26016 15988
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25700 15706 25728 15966
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25608 15502 25636 15574
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24780 15094 24808 15370
rect 25608 15162 25636 15438
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 25700 15094 25728 15642
rect 25792 15502 25820 15846
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25976 15094 26004 15982
rect 26068 15366 26096 16390
rect 26608 16176 26660 16182
rect 26608 16118 26660 16124
rect 26620 15502 26648 16118
rect 26712 16114 26740 16458
rect 27080 16454 27108 16934
rect 27448 16590 27476 17156
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 26976 16448 27028 16454
rect 26976 16390 27028 16396
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26988 15706 27016 16390
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 25688 15088 25740 15094
rect 25688 15030 25740 15036
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 26620 15026 26648 15438
rect 26988 15094 27016 15642
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 27172 15026 27200 16526
rect 27448 16250 27476 16526
rect 27632 16250 27660 16934
rect 27804 16788 27856 16794
rect 27908 16776 27936 17138
rect 27856 16748 27936 16776
rect 27804 16730 27856 16736
rect 28000 16658 28028 20198
rect 28092 20058 28120 20878
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27632 15570 27660 16186
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27724 15706 27752 15982
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27344 15564 27396 15570
rect 27344 15506 27396 15512
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27356 15162 27384 15506
rect 28000 15502 28028 16594
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28080 15972 28132 15978
rect 28080 15914 28132 15920
rect 28092 15706 28120 15914
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 28356 14952 28408 14958
rect 28354 14920 28356 14929
rect 28408 14920 28410 14929
rect 28354 14855 28410 14864
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24596 14618 24624 14758
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 12850 23704 14486
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24412 13530 24440 14282
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24504 12850 24532 14214
rect 24596 13938 24624 14350
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24964 13734 24992 14350
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13138 24992 13670
rect 25056 13462 25084 13874
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 25148 13410 25176 13670
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25056 13274 25084 13398
rect 25148 13382 25268 13410
rect 25056 13258 25176 13274
rect 25056 13252 25188 13258
rect 25056 13246 25136 13252
rect 25136 13194 25188 13200
rect 24964 13110 25084 13138
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 23860 12442 23888 12718
rect 23308 12406 23428 12434
rect 23848 12436 23900 12442
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22558 10503 22614 10512
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21640 9716 21692 9722
rect 22204 9704 22232 9862
rect 21640 9658 21692 9664
rect 22112 9676 22232 9704
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 9110 21864 9318
rect 21732 9104 21784 9110
rect 21652 9064 21732 9092
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21364 8900 21416 8906
rect 21364 8842 21416 8848
rect 21468 8294 21496 8978
rect 21652 8498 21680 9064
rect 21732 9046 21784 9052
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 22112 8974 22140 9676
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 22204 8634 22232 9318
rect 22296 9178 22324 9454
rect 22480 9217 22508 9930
rect 22664 9654 22692 10202
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22466 9208 22522 9217
rect 22284 9172 22336 9178
rect 22466 9143 22522 9152
rect 22284 9114 22336 9120
rect 22572 9110 22600 9522
rect 22756 9450 22784 11562
rect 22848 11354 22876 11834
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 23124 11218 23152 12174
rect 23308 12170 23336 12406
rect 24412 12434 24440 12718
rect 23848 12378 23900 12384
rect 24136 12406 24440 12434
rect 24136 12306 24164 12406
rect 24780 12306 24808 12786
rect 25056 12646 25084 13110
rect 25240 12714 25268 13382
rect 25608 13326 25636 13874
rect 25872 13388 25924 13394
rect 25872 13330 25924 13336
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25332 12986 25360 13262
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25700 12782 25728 13126
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22848 9450 22876 9998
rect 22940 9586 22968 10678
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23308 10577 23336 10610
rect 23294 10568 23350 10577
rect 23294 10503 23350 10512
rect 23112 10192 23164 10198
rect 23112 10134 23164 10140
rect 23124 9586 23152 10134
rect 23308 9674 23336 10503
rect 23400 10062 23428 12038
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23492 10130 23520 11698
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23400 9926 23428 9998
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23216 9646 23336 9674
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23216 9450 23244 9646
rect 22744 9444 22796 9450
rect 22744 9386 22796 9392
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22756 9330 22784 9386
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 21008 6254 21036 7686
rect 21100 6322 21128 7754
rect 21560 7274 21588 7822
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22296 7478 22324 7754
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22572 7410 22600 9046
rect 22664 8838 22692 9318
rect 22756 9302 22876 9330
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 7818 22692 8774
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22756 7410 22784 9114
rect 22848 8498 22876 9302
rect 23216 9178 23244 9386
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23400 9110 23428 9862
rect 23584 9602 23612 11154
rect 23676 11150 23704 11494
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23676 10538 23704 11086
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23768 10606 23796 10950
rect 24136 10742 24164 12242
rect 24964 12238 24992 12582
rect 25056 12374 25084 12582
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25412 12368 25464 12374
rect 25412 12310 25464 12316
rect 25424 12238 25452 12310
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23492 9574 23612 9602
rect 23492 9518 23520 9574
rect 23952 9518 23980 9930
rect 24136 9926 24164 10678
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23940 9512 23992 9518
rect 23940 9454 23992 9460
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23388 9104 23440 9110
rect 23308 9064 23388 9092
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8566 23244 8774
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 23308 7954 23336 9064
rect 23388 9046 23440 9052
rect 23492 8974 23520 9318
rect 23570 9208 23626 9217
rect 23570 9143 23626 9152
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23400 8090 23428 8910
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23584 7546 23612 9143
rect 23860 9042 23888 9318
rect 24044 9042 24072 9522
rect 24136 9450 24164 9590
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24136 8634 24164 9386
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24136 8090 24164 8570
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24228 8022 24256 11018
rect 24320 10606 24348 11154
rect 24412 11150 24440 11562
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24596 10810 24624 12106
rect 24688 11354 24716 12106
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11354 24900 11630
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24768 11144 24820 11150
rect 25056 11132 25084 12174
rect 25608 12170 25636 12718
rect 25136 12164 25188 12170
rect 25136 12106 25188 12112
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25148 11354 25176 12106
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25240 11830 25268 12038
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 24768 11086 24820 11092
rect 24964 11104 25084 11132
rect 25136 11144 25188 11150
rect 24584 10804 24636 10810
rect 24584 10746 24636 10752
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 9586 24624 10542
rect 24688 10266 24716 10610
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24688 9722 24716 10202
rect 24780 9994 24808 11086
rect 24964 10470 24992 11104
rect 25136 11086 25188 11092
rect 25688 11144 25740 11150
rect 25792 11132 25820 12786
rect 25884 11694 25912 13330
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25976 12918 26004 13262
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25964 12708 26016 12714
rect 25964 12650 26016 12656
rect 25976 12238 26004 12650
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 25740 11104 25820 11132
rect 25872 11144 25924 11150
rect 25688 11086 25740 11092
rect 25976 11132 26004 11834
rect 26068 11762 26096 12922
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 25924 11104 26004 11132
rect 25872 11086 25924 11092
rect 25148 11014 25176 11086
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24872 10062 24900 10406
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24596 8430 24624 9522
rect 24688 9178 24716 9522
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24780 9110 24808 9454
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24780 8498 24808 9046
rect 24872 8906 24900 9998
rect 24964 9450 24992 10406
rect 25148 10266 25176 10950
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 25056 9722 25084 9930
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 25056 9217 25084 9658
rect 25148 9586 25176 10202
rect 25884 10198 25912 11086
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 26160 10266 26188 10678
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 25872 10192 25924 10198
rect 25872 10134 25924 10140
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25042 9208 25098 9217
rect 25261 9211 25569 9220
rect 25608 9178 25636 9862
rect 25884 9722 25912 10134
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 26252 9518 26280 9862
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 25042 9143 25098 9152
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 25148 8430 25176 8774
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 22572 6798 22600 7346
rect 22756 7206 22784 7346
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20640 5166 20668 5646
rect 21008 5642 21036 6190
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 21008 5234 21036 5578
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20272 2514 20300 3878
rect 20364 3738 20392 4558
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4146 20576 4490
rect 20640 4282 20668 4966
rect 21008 4622 21036 5170
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20732 3738 20760 4150
rect 20916 4078 20944 4422
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 20456 800 20484 2450
rect 20732 2446 20760 3674
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21008 3058 21036 3334
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21376 2854 21404 3946
rect 21468 3466 21496 4422
rect 21652 4214 21680 5170
rect 22204 4622 22232 6122
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22296 5370 22324 5510
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22468 5296 22520 5302
rect 22468 5238 22520 5244
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21640 4208 21692 4214
rect 22204 4162 22232 4558
rect 22296 4214 22324 4966
rect 21640 4150 21692 4156
rect 22020 4146 22232 4162
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22008 4140 22232 4146
rect 22060 4134 22232 4140
rect 22008 4082 22060 4088
rect 22204 3738 22232 4134
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 21468 3058 21496 3402
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 22204 3074 22232 3674
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22112 3058 22232 3074
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 22100 3052 22232 3058
rect 22152 3046 22232 3052
rect 22100 2994 22152 3000
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21468 2582 21496 2994
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 21560 800 21588 2586
rect 22388 2582 22416 3334
rect 22480 3194 22508 5238
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22756 3534 22784 4422
rect 22940 3942 22968 4558
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 23204 4004 23256 4010
rect 23204 3946 23256 3952
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 23110 3768 23166 3777
rect 23110 3703 23112 3712
rect 23164 3703 23166 3712
rect 23112 3674 23164 3680
rect 23216 3618 23244 3946
rect 23400 3754 23428 3946
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23400 3726 23520 3754
rect 23124 3590 23244 3618
rect 23388 3596 23440 3602
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22376 2576 22428 2582
rect 22376 2518 22428 2524
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 22664 800 22692 2790
rect 23124 2774 23152 3590
rect 23388 3538 23440 3544
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 23216 3058 23244 3402
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23124 2746 23244 2774
rect 22928 2576 22980 2582
rect 22980 2524 23152 2530
rect 22928 2518 23152 2524
rect 22940 2514 23152 2518
rect 22940 2508 23164 2514
rect 22940 2502 23112 2508
rect 23112 2450 23164 2456
rect 23216 2446 23244 2746
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23308 2378 23336 3334
rect 23400 2446 23428 3538
rect 23492 3534 23520 3726
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23584 3194 23612 3538
rect 23952 3194 23980 3878
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 23756 2576 23808 2582
rect 23756 2518 23808 2524
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23296 2372 23348 2378
rect 23296 2314 23348 2320
rect 23768 800 23796 2518
rect 23860 2446 23888 3130
rect 24504 2922 24532 4490
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 3126 24624 3334
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 24780 2310 24808 2994
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24872 800 24900 2382
rect 25976 800 26004 2382
rect 27080 800 27108 2382
rect 28184 800 28212 2382
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 29288 800 29316 2926
rect 16132 734 16436 762
rect 17130 0 17186 800
rect 18234 0 18290 800
rect 19338 0 19394 800
rect 20442 0 20498 800
rect 21546 0 21602 800
rect 22650 0 22706 800
rect 23754 0 23810 800
rect 24858 0 24914 800
rect 25962 0 26018 800
rect 27066 0 27122 800
rect 28170 0 28226 800
rect 29274 0 29330 800
<< via2 >>
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4158 26288 4214 26344
rect 1858 19624 1914 19680
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 1950 13776 2006 13832
rect 3330 20476 3332 20496
rect 3332 20476 3384 20496
rect 3384 20476 3386 20496
rect 3330 20440 3386 20476
rect 2502 9424 2558 9480
rect 4710 25100 4712 25120
rect 4712 25100 4764 25120
rect 4764 25100 4766 25120
rect 4710 25064 4766 25100
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4158 19352 4214 19408
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4710 20712 4766 20768
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4434 19488 4490 19544
rect 4802 19488 4858 19544
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4986 17584 5042 17640
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4618 15444 4620 15464
rect 4620 15444 4672 15464
rect 4672 15444 4674 15464
rect 4618 15408 4674 15444
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4434 12688 4490 12744
rect 4710 12844 4766 12880
rect 4710 12824 4712 12844
rect 4712 12824 4764 12844
rect 4764 12824 4766 12844
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 3882 10648 3938 10704
rect 3422 7948 3478 7984
rect 3422 7928 3424 7948
rect 3424 7928 3476 7948
rect 3476 7928 3478 7948
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 5446 20304 5502 20360
rect 5446 19624 5502 19680
rect 5170 12688 5226 12744
rect 5078 12416 5134 12472
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 6458 25200 6514 25256
rect 5078 10920 5134 10976
rect 7654 25200 7710 25256
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 6550 19796 6552 19816
rect 6552 19796 6604 19816
rect 6604 19796 6606 19816
rect 6550 19760 6606 19796
rect 6366 19488 6422 19544
rect 6642 17448 6698 17504
rect 8298 23060 8300 23080
rect 8300 23060 8352 23080
rect 8352 23060 8354 23080
rect 7378 20848 7434 20904
rect 8298 23024 8354 23060
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 5078 8064 5134 8120
rect 5078 7928 5134 7984
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4986 6860 5042 6896
rect 4986 6840 4988 6860
rect 4988 6840 5040 6860
rect 5040 6840 5042 6860
rect 5998 12688 6054 12744
rect 5722 10668 5778 10704
rect 5722 10648 5724 10668
rect 5724 10648 5776 10668
rect 5776 10648 5778 10668
rect 5814 9560 5870 9616
rect 5538 8336 5594 8392
rect 5722 8492 5778 8528
rect 5722 8472 5724 8492
rect 5724 8472 5776 8492
rect 5776 8472 5778 8492
rect 6458 13932 6514 13968
rect 6458 13912 6460 13932
rect 6460 13912 6512 13932
rect 6512 13912 6514 13932
rect 6826 12824 6882 12880
rect 7286 14320 7342 14376
rect 7102 12824 7158 12880
rect 7010 12552 7066 12608
rect 6550 10648 6606 10704
rect 6550 8472 6606 8528
rect 8298 20848 8354 20904
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 8114 20440 8170 20496
rect 7838 20304 7894 20360
rect 8022 20304 8078 20360
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 8666 22616 8722 22672
rect 9402 25200 9458 25256
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 8482 20848 8538 20904
rect 8482 19780 8538 19816
rect 8482 19760 8484 19780
rect 8484 19760 8536 19780
rect 8536 19760 8538 19780
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7930 17620 7932 17640
rect 7932 17620 7984 17640
rect 7984 17620 7986 17640
rect 7930 17584 7986 17620
rect 8390 17620 8392 17640
rect 8392 17620 8444 17640
rect 8444 17620 8446 17640
rect 8390 17584 8446 17620
rect 7746 17448 7802 17504
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7838 15408 7894 15464
rect 8022 15444 8024 15464
rect 8024 15444 8076 15464
rect 8076 15444 8078 15464
rect 8022 15408 8078 15444
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7654 13776 7710 13832
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 7378 12552 7434 12608
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 8666 12416 8722 12472
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 8206 8064 8262 8120
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 9310 20304 9366 20360
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 10874 22480 10930 22536
rect 9126 19352 9182 19408
rect 9218 15408 9274 15464
rect 9126 13912 9182 13968
rect 8942 12416 8998 12472
rect 8850 12280 8906 12336
rect 9862 17040 9918 17096
rect 10046 17040 10102 17096
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11978 22480 12034 22536
rect 12714 22072 12770 22128
rect 11978 20340 11980 20360
rect 11980 20340 12032 20360
rect 12032 20340 12034 20360
rect 11978 20304 12034 20340
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 10230 17040 10286 17096
rect 9494 12280 9550 12336
rect 10138 13776 10194 13832
rect 8574 9036 8630 9072
rect 8574 9016 8576 9036
rect 8576 9016 8628 9036
rect 8628 9016 8630 9036
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 10506 10512 10562 10568
rect 10690 13932 10746 13968
rect 10690 13912 10692 13932
rect 10692 13912 10744 13932
rect 10744 13912 10746 13932
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 10690 11056 10746 11112
rect 10230 6704 10286 6760
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 10966 10684 10968 10704
rect 10968 10684 11020 10704
rect 11020 10684 11022 10704
rect 10966 10648 11022 10684
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11886 12688 11942 12744
rect 12714 19352 12770 19408
rect 12438 14864 12494 14920
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11978 10648 12034 10704
rect 13174 20340 13176 20360
rect 13176 20340 13228 20360
rect 13228 20340 13230 20360
rect 13174 20304 13230 20340
rect 14002 22636 14058 22672
rect 14002 22616 14004 22636
rect 14004 22616 14056 22636
rect 14056 22616 14058 22636
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14462 20712 14518 20768
rect 13634 19352 13690 19408
rect 13542 19116 13544 19136
rect 13544 19116 13596 19136
rect 13596 19116 13598 19136
rect 13542 19080 13598 19116
rect 11886 10512 11942 10568
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 12438 7384 12494 7440
rect 13450 17040 13506 17096
rect 13266 13912 13322 13968
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14830 19760 14886 19816
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 15290 13776 15346 13832
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 15934 22480 15990 22536
rect 13726 7384 13782 7440
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 15842 13932 15898 13968
rect 15842 13912 15844 13932
rect 15844 13912 15896 13932
rect 15896 13912 15898 13932
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 19522 26308 19578 26344
rect 19522 26288 19524 26308
rect 19524 26288 19576 26308
rect 19576 26288 19578 26308
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 18694 25644 18696 25664
rect 18696 25644 18748 25664
rect 18748 25644 18750 25664
rect 16946 24928 17002 24984
rect 18694 25608 18750 25644
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 16762 19080 16818 19136
rect 16578 15272 16634 15328
rect 16486 15000 16542 15056
rect 16946 14864 17002 14920
rect 16854 13776 16910 13832
rect 17314 14864 17370 14920
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 15106 7948 15162 7984
rect 15106 7928 15108 7948
rect 15108 7928 15160 7948
rect 15160 7928 15162 7948
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 15382 8780 15384 8800
rect 15384 8780 15436 8800
rect 15436 8780 15438 8800
rect 15382 8744 15438 8780
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18510 19796 18512 19816
rect 18512 19796 18564 19816
rect 18564 19796 18566 19816
rect 18510 19760 18566 19796
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18326 17720 18382 17776
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18694 16108 18750 16144
rect 18694 16088 18696 16108
rect 18696 16088 18748 16108
rect 18748 16088 18750 16108
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18326 15136 18382 15192
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 22282 23704 22338 23760
rect 21546 21936 21602 21992
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 23662 23704 23718 23760
rect 21914 21956 21970 21992
rect 21914 21936 21916 21956
rect 21916 21936 21968 21956
rect 21968 21936 21970 21956
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 19890 17196 19946 17232
rect 19890 17176 19892 17196
rect 19892 17176 19944 17196
rect 19944 17176 19946 17196
rect 19982 15020 20038 15056
rect 19982 15000 19984 15020
rect 19984 15000 20036 15020
rect 20036 15000 20038 15020
rect 18786 13776 18842 13832
rect 19062 13776 19118 13832
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18050 12280 18106 12336
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 17406 8336 17462 8392
rect 17406 6724 17462 6760
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18142 7964 18144 7984
rect 18144 7964 18196 7984
rect 18196 7964 18198 7984
rect 18142 7928 18198 7964
rect 19062 8744 19118 8800
rect 19798 11772 19800 11792
rect 19800 11772 19852 11792
rect 19852 11772 19854 11792
rect 19798 11736 19854 11772
rect 20994 17176 21050 17232
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21270 17212 21272 17232
rect 21272 17212 21324 17232
rect 21324 17212 21326 17232
rect 21270 17176 21326 17212
rect 20626 15272 20682 15328
rect 20810 15136 20866 15192
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 20074 11500 20076 11520
rect 20076 11500 20128 11520
rect 20128 11500 20130 11520
rect 20074 11464 20130 11500
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 19706 10512 19762 10568
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 17406 6704 17408 6724
rect 17408 6704 17460 6724
rect 17460 6704 17462 6724
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 21546 12280 21602 12336
rect 20810 11464 20866 11520
rect 20902 9172 20958 9208
rect 20902 9152 20904 9172
rect 20904 9152 20956 9172
rect 20956 9152 20958 9172
rect 20902 8336 20958 8392
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 22466 13776 22522 13832
rect 22190 11756 22246 11792
rect 22190 11736 22192 11756
rect 22192 11736 22244 11756
rect 22244 11736 22246 11756
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 22558 10512 22614 10568
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28354 14900 28356 14920
rect 28356 14900 28408 14920
rect 28408 14900 28410 14920
rect 28354 14864 28410 14900
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 22466 9152 22522 9208
rect 23294 10512 23350 10568
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 23570 9152 23626 9208
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25042 9152 25098 9208
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 23110 3732 23166 3768
rect 23110 3712 23112 3732
rect 23112 3712 23164 3732
rect 23164 3712 23166 3732
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 4153 26346 4219 26349
rect 19517 26348 19583 26349
rect 6126 26346 6132 26348
rect 4153 26344 6132 26346
rect 4153 26288 4158 26344
rect 4214 26288 6132 26344
rect 4153 26286 6132 26288
rect 4153 26283 4219 26286
rect 6126 26284 6132 26286
rect 6196 26284 6202 26348
rect 19517 26344 19564 26348
rect 19628 26346 19634 26348
rect 19517 26288 19522 26344
rect 19517 26284 19564 26288
rect 19628 26286 19674 26346
rect 19628 26284 19634 26286
rect 19517 26283 19583 26284
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 18689 25666 18755 25669
rect 18822 25666 18828 25668
rect 18689 25664 18828 25666
rect 18689 25608 18694 25664
rect 18750 25608 18828 25664
rect 18689 25606 18828 25608
rect 18689 25603 18755 25606
rect 18822 25604 18828 25606
rect 18892 25604 18898 25668
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 6453 25258 6519 25261
rect 7649 25258 7715 25261
rect 9397 25258 9463 25261
rect 6453 25256 9463 25258
rect 6453 25200 6458 25256
rect 6514 25200 7654 25256
rect 7710 25200 9402 25256
rect 9458 25200 9463 25256
rect 6453 25198 9463 25200
rect 6453 25195 6519 25198
rect 7649 25195 7715 25198
rect 9397 25195 9463 25198
rect 4705 25122 4771 25125
rect 5022 25122 5028 25124
rect 4705 25120 5028 25122
rect 4705 25064 4710 25120
rect 4766 25064 5028 25120
rect 4705 25062 5028 25064
rect 4705 25059 4771 25062
rect 5022 25060 5028 25062
rect 5092 25060 5098 25124
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 16941 24988 17007 24989
rect 16941 24984 16988 24988
rect 17052 24986 17058 24988
rect 16941 24928 16946 24984
rect 16941 24924 16988 24928
rect 17052 24926 17098 24986
rect 17052 24924 17058 24926
rect 16941 24923 17007 24924
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 22277 23762 22343 23765
rect 23657 23762 23723 23765
rect 22277 23760 23723 23762
rect 22277 23704 22282 23760
rect 22338 23704 23662 23760
rect 23718 23704 23723 23760
rect 22277 23702 23723 23704
rect 22277 23699 22343 23702
rect 23657 23699 23723 23702
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 5022 23020 5028 23084
rect 5092 23082 5098 23084
rect 8293 23082 8359 23085
rect 5092 23080 8359 23082
rect 5092 23024 8298 23080
rect 8354 23024 8359 23080
rect 5092 23022 8359 23024
rect 5092 23020 5098 23022
rect 8293 23019 8359 23022
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 8661 22674 8727 22677
rect 13997 22674 14063 22677
rect 8661 22672 14063 22674
rect 8661 22616 8666 22672
rect 8722 22616 14002 22672
rect 14058 22616 14063 22672
rect 8661 22614 14063 22616
rect 8661 22611 8727 22614
rect 13997 22611 14063 22614
rect 10869 22538 10935 22541
rect 11973 22538 12039 22541
rect 15929 22538 15995 22541
rect 10869 22536 15995 22538
rect 10869 22480 10874 22536
rect 10930 22480 11978 22536
rect 12034 22480 15934 22536
rect 15990 22480 15995 22536
rect 10869 22478 15995 22480
rect 10869 22475 10935 22478
rect 11973 22475 12039 22478
rect 15929 22475 15995 22478
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 12709 22132 12775 22133
rect 12709 22128 12756 22132
rect 12820 22130 12826 22132
rect 12709 22072 12714 22128
rect 12709 22068 12756 22072
rect 12820 22070 12866 22130
rect 12820 22068 12826 22070
rect 12709 22067 12775 22068
rect 21541 21994 21607 21997
rect 21909 21994 21975 21997
rect 21541 21992 21975 21994
rect 21541 21936 21546 21992
rect 21602 21936 21914 21992
rect 21970 21936 21975 21992
rect 21541 21934 21975 21936
rect 21541 21931 21607 21934
rect 21909 21931 21975 21934
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 7373 20906 7439 20909
rect 8293 20906 8359 20909
rect 8477 20906 8543 20909
rect 7373 20904 8543 20906
rect 7373 20848 7378 20904
rect 7434 20848 8298 20904
rect 8354 20848 8482 20904
rect 8538 20848 8543 20904
rect 7373 20846 8543 20848
rect 7373 20843 7439 20846
rect 8293 20843 8359 20846
rect 8477 20843 8543 20846
rect 4705 20770 4771 20773
rect 5022 20770 5028 20772
rect 4705 20768 5028 20770
rect 4705 20712 4710 20768
rect 4766 20712 5028 20768
rect 4705 20710 5028 20712
rect 4705 20707 4771 20710
rect 5022 20708 5028 20710
rect 5092 20708 5098 20772
rect 14457 20770 14523 20773
rect 14590 20770 14596 20772
rect 14457 20768 14596 20770
rect 14457 20712 14462 20768
rect 14518 20712 14596 20768
rect 14457 20710 14596 20712
rect 14457 20707 14523 20710
rect 14590 20708 14596 20710
rect 14660 20708 14666 20772
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 3325 20498 3391 20501
rect 8109 20498 8175 20501
rect 3325 20496 8175 20498
rect 3325 20440 3330 20496
rect 3386 20440 8114 20496
rect 8170 20440 8175 20496
rect 3325 20438 8175 20440
rect 3325 20435 3391 20438
rect 8109 20435 8175 20438
rect 5441 20362 5507 20365
rect 7833 20362 7899 20365
rect 5441 20360 7899 20362
rect 5441 20304 5446 20360
rect 5502 20304 7838 20360
rect 7894 20304 7899 20360
rect 5441 20302 7899 20304
rect 5441 20299 5507 20302
rect 7833 20299 7899 20302
rect 8017 20362 8083 20365
rect 9305 20362 9371 20365
rect 8017 20360 9371 20362
rect 8017 20304 8022 20360
rect 8078 20304 9310 20360
rect 9366 20304 9371 20360
rect 8017 20302 9371 20304
rect 8017 20299 8083 20302
rect 9305 20299 9371 20302
rect 11973 20362 12039 20365
rect 13169 20362 13235 20365
rect 11973 20360 13235 20362
rect 11973 20304 11978 20360
rect 12034 20304 13174 20360
rect 13230 20304 13235 20360
rect 11973 20302 13235 20304
rect 11973 20299 12039 20302
rect 13169 20299 13235 20302
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 6545 19818 6611 19821
rect 8477 19818 8543 19821
rect 6545 19816 8543 19818
rect 6545 19760 6550 19816
rect 6606 19760 8482 19816
rect 8538 19760 8543 19816
rect 6545 19758 8543 19760
rect 6545 19755 6611 19758
rect 8477 19755 8543 19758
rect 14825 19818 14891 19821
rect 18505 19818 18571 19821
rect 14825 19816 18571 19818
rect 14825 19760 14830 19816
rect 14886 19760 18510 19816
rect 18566 19760 18571 19816
rect 14825 19758 18571 19760
rect 14825 19755 14891 19758
rect 18505 19755 18571 19758
rect 1853 19682 1919 19685
rect 5441 19682 5507 19685
rect 1853 19680 5507 19682
rect 1853 19624 1858 19680
rect 1914 19624 5446 19680
rect 5502 19624 5507 19680
rect 1853 19622 5507 19624
rect 1853 19619 1919 19622
rect 5441 19619 5507 19622
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 4429 19546 4495 19549
rect 4797 19546 4863 19549
rect 6361 19546 6427 19549
rect 4429 19544 6427 19546
rect 4429 19488 4434 19544
rect 4490 19488 4802 19544
rect 4858 19488 6366 19544
rect 6422 19488 6427 19544
rect 4429 19486 6427 19488
rect 4429 19483 4495 19486
rect 4797 19483 4863 19486
rect 6361 19483 6427 19486
rect 4153 19410 4219 19413
rect 9121 19410 9187 19413
rect 4153 19408 9187 19410
rect 4153 19352 4158 19408
rect 4214 19352 9126 19408
rect 9182 19352 9187 19408
rect 4153 19350 9187 19352
rect 4153 19347 4219 19350
rect 9121 19347 9187 19350
rect 12709 19410 12775 19413
rect 13629 19412 13695 19413
rect 13486 19410 13492 19412
rect 12709 19408 13492 19410
rect 12709 19352 12714 19408
rect 12770 19352 13492 19408
rect 12709 19350 13492 19352
rect 12709 19347 12775 19350
rect 13486 19348 13492 19350
rect 13556 19348 13562 19412
rect 13629 19408 13676 19412
rect 13740 19410 13746 19412
rect 13629 19352 13634 19408
rect 13629 19348 13676 19352
rect 13740 19350 13786 19410
rect 13740 19348 13746 19350
rect 13629 19347 13695 19348
rect 13537 19138 13603 19141
rect 16757 19138 16823 19141
rect 13537 19136 16823 19138
rect 13537 19080 13542 19136
rect 13598 19080 16762 19136
rect 16818 19080 16823 19136
rect 13537 19078 16823 19080
rect 13537 19075 13603 19078
rect 16757 19075 16823 19078
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 14590 17716 14596 17780
rect 14660 17778 14666 17780
rect 18321 17778 18387 17781
rect 14660 17776 18387 17778
rect 14660 17720 18326 17776
rect 18382 17720 18387 17776
rect 14660 17718 18387 17720
rect 14660 17716 14666 17718
rect 18321 17715 18387 17718
rect 4981 17642 5047 17645
rect 7925 17642 7991 17645
rect 4981 17640 7991 17642
rect 4981 17584 4986 17640
rect 5042 17584 7930 17640
rect 7986 17584 7991 17640
rect 4981 17582 7991 17584
rect 4981 17579 5047 17582
rect 7925 17579 7991 17582
rect 8385 17642 8451 17645
rect 8518 17642 8524 17644
rect 8385 17640 8524 17642
rect 8385 17584 8390 17640
rect 8446 17584 8524 17640
rect 8385 17582 8524 17584
rect 8385 17579 8451 17582
rect 8518 17580 8524 17582
rect 8588 17580 8594 17644
rect 6637 17506 6703 17509
rect 7741 17506 7807 17509
rect 6637 17504 7807 17506
rect 6637 17448 6642 17504
rect 6698 17448 7746 17504
rect 7802 17448 7807 17504
rect 6637 17446 7807 17448
rect 6637 17443 6703 17446
rect 7741 17443 7807 17446
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 19885 17234 19951 17237
rect 20989 17234 21055 17237
rect 21265 17234 21331 17237
rect 19885 17232 21331 17234
rect 19885 17176 19890 17232
rect 19946 17176 20994 17232
rect 21050 17176 21270 17232
rect 21326 17176 21331 17232
rect 19885 17174 21331 17176
rect 19885 17171 19951 17174
rect 20989 17171 21055 17174
rect 21265 17171 21331 17174
rect 9857 17098 9923 17101
rect 10041 17098 10107 17101
rect 9857 17096 10107 17098
rect 9857 17040 9862 17096
rect 9918 17040 10046 17096
rect 10102 17040 10107 17096
rect 9857 17038 10107 17040
rect 9857 17035 9923 17038
rect 10041 17035 10107 17038
rect 10225 17098 10291 17101
rect 13445 17098 13511 17101
rect 10225 17096 13511 17098
rect 10225 17040 10230 17096
rect 10286 17040 13450 17096
rect 13506 17040 13511 17096
rect 10225 17038 13511 17040
rect 10225 17035 10291 17038
rect 13445 17035 13511 17038
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 13486 16084 13492 16148
rect 13556 16146 13562 16148
rect 18689 16146 18755 16149
rect 13556 16144 18755 16146
rect 13556 16088 18694 16144
rect 18750 16088 18755 16144
rect 13556 16086 18755 16088
rect 13556 16084 13562 16086
rect 18689 16083 18755 16086
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 4613 15466 4679 15469
rect 5022 15466 5028 15468
rect 4613 15464 5028 15466
rect 4613 15408 4618 15464
rect 4674 15408 5028 15464
rect 4613 15406 5028 15408
rect 4613 15403 4679 15406
rect 5022 15404 5028 15406
rect 5092 15404 5098 15468
rect 7414 15404 7420 15468
rect 7484 15466 7490 15468
rect 7833 15466 7899 15469
rect 7484 15464 7899 15466
rect 7484 15408 7838 15464
rect 7894 15408 7899 15464
rect 7484 15406 7899 15408
rect 7484 15404 7490 15406
rect 7833 15403 7899 15406
rect 8017 15466 8083 15469
rect 9213 15466 9279 15469
rect 8017 15464 9279 15466
rect 8017 15408 8022 15464
rect 8078 15408 9218 15464
rect 9274 15408 9279 15464
rect 8017 15406 9279 15408
rect 8017 15403 8083 15406
rect 9213 15403 9279 15406
rect 16573 15330 16639 15333
rect 16982 15330 16988 15332
rect 16573 15328 16988 15330
rect 16573 15272 16578 15328
rect 16634 15272 16988 15328
rect 16573 15270 16988 15272
rect 16573 15267 16639 15270
rect 16982 15268 16988 15270
rect 17052 15330 17058 15332
rect 20621 15330 20687 15333
rect 17052 15328 20687 15330
rect 17052 15272 20626 15328
rect 20682 15272 20687 15328
rect 17052 15270 20687 15272
rect 17052 15268 17058 15270
rect 20621 15267 20687 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 18321 15194 18387 15197
rect 19558 15194 19564 15196
rect 18321 15192 19564 15194
rect 18321 15136 18326 15192
rect 18382 15136 19564 15192
rect 18321 15134 19564 15136
rect 18321 15131 18387 15134
rect 19558 15132 19564 15134
rect 19628 15132 19634 15196
rect 20805 15194 20871 15197
rect 20670 15192 20871 15194
rect 20670 15136 20810 15192
rect 20866 15136 20871 15192
rect 20670 15134 20871 15136
rect 16481 15058 16547 15061
rect 19977 15058 20043 15061
rect 16481 15056 20043 15058
rect 16481 15000 16486 15056
rect 16542 15000 19982 15056
rect 20038 15000 20043 15056
rect 16481 14998 20043 15000
rect 16481 14995 16547 14998
rect 19977 14995 20043 14998
rect 12433 14922 12499 14925
rect 16941 14922 17007 14925
rect 12433 14920 17007 14922
rect 12433 14864 12438 14920
rect 12494 14864 16946 14920
rect 17002 14864 17007 14920
rect 12433 14862 17007 14864
rect 12433 14859 12499 14862
rect 16941 14859 17007 14862
rect 17309 14922 17375 14925
rect 20670 14922 20730 15134
rect 20805 15131 20871 15134
rect 17309 14920 20730 14922
rect 17309 14864 17314 14920
rect 17370 14864 20730 14920
rect 17309 14862 20730 14864
rect 28349 14922 28415 14925
rect 29200 14922 30000 14952
rect 28349 14920 30000 14922
rect 28349 14864 28354 14920
rect 28410 14864 30000 14920
rect 28349 14862 30000 14864
rect 17309 14859 17375 14862
rect 28349 14859 28415 14862
rect 29200 14832 30000 14862
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 7281 14378 7347 14381
rect 12750 14378 12756 14380
rect 7281 14376 12756 14378
rect 7281 14320 7286 14376
rect 7342 14320 12756 14376
rect 7281 14318 12756 14320
rect 7281 14315 7347 14318
rect 12750 14316 12756 14318
rect 12820 14316 12826 14380
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 6453 13970 6519 13973
rect 9121 13970 9187 13973
rect 6453 13968 9187 13970
rect 6453 13912 6458 13968
rect 6514 13912 9126 13968
rect 9182 13912 9187 13968
rect 6453 13910 9187 13912
rect 6453 13907 6519 13910
rect 9121 13907 9187 13910
rect 10685 13970 10751 13973
rect 13261 13970 13327 13973
rect 10685 13968 13327 13970
rect 10685 13912 10690 13968
rect 10746 13912 13266 13968
rect 13322 13912 13327 13968
rect 10685 13910 13327 13912
rect 10685 13907 10751 13910
rect 13261 13907 13327 13910
rect 13670 13908 13676 13972
rect 13740 13970 13746 13972
rect 15837 13970 15903 13973
rect 13740 13968 15903 13970
rect 13740 13912 15842 13968
rect 15898 13912 15903 13968
rect 13740 13910 15903 13912
rect 13740 13908 13746 13910
rect 15837 13907 15903 13910
rect 1945 13834 2011 13837
rect 7649 13834 7715 13837
rect 1945 13832 7715 13834
rect 1945 13776 1950 13832
rect 2006 13776 7654 13832
rect 7710 13776 7715 13832
rect 1945 13774 7715 13776
rect 1945 13771 2011 13774
rect 7649 13771 7715 13774
rect 10133 13834 10199 13837
rect 15285 13834 15351 13837
rect 16849 13834 16915 13837
rect 10133 13832 16915 13834
rect 10133 13776 10138 13832
rect 10194 13776 15290 13832
rect 15346 13776 16854 13832
rect 16910 13776 16915 13832
rect 10133 13774 16915 13776
rect 10133 13771 10199 13774
rect 15285 13771 15351 13774
rect 16849 13771 16915 13774
rect 18781 13834 18847 13837
rect 19057 13834 19123 13837
rect 22461 13834 22527 13837
rect 18781 13832 22527 13834
rect 18781 13776 18786 13832
rect 18842 13776 19062 13832
rect 19118 13776 22466 13832
rect 22522 13776 22527 13832
rect 18781 13774 22527 13776
rect 18781 13771 18847 13774
rect 19057 13771 19123 13774
rect 22461 13771 22527 13774
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 4705 12882 4771 12885
rect 6821 12882 6887 12885
rect 7097 12882 7163 12885
rect 4705 12880 7163 12882
rect 4705 12824 4710 12880
rect 4766 12824 6826 12880
rect 6882 12824 7102 12880
rect 7158 12824 7163 12880
rect 4705 12822 7163 12824
rect 4705 12819 4771 12822
rect 6821 12819 6887 12822
rect 7097 12819 7163 12822
rect 4429 12746 4495 12749
rect 5165 12746 5231 12749
rect 5993 12746 6059 12749
rect 6310 12746 6316 12748
rect 4429 12744 6316 12746
rect 4429 12688 4434 12744
rect 4490 12688 5170 12744
rect 5226 12688 5998 12744
rect 6054 12688 6316 12744
rect 4429 12686 6316 12688
rect 4429 12683 4495 12686
rect 5165 12683 5231 12686
rect 5993 12683 6059 12686
rect 6310 12684 6316 12686
rect 6380 12746 6386 12748
rect 11881 12746 11947 12749
rect 6380 12744 11947 12746
rect 6380 12688 11886 12744
rect 11942 12688 11947 12744
rect 6380 12686 11947 12688
rect 6380 12684 6386 12686
rect 11881 12683 11947 12686
rect 7005 12610 7071 12613
rect 7373 12610 7439 12613
rect 7005 12608 7439 12610
rect 7005 12552 7010 12608
rect 7066 12552 7378 12608
rect 7434 12552 7439 12608
rect 7005 12550 7439 12552
rect 7005 12547 7071 12550
rect 7373 12547 7439 12550
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 5073 12474 5139 12477
rect 8661 12474 8727 12477
rect 8937 12474 9003 12477
rect 5073 12472 9003 12474
rect 5073 12416 5078 12472
rect 5134 12416 8666 12472
rect 8722 12416 8942 12472
rect 8998 12416 9003 12472
rect 5073 12414 9003 12416
rect 5073 12411 5139 12414
rect 8661 12411 8727 12414
rect 8937 12411 9003 12414
rect 8845 12338 8911 12341
rect 9489 12338 9555 12341
rect 8845 12336 9555 12338
rect 8845 12280 8850 12336
rect 8906 12280 9494 12336
rect 9550 12280 9555 12336
rect 8845 12278 9555 12280
rect 8845 12275 8911 12278
rect 9489 12275 9555 12278
rect 18045 12338 18111 12341
rect 21541 12338 21607 12341
rect 18045 12336 21607 12338
rect 18045 12280 18050 12336
rect 18106 12280 21546 12336
rect 21602 12280 21607 12336
rect 18045 12278 21607 12280
rect 18045 12275 18111 12278
rect 21541 12275 21607 12278
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 19793 11794 19859 11797
rect 22185 11794 22251 11797
rect 19793 11792 22251 11794
rect 19793 11736 19798 11792
rect 19854 11736 22190 11792
rect 22246 11736 22251 11792
rect 19793 11734 22251 11736
rect 19793 11731 19859 11734
rect 22185 11731 22251 11734
rect 20069 11522 20135 11525
rect 20805 11522 20871 11525
rect 20069 11520 20871 11522
rect 20069 11464 20074 11520
rect 20130 11464 20810 11520
rect 20866 11464 20871 11520
rect 20069 11462 20871 11464
rect 20069 11459 20135 11462
rect 20805 11459 20871 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 8518 11114 8524 11116
rect 5582 11054 8524 11114
rect 4102 10916 4108 10980
rect 4172 10978 4178 10980
rect 5073 10978 5139 10981
rect 5582 10978 5642 11054
rect 8518 11052 8524 11054
rect 8588 11114 8594 11116
rect 10685 11114 10751 11117
rect 8588 11112 10751 11114
rect 8588 11056 10690 11112
rect 10746 11056 10751 11112
rect 8588 11054 10751 11056
rect 8588 11052 8594 11054
rect 10685 11051 10751 11054
rect 4172 10976 5642 10978
rect 4172 10920 5078 10976
rect 5134 10920 5642 10976
rect 4172 10918 5642 10920
rect 4172 10916 4178 10918
rect 5073 10915 5139 10918
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 3877 10706 3943 10709
rect 5717 10706 5783 10709
rect 6545 10706 6611 10709
rect 3877 10704 6611 10706
rect 3877 10648 3882 10704
rect 3938 10648 5722 10704
rect 5778 10648 6550 10704
rect 6606 10648 6611 10704
rect 3877 10646 6611 10648
rect 3877 10643 3943 10646
rect 5717 10643 5783 10646
rect 6545 10643 6611 10646
rect 10961 10706 11027 10709
rect 11973 10706 12039 10709
rect 10961 10704 12039 10706
rect 10961 10648 10966 10704
rect 11022 10648 11978 10704
rect 12034 10648 12039 10704
rect 10961 10646 12039 10648
rect 10961 10643 11027 10646
rect 11973 10643 12039 10646
rect 10501 10570 10567 10573
rect 11881 10570 11947 10573
rect 10501 10568 11947 10570
rect 10501 10512 10506 10568
rect 10562 10512 11886 10568
rect 11942 10512 11947 10568
rect 10501 10510 11947 10512
rect 10501 10507 10567 10510
rect 11881 10507 11947 10510
rect 19701 10570 19767 10573
rect 22553 10570 22619 10573
rect 23289 10570 23355 10573
rect 19701 10568 23355 10570
rect 19701 10512 19706 10568
rect 19762 10512 22558 10568
rect 22614 10512 23294 10568
rect 23350 10512 23355 10568
rect 19701 10510 23355 10512
rect 19701 10507 19767 10510
rect 22553 10507 22619 10510
rect 23289 10507 23355 10510
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 5809 9618 5875 9621
rect 6310 9618 6316 9620
rect 5809 9616 6316 9618
rect 5809 9560 5814 9616
rect 5870 9560 6316 9616
rect 5809 9558 6316 9560
rect 5809 9555 5875 9558
rect 6310 9556 6316 9558
rect 6380 9556 6386 9620
rect 2497 9482 2563 9485
rect 7414 9482 7420 9484
rect 2497 9480 7420 9482
rect 2497 9424 2502 9480
rect 2558 9424 7420 9480
rect 2497 9422 7420 9424
rect 2497 9419 2563 9422
rect 7414 9420 7420 9422
rect 7484 9420 7490 9484
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 20897 9210 20963 9213
rect 22461 9210 22527 9213
rect 23565 9210 23631 9213
rect 25037 9210 25103 9213
rect 20897 9208 25103 9210
rect 20897 9152 20902 9208
rect 20958 9152 22466 9208
rect 22522 9152 23570 9208
rect 23626 9152 25042 9208
rect 25098 9152 25103 9208
rect 20897 9150 25103 9152
rect 20897 9147 20963 9150
rect 22461 9147 22527 9150
rect 23565 9147 23631 9150
rect 25037 9147 25103 9150
rect 6126 9012 6132 9076
rect 6196 9074 6202 9076
rect 8569 9074 8635 9077
rect 6196 9072 8635 9074
rect 6196 9016 8574 9072
rect 8630 9016 8635 9072
rect 6196 9014 8635 9016
rect 6196 9012 6202 9014
rect 8569 9011 8635 9014
rect 15377 8802 15443 8805
rect 19057 8802 19123 8805
rect 15377 8800 19123 8802
rect 15377 8744 15382 8800
rect 15438 8744 19062 8800
rect 19118 8744 19123 8800
rect 15377 8742 19123 8744
rect 15377 8739 15443 8742
rect 19057 8739 19123 8742
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 5717 8530 5783 8533
rect 6545 8530 6611 8533
rect 5717 8528 6611 8530
rect 5717 8472 5722 8528
rect 5778 8472 6550 8528
rect 6606 8472 6611 8528
rect 5717 8470 6611 8472
rect 5717 8467 5783 8470
rect 6545 8467 6611 8470
rect 5533 8394 5599 8397
rect 6310 8394 6316 8396
rect 5533 8392 6316 8394
rect 5533 8336 5538 8392
rect 5594 8336 6316 8392
rect 5533 8334 6316 8336
rect 5533 8331 5599 8334
rect 6310 8332 6316 8334
rect 6380 8332 6386 8396
rect 17401 8394 17467 8397
rect 20897 8394 20963 8397
rect 17401 8392 20963 8394
rect 17401 8336 17406 8392
rect 17462 8336 20902 8392
rect 20958 8336 20963 8392
rect 17401 8334 20963 8336
rect 17401 8331 17467 8334
rect 20897 8331 20963 8334
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 5073 8122 5139 8125
rect 8201 8122 8267 8125
rect 5073 8120 8267 8122
rect 5073 8064 5078 8120
rect 5134 8064 8206 8120
rect 8262 8064 8267 8120
rect 5073 8062 8267 8064
rect 5073 8059 5139 8062
rect 8201 8059 8267 8062
rect 3417 7986 3483 7989
rect 4102 7986 4108 7988
rect 3417 7984 4108 7986
rect 3417 7928 3422 7984
rect 3478 7928 4108 7984
rect 3417 7926 4108 7928
rect 3417 7923 3483 7926
rect 4102 7924 4108 7926
rect 4172 7986 4178 7988
rect 5073 7986 5139 7989
rect 4172 7984 5139 7986
rect 4172 7928 5078 7984
rect 5134 7928 5139 7984
rect 4172 7926 5139 7928
rect 4172 7924 4178 7926
rect 5073 7923 5139 7926
rect 15101 7986 15167 7989
rect 18137 7986 18203 7989
rect 15101 7984 18203 7986
rect 15101 7928 15106 7984
rect 15162 7928 18142 7984
rect 18198 7928 18203 7984
rect 15101 7926 18203 7928
rect 15101 7923 15167 7926
rect 18137 7923 18203 7926
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 12433 7442 12499 7445
rect 13721 7442 13787 7445
rect 12433 7440 13787 7442
rect 12433 7384 12438 7440
rect 12494 7384 13726 7440
rect 13782 7384 13787 7440
rect 12433 7382 13787 7384
rect 12433 7379 12499 7382
rect 13721 7379 13787 7382
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 4981 6900 5047 6901
rect 4981 6898 5028 6900
rect 4936 6896 5028 6898
rect 4936 6840 4986 6896
rect 4936 6838 5028 6840
rect 4981 6836 5028 6838
rect 5092 6836 5098 6900
rect 4981 6835 5047 6836
rect 10225 6762 10291 6765
rect 17401 6762 17467 6765
rect 10225 6760 17467 6762
rect 10225 6704 10230 6760
rect 10286 6704 17406 6760
rect 17462 6704 17467 6760
rect 10225 6702 17467 6704
rect 10225 6699 10291 6702
rect 17401 6699 17467 6702
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 18822 3708 18828 3772
rect 18892 3770 18898 3772
rect 23105 3770 23171 3773
rect 18892 3768 23171 3770
rect 18892 3712 23110 3768
rect 23166 3712 23171 3768
rect 18892 3710 23171 3712
rect 18892 3708 18898 3710
rect 23105 3707 23171 3710
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 6132 26284 6196 26348
rect 19564 26344 19628 26348
rect 19564 26288 19578 26344
rect 19578 26288 19628 26344
rect 19564 26284 19628 26288
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 18828 25604 18892 25668
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 5028 25060 5092 25124
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 16988 24984 17052 24988
rect 16988 24928 17002 24984
rect 17002 24928 17052 24984
rect 16988 24924 17052 24928
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 5028 23020 5092 23084
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 12756 22128 12820 22132
rect 12756 22072 12770 22128
rect 12770 22072 12820 22128
rect 12756 22068 12820 22072
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 5028 20708 5092 20772
rect 14596 20708 14660 20772
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 13492 19348 13556 19412
rect 13676 19408 13740 19412
rect 13676 19352 13690 19408
rect 13690 19352 13740 19408
rect 13676 19348 13740 19352
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 14596 17716 14660 17780
rect 8524 17580 8588 17644
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 13492 16084 13556 16148
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 5028 15404 5092 15468
rect 7420 15404 7484 15468
rect 16988 15268 17052 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 19564 15132 19628 15196
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 12756 14316 12820 14380
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 13676 13908 13740 13972
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 6316 12684 6380 12748
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 4108 10916 4172 10980
rect 8524 11052 8588 11116
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 6316 9556 6380 9620
rect 7420 9420 7484 9484
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 6132 9012 6196 9076
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 6316 8332 6380 8396
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 4108 7924 4172 7988
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 5028 6896 5092 6900
rect 5028 6840 5042 6896
rect 5042 6840 5092 6896
rect 5028 6836 5092 6840
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 18828 3708 18892 3772
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 7890 27232 8210 27792
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 6131 26348 6197 26349
rect 6131 26284 6132 26348
rect 6196 26284 6197 26348
rect 6131 26283 6197 26284
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 5027 25124 5093 25125
rect 5027 25060 5028 25124
rect 5092 25060 5093 25124
rect 5027 25059 5093 25060
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 5030 23085 5090 25059
rect 5027 23084 5093 23085
rect 5027 23020 5028 23084
rect 5092 23020 5093 23084
rect 5027 23019 5093 23020
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 5030 20773 5090 23019
rect 5027 20772 5093 20773
rect 5027 20708 5028 20772
rect 5092 20708 5093 20772
rect 5027 20707 5093 20708
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 5030 15469 5090 20707
rect 5027 15468 5093 15469
rect 5027 15404 5028 15468
rect 5092 15404 5093 15468
rect 5027 15403 5093 15404
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4107 10980 4173 10981
rect 4107 10916 4108 10980
rect 4172 10916 4173 10980
rect 4107 10915 4173 10916
rect 4110 7989 4170 10915
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4107 7988 4173 7989
rect 4107 7924 4108 7988
rect 4172 7924 4173 7988
rect 4107 7923 4173 7924
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 5030 6901 5090 15403
rect 6134 9077 6194 26283
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 14836 27232 15156 27792
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 21782 27232 22102 27792
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 19563 26348 19629 26349
rect 19563 26284 19564 26348
rect 19628 26284 19629 26348
rect 19563 26283 19629 26284
rect 18827 25668 18893 25669
rect 18827 25604 18828 25668
rect 18892 25604 18893 25668
rect 18827 25603 18893 25604
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 16987 24988 17053 24989
rect 16987 24924 16988 24988
rect 17052 24924 17053 24988
rect 16987 24923 17053 24924
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 12755 22132 12821 22133
rect 12755 22068 12756 22132
rect 12820 22068 12821 22132
rect 12755 22067 12821 22068
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 8523 17644 8589 17645
rect 8523 17580 8524 17644
rect 8588 17580 8589 17644
rect 8523 17579 8589 17580
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7419 15468 7485 15469
rect 7419 15404 7420 15468
rect 7484 15404 7485 15468
rect 7419 15403 7485 15404
rect 6315 12748 6381 12749
rect 6315 12684 6316 12748
rect 6380 12684 6381 12748
rect 6315 12683 6381 12684
rect 6318 9621 6378 12683
rect 6315 9620 6381 9621
rect 6315 9556 6316 9620
rect 6380 9556 6381 9620
rect 6315 9555 6381 9556
rect 6131 9076 6197 9077
rect 6131 9012 6132 9076
rect 6196 9012 6197 9076
rect 6131 9011 6197 9012
rect 6318 8397 6378 9555
rect 7422 9485 7482 15403
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 8526 11117 8586 17579
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 12758 14381 12818 22067
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14595 20772 14661 20773
rect 14595 20708 14596 20772
rect 14660 20708 14661 20772
rect 14595 20707 14661 20708
rect 13491 19412 13557 19413
rect 13491 19348 13492 19412
rect 13556 19348 13557 19412
rect 13491 19347 13557 19348
rect 13675 19412 13741 19413
rect 13675 19348 13676 19412
rect 13740 19348 13741 19412
rect 13675 19347 13741 19348
rect 13494 16149 13554 19347
rect 13491 16148 13557 16149
rect 13491 16084 13492 16148
rect 13556 16084 13557 16148
rect 13491 16083 13557 16084
rect 12755 14380 12821 14381
rect 12755 14316 12756 14380
rect 12820 14316 12821 14380
rect 12755 14315 12821 14316
rect 13678 13973 13738 19347
rect 14598 17781 14658 20707
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14595 17780 14661 17781
rect 14595 17716 14596 17780
rect 14660 17716 14661 17780
rect 14595 17715 14661 17716
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 16990 15333 17050 24923
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 16987 15332 17053 15333
rect 16987 15268 16988 15332
rect 17052 15268 17053 15332
rect 16987 15267 17053 15268
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 13675 13972 13741 13973
rect 13675 13908 13676 13972
rect 13740 13908 13741 13972
rect 13675 13907 13741 13908
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 8523 11116 8589 11117
rect 8523 11052 8524 11116
rect 8588 11052 8589 11116
rect 8523 11051 8589 11052
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7419 9484 7485 9485
rect 7419 9420 7420 9484
rect 7484 9420 7485 9484
rect 7419 9419 7485 9420
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 6315 8396 6381 8397
rect 6315 8332 6316 8396
rect 6380 8332 6381 8396
rect 6315 8331 6381 8332
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 5027 6900 5093 6901
rect 5027 6836 5028 6900
rect 5092 6836 5093 6900
rect 5027 6835 5093 6836
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18830 3773 18890 25603
rect 19566 15197 19626 26283
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 19563 15196 19629 15197
rect 19563 15132 19564 15196
rect 19628 15132 19629 15196
rect 19563 15131 19629 15132
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 18827 3772 18893 3773
rect 18827 3708 18828 3772
rect 18892 3708 18893 3772
rect 18827 3707 18893 3708
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 27232 29048 27792
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__C
timestamp 1666464484
transform -1 0 26312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__D
timestamp 1666464484
transform 1 0 23368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1666464484
transform -1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A0
timestamp 1666464484
transform -1 0 8004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A0
timestamp 1666464484
transform -1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A0
timestamp 1666464484
transform -1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1666464484
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A
timestamp 1666464484
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1666464484
transform -1 0 15916 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__S
timestamp 1666464484
transform 1 0 18584 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1666464484
transform -1 0 17112 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1666464484
transform -1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B1
timestamp 1666464484
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 1666464484
transform -1 0 26404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A3
timestamp 1666464484
transform -1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1666464484
transform 1 0 25668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1666464484
transform -1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B
timestamp 1666464484
transform -1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1666464484
transform -1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B
timestamp 1666464484
transform 1 0 23552 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B
timestamp 1666464484
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1666464484
transform -1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1666464484
transform 1 0 24196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1666464484
transform -1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1666464484
transform -1 0 24748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B
timestamp 1666464484
transform -1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1666464484
transform 1 0 5704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A2
timestamp 1666464484
transform 1 0 5520 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1666464484
transform -1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B2
timestamp 1666464484
transform 1 0 21804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2
timestamp 1666464484
transform 1 0 4140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B2
timestamp 1666464484
transform 1 0 25208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1666464484
transform -1 0 27416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1666464484
transform 1 0 4600 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1666464484
transform 1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B1
timestamp 1666464484
transform 1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1666464484
transform 1 0 26128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1666464484
transform 1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1666464484
transform -1 0 10212 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1666464484
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1666464484
transform 1 0 26772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1666464484
transform -1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A2
timestamp 1666464484
transform 1 0 26312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A2
timestamp 1666464484
transform 1 0 24564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__C
timestamp 1666464484
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__C
timestamp 1666464484
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A0
timestamp 1666464484
transform 1 0 21252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A0
timestamp 1666464484
transform 1 0 26036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A0
timestamp 1666464484
transform 1 0 25484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1666464484
transform 1 0 22632 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 1666464484
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1666464484
transform -1 0 2760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1666464484
transform -1 0 2024 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B
timestamp 1666464484
transform -1 0 2208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1666464484
transform 1 0 5060 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1666464484
transform -1 0 4232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B
timestamp 1666464484
transform 1 0 3496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B
timestamp 1666464484
transform -1 0 22540 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1666464484
transform 1 0 14260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1666464484
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B
timestamp 1666464484
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1666464484
transform -1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1666464484
transform -1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A
timestamp 1666464484
transform 1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B
timestamp 1666464484
transform 1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B
timestamp 1666464484
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1666464484
transform 1 0 2944 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B
timestamp 1666464484
transform -1 0 2576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__C
timestamp 1666464484
transform -1 0 3128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B
timestamp 1666464484
transform -1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1666464484
transform -1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B
timestamp 1666464484
transform 1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1666464484
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1666464484
transform -1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B
timestamp 1666464484
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1666464484
transform -1 0 6072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B1
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1666464484
transform -1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1666464484
transform 1 0 22816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1666464484
transform -1 0 8556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 1666464484
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__B1
timestamp 1666464484
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1666464484
transform -1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B
timestamp 1666464484
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1666464484
transform 1 0 4508 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B1
timestamp 1666464484
transform -1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1666464484
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B1
timestamp 1666464484
transform 1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B1
timestamp 1666464484
transform 1 0 2208 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B1
timestamp 1666464484
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B1
timestamp 1666464484
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B1
timestamp 1666464484
transform 1 0 2208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1666464484
transform -1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1666464484
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1666464484
transform 1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A2
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B1
timestamp 1666464484
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1666464484
transform -1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B1
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1666464484
transform -1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1666464484
transform -1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A2
timestamp 1666464484
transform -1 0 4048 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B1
timestamp 1666464484
transform 1 0 1840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A2
timestamp 1666464484
transform 1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B1
timestamp 1666464484
transform -1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A2
timestamp 1666464484
transform 1 0 2392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B1
timestamp 1666464484
transform 1 0 2392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1666464484
transform -1 0 3496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1666464484
transform -1 0 4140 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1666464484
transform 1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1666464484
transform -1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A2
timestamp 1666464484
transform 1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B1
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1666464484
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1666464484
transform -1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B1
timestamp 1666464484
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B1
timestamp 1666464484
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B1
timestamp 1666464484
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B1
timestamp 1666464484
transform -1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B1
timestamp 1666464484
transform -1 0 25944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B1
timestamp 1666464484
transform 1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B1
timestamp 1666464484
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B1
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1666464484
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B
timestamp 1666464484
transform 1 0 21988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A_N
timestamp 1666464484
transform 1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A_N
timestamp 1666464484
transform 1 0 23828 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A_N
timestamp 1666464484
transform -1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1666464484
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B1
timestamp 1666464484
transform -1 0 5428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B1
timestamp 1666464484
transform -1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B1
timestamp 1666464484
transform -1 0 2760 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B1
timestamp 1666464484
transform 1 0 1840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B1
timestamp 1666464484
transform 1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__B1
timestamp 1666464484
transform -1 0 1840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1666464484
transform 1 0 7084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 1666464484
transform 1 0 4876 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B1
timestamp 1666464484
transform 1 0 6532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B1
timestamp 1666464484
transform 1 0 5428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1666464484
transform -1 0 24380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1666464484
transform 1 0 8740 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B1
timestamp 1666464484
transform -1 0 9936 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B1
timestamp 1666464484
transform -1 0 8004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__B1
timestamp 1666464484
transform -1 0 11040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B1
timestamp 1666464484
transform -1 0 13432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B1
timestamp 1666464484
transform 1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1666464484
transform 1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__B1
timestamp 1666464484
transform 1 0 17480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1666464484
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A2
timestamp 1666464484
transform 1 0 17296 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A2
timestamp 1666464484
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B1
timestamp 1666464484
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A2
timestamp 1666464484
transform 1 0 16836 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1666464484
transform 1 0 16836 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A2
timestamp 1666464484
transform -1 0 15640 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B1
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A2
timestamp 1666464484
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A2
timestamp 1666464484
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B1
timestamp 1666464484
transform -1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A2
timestamp 1666464484
transform -1 0 22172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__B1
timestamp 1666464484
transform -1 0 22632 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A2
timestamp 1666464484
transform 1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B1
timestamp 1666464484
transform -1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A2
timestamp 1666464484
transform 1 0 7636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A2
timestamp 1666464484
transform -1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1
timestamp 1666464484
transform -1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1666464484
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform -1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 7360 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 10488 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 15088 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 20884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 23368 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 25852 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 27784 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1666464484
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35
timestamp 1666464484
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46
timestamp 1666464484
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1666464484
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1666464484
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1666464484
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1666464484
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1666464484
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1666464484
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1666464484
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1666464484
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1666464484
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_215
timestamp 1666464484
transform 1 0 20884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1666464484
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1666464484
transform 1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1666464484
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_270
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1666464484
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1666464484
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1666464484
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1666464484
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1666464484
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1666464484
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1666464484
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1666464484
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1666464484
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1666464484
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1666464484
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1666464484
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_197
timestamp 1666464484
transform 1 0 19228 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1666464484
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1666464484
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_251
timestamp 1666464484
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1666464484
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_264
timestamp 1666464484
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1666464484
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1666464484
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_71
timestamp 1666464484
transform 1 0 7636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1666464484
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1666464484
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1666464484
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1666464484
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1666464484
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1666464484
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1666464484
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1666464484
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1666464484
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1666464484
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_258
timestamp 1666464484
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_270
timestamp 1666464484
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_282
timestamp 1666464484
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1666464484
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1666464484
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1666464484
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1666464484
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 1666464484
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1666464484
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1666464484
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_180
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1666464484
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1666464484
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1666464484
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_43
timestamp 1666464484
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_46
timestamp 1666464484
transform 1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1666464484
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1666464484
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_66
timestamp 1666464484
transform 1 0 7176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1666464484
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1666464484
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1666464484
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1666464484
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1666464484
transform 1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1666464484
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1666464484
transform 1 0 14536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1666464484
transform 1 0 15088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1666464484
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_203
timestamp 1666464484
transform 1 0 19780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1666464484
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_217
timestamp 1666464484
transform 1 0 21068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1666464484
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1666464484
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_18
timestamp 1666464484
transform 1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_24
timestamp 1666464484
transform 1 0 3312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1666464484
transform 1 0 4140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_46
timestamp 1666464484
transform 1 0 5336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1666464484
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1666464484
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_72
timestamp 1666464484
transform 1 0 7728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1666464484
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1666464484
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_136
timestamp 1666464484
transform 1 0 13616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1666464484
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1666464484
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_180
timestamp 1666464484
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1666464484
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1666464484
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1666464484
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_232
timestamp 1666464484
transform 1 0 22448 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_240
timestamp 1666464484
transform 1 0 23184 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_244
timestamp 1666464484
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_256
timestamp 1666464484
transform 1 0 24656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_268
timestamp 1666464484
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1666464484
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1666464484
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_20
timestamp 1666464484
transform 1 0 2944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1666464484
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_33
timestamp 1666464484
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1666464484
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1666464484
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_57
timestamp 1666464484
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_63
timestamp 1666464484
transform 1 0 6900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_69
timestamp 1666464484
transform 1 0 7452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1666464484
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1666464484
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_107
timestamp 1666464484
transform 1 0 10948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_113
timestamp 1666464484
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1666464484
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1666464484
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1666464484
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1666464484
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1666464484
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1666464484
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1666464484
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1666464484
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_229
timestamp 1666464484
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1666464484
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1666464484
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1666464484
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_14
timestamp 1666464484
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_22
timestamp 1666464484
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1666464484
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1666464484
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_37
timestamp 1666464484
transform 1 0 4508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_45
timestamp 1666464484
transform 1 0 5244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_48
timestamp 1666464484
transform 1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_66
timestamp 1666464484
transform 1 0 7176 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_72
timestamp 1666464484
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1666464484
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_84
timestamp 1666464484
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1666464484
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1666464484
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_120
timestamp 1666464484
transform 1 0 12144 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_128
timestamp 1666464484
transform 1 0 12880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_183
timestamp 1666464484
transform 1 0 17940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1666464484
transform 1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_203
timestamp 1666464484
transform 1 0 19780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp 1666464484
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1666464484
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1666464484
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1666464484
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1666464484
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_16
timestamp 1666464484
transform 1 0 2576 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1666464484
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_43
timestamp 1666464484
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1666464484
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1666464484
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1666464484
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1666464484
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1666464484
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_89
timestamp 1666464484
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1666464484
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1666464484
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1666464484
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1666464484
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1666464484
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1666464484
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1666464484
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1666464484
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1666464484
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1666464484
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_12
timestamp 1666464484
transform 1 0 2208 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1666464484
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1666464484
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1666464484
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_48
timestamp 1666464484
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1666464484
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_73
timestamp 1666464484
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_77
timestamp 1666464484
transform 1 0 8188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1666464484
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1666464484
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1666464484
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1666464484
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_191
timestamp 1666464484
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1666464484
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1666464484
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_231
timestamp 1666464484
transform 1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1666464484
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_244
timestamp 1666464484
transform 1 0 23552 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_256
timestamp 1666464484
transform 1 0 24656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_268
timestamp 1666464484
transform 1 0 25760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_11
timestamp 1666464484
transform 1 0 2116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1666464484
transform 1 0 2668 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1666464484
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_37
timestamp 1666464484
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1666464484
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1666464484
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1666464484
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1666464484
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1666464484
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1666464484
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1666464484
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1666464484
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_204
timestamp 1666464484
transform 1 0 19872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_213
timestamp 1666464484
transform 1 0 20700 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1666464484
transform 1 0 21528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_231
timestamp 1666464484
transform 1 0 22356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1666464484
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_244
timestamp 1666464484
transform 1 0 23552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_257
timestamp 1666464484
transform 1 0 24748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_269
timestamp 1666464484
transform 1 0 25852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_281
timestamp 1666464484
transform 1 0 26956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1666464484
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1666464484
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1666464484
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1666464484
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1666464484
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1666464484
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1666464484
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1666464484
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1666464484
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_82
timestamp 1666464484
transform 1 0 8648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1666464484
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1666464484
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1666464484
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1666464484
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1666464484
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1666464484
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1666464484
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1666464484
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_230
timestamp 1666464484
transform 1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_234
timestamp 1666464484
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1666464484
transform 1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_263
timestamp 1666464484
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1666464484
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1666464484
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1666464484
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1666464484
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1666464484
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_47
timestamp 1666464484
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1666464484
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1666464484
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1666464484
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_102
timestamp 1666464484
transform 1 0 10488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1666464484
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_132
timestamp 1666464484
transform 1 0 13248 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1666464484
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1666464484
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1666464484
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1666464484
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1666464484
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_231
timestamp 1666464484
transform 1 0 22356 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_239
timestamp 1666464484
transform 1 0 23092 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1666464484
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_262
timestamp 1666464484
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1666464484
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_281
timestamp 1666464484
transform 1 0 26956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1666464484
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 1666464484
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1666464484
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1666464484
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1666464484
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1666464484
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1666464484
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1666464484
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_153
timestamp 1666464484
transform 1 0 15180 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_159
timestamp 1666464484
transform 1 0 15732 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1666464484
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_183
timestamp 1666464484
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_196
timestamp 1666464484
transform 1 0 19136 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1666464484
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1666464484
transform 1 0 22632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_238
timestamp 1666464484
transform 1 0 23000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1666464484
transform 1 0 23828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_258
timestamp 1666464484
transform 1 0 24840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_267
timestamp 1666464484
transform 1 0 25668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1666464484
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1666464484
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1666464484
transform 1 0 4784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1666464484
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_72
timestamp 1666464484
transform 1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1666464484
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1666464484
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1666464484
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_178
timestamp 1666464484
transform 1 0 17480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1666464484
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1666464484
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1666464484
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_229
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_239
timestamp 1666464484
transform 1 0 23092 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1666464484
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_260
timestamp 1666464484
transform 1 0 25024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_268
timestamp 1666464484
transform 1 0 25760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_274
timestamp 1666464484
transform 1 0 26312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_280
timestamp 1666464484
transform 1 0 26864 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_286
timestamp 1666464484
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1666464484
transform 1 0 28520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1666464484
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1666464484
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp 1666464484
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_44
timestamp 1666464484
transform 1 0 5152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1666464484
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1666464484
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1666464484
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_128
timestamp 1666464484
transform 1 0 12880 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1666464484
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_191
timestamp 1666464484
transform 1 0 18676 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1666464484
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1666464484
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1666464484
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1666464484
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_236
timestamp 1666464484
transform 1 0 22816 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1666464484
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_253
timestamp 1666464484
transform 1 0 24380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1666464484
transform 1 0 25668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1666464484
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1666464484
transform 1 0 5796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1666464484
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1666464484
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_107
timestamp 1666464484
transform 1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1666464484
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1666464484
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1666464484
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1666464484
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1666464484
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1666464484
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1666464484
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1666464484
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_232
timestamp 1666464484
transform 1 0 22448 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_238
timestamp 1666464484
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_244
timestamp 1666464484
transform 1 0 23552 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1666464484
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_262
timestamp 1666464484
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1666464484
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1666464484
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_281
timestamp 1666464484
transform 1 0 26956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1666464484
transform 1 0 2208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_65
timestamp 1666464484
transform 1 0 7084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1666464484
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1666464484
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_154
timestamp 1666464484
transform 1 0 15272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1666464484
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1666464484
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1666464484
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1666464484
transform 1 0 20976 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1666464484
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1666464484
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_234
timestamp 1666464484
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_238
timestamp 1666464484
transform 1 0 23000 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_259
timestamp 1666464484
transform 1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_270
timestamp 1666464484
transform 1 0 25944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1666464484
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1666464484
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1666464484
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1666464484
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1666464484
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1666464484
transform 1 0 9660 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1666464484
transform 1 0 10212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1666464484
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_129
timestamp 1666464484
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_149
timestamp 1666464484
transform 1 0 14812 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1666464484
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1666464484
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1666464484
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_227
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1666464484
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_271
timestamp 1666464484
transform 1 0 26036 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_283
timestamp 1666464484
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_295
timestamp 1666464484
transform 1 0 28244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1666464484
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_36
timestamp 1666464484
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_44
timestamp 1666464484
transform 1 0 5152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1666464484
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1666464484
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1666464484
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1666464484
transform 1 0 15548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1666464484
transform 1 0 17296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1666464484
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1666464484
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_231
timestamp 1666464484
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1666464484
transform 1 0 23092 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_248
timestamp 1666464484
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_259
timestamp 1666464484
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_268
timestamp 1666464484
transform 1 0 25760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1666464484
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1666464484
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1666464484
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1666464484
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_75
timestamp 1666464484
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_95
timestamp 1666464484
transform 1 0 9844 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1666464484
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1666464484
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1666464484
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1666464484
transform 1 0 18032 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1666464484
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1666464484
transform 1 0 20424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1666464484
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_225
timestamp 1666464484
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1666464484
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1666464484
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1666464484
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_10
timestamp 1666464484
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1666464484
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1666464484
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_72
timestamp 1666464484
transform 1 0 7728 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1666464484
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1666464484
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1666464484
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1666464484
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1666464484
transform 1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_185
timestamp 1666464484
transform 1 0 18124 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_196
timestamp 1666464484
transform 1 0 19136 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1666464484
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_210
timestamp 1666464484
transform 1 0 20424 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1666464484
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1666464484
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1666464484
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1666464484
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1666464484
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1666464484
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1666464484
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1666464484
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1666464484
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1666464484
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1666464484
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_94
timestamp 1666464484
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1666464484
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1666464484
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1666464484
transform 1 0 14720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_185
timestamp 1666464484
transform 1 0 18124 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1666464484
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1666464484
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1666464484
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1666464484
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_227
timestamp 1666464484
transform 1 0 21988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_235
timestamp 1666464484
transform 1 0 22724 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1666464484
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1666464484
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1666464484
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1666464484
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_270
timestamp 1666464484
transform 1 0 25944 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_282
timestamp 1666464484
transform 1 0 27048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1666464484
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1666464484
transform 1 0 28520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1666464484
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1666464484
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_37
timestamp 1666464484
transform 1 0 4508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1666464484
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1666464484
transform 1 0 7176 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1666464484
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_101
timestamp 1666464484
transform 1 0 10396 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1666464484
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1666464484
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1666464484
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_151
timestamp 1666464484
transform 1 0 14996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_160
timestamp 1666464484
transform 1 0 15824 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1666464484
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1666464484
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1666464484
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1666464484
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1666464484
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_229
timestamp 1666464484
transform 1 0 22172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1666464484
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1666464484
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_257
timestamp 1666464484
transform 1 0 24748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_265
timestamp 1666464484
transform 1 0 25484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1666464484
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1666464484
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_286
timestamp 1666464484
transform 1 0 27416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1666464484
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1666464484
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_95
timestamp 1666464484
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1666464484
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_145
timestamp 1666464484
transform 1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1666464484
transform 1 0 15272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_178
timestamp 1666464484
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1666464484
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_205
timestamp 1666464484
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_212
timestamp 1666464484
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_224
timestamp 1666464484
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_234
timestamp 1666464484
transform 1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1666464484
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1666464484
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1666464484
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1666464484
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1666464484
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1666464484
transform 1 0 28336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_25
timestamp 1666464484
transform 1 0 3404 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1666464484
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_66
timestamp 1666464484
transform 1 0 7176 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_72
timestamp 1666464484
transform 1 0 7728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1666464484
transform 1 0 10028 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1666464484
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_122
timestamp 1666464484
transform 1 0 12328 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1666464484
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1666464484
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1666464484
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1666464484
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1666464484
transform 1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_194
timestamp 1666464484
transform 1 0 18952 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1666464484
transform 1 0 19504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_208
timestamp 1666464484
transform 1 0 20240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1666464484
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1666464484
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1666464484
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_253
timestamp 1666464484
transform 1 0 24380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_263
timestamp 1666464484
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_292
timestamp 1666464484
transform 1 0 27968 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1666464484
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1666464484
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_38
timestamp 1666464484
transform 1 0 4600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1666464484
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1666464484
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_105
timestamp 1666464484
transform 1 0 10764 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_127
timestamp 1666464484
transform 1 0 12788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_148
timestamp 1666464484
transform 1 0 14720 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1666464484
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1666464484
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1666464484
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1666464484
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1666464484
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_232
timestamp 1666464484
transform 1 0 22448 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_238
timestamp 1666464484
transform 1 0 23000 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_257
timestamp 1666464484
transform 1 0 24748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_273
timestamp 1666464484
transform 1 0 26220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1666464484
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1666464484
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_67
timestamp 1666464484
transform 1 0 7268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1666464484
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1666464484
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1666464484
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_199
timestamp 1666464484
transform 1 0 19412 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1666464484
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1666464484
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1666464484
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1666464484
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1666464484
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1666464484
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1666464484
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1666464484
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1666464484
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1666464484
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_38
timestamp 1666464484
transform 1 0 4600 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1666464484
transform 1 0 5152 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1666464484
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1666464484
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1666464484
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_100
timestamp 1666464484
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_124
timestamp 1666464484
transform 1 0 12512 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_130
timestamp 1666464484
transform 1 0 13064 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1666464484
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1666464484
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1666464484
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_180
timestamp 1666464484
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1666464484
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_213
timestamp 1666464484
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1666464484
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_238
timestamp 1666464484
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1666464484
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_258
timestamp 1666464484
transform 1 0 24840 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_266
timestamp 1666464484
transform 1 0 25576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_273
timestamp 1666464484
transform 1 0 26220 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_284
timestamp 1666464484
transform 1 0 27232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1666464484
transform 1 0 28336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_12
timestamp 1666464484
transform 1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_36
timestamp 1666464484
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_48
timestamp 1666464484
transform 1 0 5520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1666464484
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_77
timestamp 1666464484
transform 1 0 8188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1666464484
transform 1 0 9108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1666464484
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_123
timestamp 1666464484
transform 1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1666464484
transform 1 0 15548 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1666464484
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1666464484
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_207
timestamp 1666464484
transform 1 0 20148 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_213
timestamp 1666464484
transform 1 0 20700 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1666464484
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_234
timestamp 1666464484
transform 1 0 22632 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1666464484
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1666464484
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_290
timestamp 1666464484
transform 1 0 27784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1666464484
transform 1 0 28520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_35
timestamp 1666464484
transform 1 0 4324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1666464484
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1666464484
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1666464484
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_108
timestamp 1666464484
transform 1 0 11040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_114
timestamp 1666464484
transform 1 0 11592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_131
timestamp 1666464484
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1666464484
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1666464484
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1666464484
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1666464484
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1666464484
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_206
timestamp 1666464484
transform 1 0 20056 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1666464484
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_225
timestamp 1666464484
transform 1 0 21804 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_237
timestamp 1666464484
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_244
timestamp 1666464484
transform 1 0 23552 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1666464484
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1666464484
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_291
timestamp 1666464484
transform 1 0 27876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1666464484
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_26
timestamp 1666464484
transform 1 0 3496 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_32
timestamp 1666464484
transform 1 0 4048 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1666464484
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_76
timestamp 1666464484
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1666464484
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1666464484
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1666464484
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_127
timestamp 1666464484
transform 1 0 12788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_133
timestamp 1666464484
transform 1 0 13340 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1666464484
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1666464484
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_190
timestamp 1666464484
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1666464484
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1666464484
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1666464484
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_232
timestamp 1666464484
transform 1 0 22448 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1666464484
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1666464484
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1666464484
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1666464484
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1666464484
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_288
timestamp 1666464484
transform 1 0 27600 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_296
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1666464484
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_69
timestamp 1666464484
transform 1 0 7452 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1666464484
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_96
timestamp 1666464484
transform 1 0 9936 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_104
timestamp 1666464484
transform 1 0 10672 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1666464484
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1666464484
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1666464484
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1666464484
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1666464484
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1666464484
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_188
timestamp 1666464484
transform 1 0 18400 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1666464484
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1666464484
transform 1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_223
timestamp 1666464484
transform 1 0 21620 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1666464484
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_234
timestamp 1666464484
transform 1 0 22632 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1666464484
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1666464484
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_272
timestamp 1666464484
transform 1 0 26128 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_287
timestamp 1666464484
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1666464484
transform 1 0 28244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1666464484
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1666464484
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_48
timestamp 1666464484
transform 1 0 5520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1666464484
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_61
timestamp 1666464484
transform 1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1666464484
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_83
timestamp 1666464484
transform 1 0 8740 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1666464484
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1666464484
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_133
timestamp 1666464484
transform 1 0 13340 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1666464484
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_148
timestamp 1666464484
transform 1 0 14720 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1666464484
transform 1 0 15456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1666464484
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1666464484
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 1666464484
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_207
timestamp 1666464484
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_214
timestamp 1666464484
transform 1 0 20792 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1666464484
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 1666464484
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_257
timestamp 1666464484
transform 1 0 24748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_264
timestamp 1666464484
transform 1 0 25392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_272
timestamp 1666464484
transform 1 0 26128 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1666464484
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1666464484
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_72
timestamp 1666464484
transform 1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1666464484
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_93
timestamp 1666464484
transform 1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_129
timestamp 1666464484
transform 1 0 12972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_151
timestamp 1666464484
transform 1 0 14996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1666464484
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_178
timestamp 1666464484
transform 1 0 17480 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_186
timestamp 1666464484
transform 1 0 18216 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1666464484
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1666464484
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_213
timestamp 1666464484
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1666464484
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1666464484
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_268
timestamp 1666464484
transform 1 0 25760 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1666464484
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1666464484
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_298
timestamp 1666464484
transform 1 0 28520 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1666464484
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1666464484
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_24
timestamp 1666464484
transform 1 0 3312 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1666464484
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_63
timestamp 1666464484
transform 1 0 6900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1666464484
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_90
timestamp 1666464484
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1666464484
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_131
timestamp 1666464484
transform 1 0 13156 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_142
timestamp 1666464484
transform 1 0 14168 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1666464484
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1666464484
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1666464484
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1666464484
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1666464484
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1666464484
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_229
timestamp 1666464484
transform 1 0 22172 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_235
timestamp 1666464484
transform 1 0 22724 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_243
timestamp 1666464484
transform 1 0 23460 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_251
timestamp 1666464484
transform 1 0 24196 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_258
timestamp 1666464484
transform 1 0 24840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_269
timestamp 1666464484
transform 1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1666464484
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_286
timestamp 1666464484
transform 1 0 27416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1666464484
transform 1 0 28520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1666464484
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1666464484
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_48
timestamp 1666464484
transform 1 0 5520 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1666464484
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_74
timestamp 1666464484
transform 1 0 7912 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_94
timestamp 1666464484
transform 1 0 9752 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_100
timestamp 1666464484
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_130
timestamp 1666464484
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_134
timestamp 1666464484
transform 1 0 13432 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1666464484
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_147
timestamp 1666464484
transform 1 0 14628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_167
timestamp 1666464484
transform 1 0 16468 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1666464484
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1666464484
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1666464484
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1666464484
transform 1 0 22080 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_234
timestamp 1666464484
transform 1 0 22632 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_242
timestamp 1666464484
transform 1 0 23368 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1666464484
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1666464484
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1666464484
transform 1 0 25944 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_283
timestamp 1666464484
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1666464484
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_8
timestamp 1666464484
transform 1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_18
timestamp 1666464484
transform 1 0 2760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1666464484
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1666464484
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1666464484
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_75
timestamp 1666464484
transform 1 0 8004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1666464484
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_100
timestamp 1666464484
transform 1 0 10304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_121
timestamp 1666464484
transform 1 0 12236 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1666464484
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1666464484
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1666464484
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1666464484
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1666464484
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1666464484
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1666464484
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1666464484
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1666464484
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_232
timestamp 1666464484
transform 1 0 22448 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_239
timestamp 1666464484
transform 1 0 23092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1666464484
transform 1 0 23460 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_250
timestamp 1666464484
transform 1 0 24104 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1666464484
transform 1 0 24840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_266
timestamp 1666464484
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1666464484
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1666464484
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1666464484
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1666464484
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_72
timestamp 1666464484
transform 1 0 7728 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_93
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_99
timestamp 1666464484
transform 1 0 10212 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1666464484
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_113
timestamp 1666464484
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_124
timestamp 1666464484
transform 1 0 12512 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_130
timestamp 1666464484
transform 1 0 13064 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1666464484
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1666464484
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1666464484
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_178
timestamp 1666464484
transform 1 0 17480 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1666464484
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1666464484
transform 1 0 20056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_214
timestamp 1666464484
transform 1 0 20792 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_220
timestamp 1666464484
transform 1 0 21344 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_232
timestamp 1666464484
transform 1 0 22448 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1666464484
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_259
timestamp 1666464484
transform 1 0 24932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1666464484
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_276
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_288
timestamp 1666464484
transform 1 0 27600 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_296
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_12
timestamp 1666464484
transform 1 0 2208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_36
timestamp 1666464484
transform 1 0 4416 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_44
timestamp 1666464484
transform 1 0 5152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1666464484
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1666464484
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_92
timestamp 1666464484
transform 1 0 9568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1666464484
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_103
timestamp 1666464484
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1666464484
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_155
timestamp 1666464484
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1666464484
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_179
timestamp 1666464484
transform 1 0 17572 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1666464484
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1666464484
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1666464484
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_209
timestamp 1666464484
transform 1 0 20332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1666464484
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1666464484
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1666464484
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_259
timestamp 1666464484
transform 1 0 24932 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_263
timestamp 1666464484
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1666464484
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_8
timestamp 1666464484
transform 1 0 1840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_14
timestamp 1666464484
transform 1 0 2392 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1666464484
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_35
timestamp 1666464484
transform 1 0 4324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_45
timestamp 1666464484
transform 1 0 5244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_51
timestamp 1666464484
transform 1 0 5796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_61
timestamp 1666464484
transform 1 0 6716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1666464484
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_94
timestamp 1666464484
transform 1 0 9752 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1666464484
transform 1 0 10580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_110
timestamp 1666464484
transform 1 0 11224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_116
timestamp 1666464484
transform 1 0 11776 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1666464484
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_128
timestamp 1666464484
transform 1 0 12880 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_131
timestamp 1666464484
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1666464484
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1666464484
transform 1 0 14444 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_169
timestamp 1666464484
transform 1 0 16652 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_175
timestamp 1666464484
transform 1 0 17204 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_182
timestamp 1666464484
transform 1 0 17848 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1666464484
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_212
timestamp 1666464484
transform 1 0 20608 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1666464484
transform 1 0 22080 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1666464484
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_262
timestamp 1666464484
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_274
timestamp 1666464484
transform 1 0 26312 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_286
timestamp 1666464484
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1666464484
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1666464484
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_10
timestamp 1666464484
transform 1 0 2024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_16
timestamp 1666464484
transform 1 0 2576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_22
timestamp 1666464484
transform 1 0 3128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_28
timestamp 1666464484
transform 1 0 3680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1666464484
transform 1 0 4232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_40
timestamp 1666464484
transform 1 0 4784 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1666464484
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_63
timestamp 1666464484
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1666464484
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_84
timestamp 1666464484
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_91
timestamp 1666464484
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1666464484
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1666464484
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1666464484
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_143
timestamp 1666464484
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_146
timestamp 1666464484
transform 1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_173
timestamp 1666464484
transform 1 0 17020 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_184
timestamp 1666464484
transform 1 0 18032 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_190
timestamp 1666464484
transform 1 0 18584 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1666464484
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_202
timestamp 1666464484
transform 1 0 19688 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_214
timestamp 1666464484
transform 1 0 20792 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_218
timestamp 1666464484
transform 1 0 21160 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_235
timestamp 1666464484
transform 1 0 22724 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_246
timestamp 1666464484
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_258
timestamp 1666464484
transform 1 0 24840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1666464484
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1666464484
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1666464484
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1666464484
transform 1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_16
timestamp 1666464484
transform 1 0 2576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1666464484
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_33
timestamp 1666464484
transform 1 0 4140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_39
timestamp 1666464484
transform 1 0 4692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_45
timestamp 1666464484
transform 1 0 5244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_49
timestamp 1666464484
transform 1 0 5612 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_52
timestamp 1666464484
transform 1 0 5888 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_61
timestamp 1666464484
transform 1 0 6716 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_67
timestamp 1666464484
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_73
timestamp 1666464484
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1666464484
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_92
timestamp 1666464484
transform 1 0 9568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_98
timestamp 1666464484
transform 1 0 10120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_108
timestamp 1666464484
transform 1 0 11040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_114
timestamp 1666464484
transform 1 0 11592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_118
timestamp 1666464484
transform 1 0 11960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_129
timestamp 1666464484
transform 1 0 12972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1666464484
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_150
timestamp 1666464484
transform 1 0 14904 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_156
timestamp 1666464484
transform 1 0 15456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1666464484
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_163
timestamp 1666464484
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1666464484
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_171
timestamp 1666464484
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1666464484
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_182
timestamp 1666464484
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1666464484
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_10
timestamp 1666464484
transform 1 0 2024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_16
timestamp 1666464484
transform 1 0 2576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_26
timestamp 1666464484
transform 1 0 3496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_32
timestamp 1666464484
transform 1 0 4048 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_40
timestamp 1666464484
transform 1 0 4784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_43
timestamp 1666464484
transform 1 0 5060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1666464484
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_67
timestamp 1666464484
transform 1 0 7268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_73
timestamp 1666464484
transform 1 0 7820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_80
timestamp 1666464484
transform 1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_89
timestamp 1666464484
transform 1 0 9292 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1666464484
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1666464484
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1666464484
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1666464484
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1666464484
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1666464484
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1666464484
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1666464484
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_173
timestamp 1666464484
transform 1 0 17020 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_186
timestamp 1666464484
transform 1 0 18216 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_192
timestamp 1666464484
transform 1 0 18768 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_204
timestamp 1666464484
transform 1 0 19872 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1666464484
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1666464484
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_12
timestamp 1666464484
transform 1 0 2208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_18
timestamp 1666464484
transform 1 0 2760 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1666464484
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_33
timestamp 1666464484
transform 1 0 4140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_47
timestamp 1666464484
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_59
timestamp 1666464484
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_71
timestamp 1666464484
transform 1 0 7636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_75
timestamp 1666464484
transform 1 0 8004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1666464484
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1666464484
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1666464484
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1666464484
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1666464484
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_118
timestamp 1666464484
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_123
timestamp 1666464484
transform 1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1666464484
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1666464484
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_159
timestamp 1666464484
transform 1 0 15732 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_172
timestamp 1666464484
transform 1 0 16928 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1666464484
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1666464484
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_202
timestamp 1666464484
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_214
timestamp 1666464484
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_226
timestamp 1666464484
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_238
timestamp 1666464484
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1666464484
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_261
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1666464484
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1666464484
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_99
timestamp 1666464484
transform 1 0 10212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1666464484
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_123
timestamp 1666464484
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1666464484
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_142
timestamp 1666464484
transform 1 0 14168 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_154
timestamp 1666464484
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_158
timestamp 1666464484
transform 1 0 15640 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_174
timestamp 1666464484
transform 1 0 17112 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_186
timestamp 1666464484
transform 1 0 18216 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_198
timestamp 1666464484
transform 1 0 19320 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_210
timestamp 1666464484
transform 1 0 20424 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_23
timestamp 1666464484
transform 1 0 3220 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1666464484
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_35
timestamp 1666464484
transform 1 0 4324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_47
timestamp 1666464484
transform 1 0 5428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_55
timestamp 1666464484
transform 1 0 6164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_57
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1666464484
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_68
timestamp 1666464484
transform 1 0 7360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1666464484
transform 1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1666464484
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_102
timestamp 1666464484
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1666464484
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1666464484
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_118
timestamp 1666464484
transform 1 0 11960 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_124
timestamp 1666464484
transform 1 0 12512 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_128
timestamp 1666464484
transform 1 0 12880 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1666464484
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_152
timestamp 1666464484
transform 1 0 15088 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1666464484
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1666464484
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1666464484
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_180
timestamp 1666464484
transform 1 0 17664 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1666464484
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1666464484
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1666464484
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_212
timestamp 1666464484
transform 1 0 20608 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1666464484
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_222
timestamp 1666464484
transform 1 0 21528 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1666464484
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_237
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_242
timestamp 1666464484
transform 1 0 23368 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1666464484
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_269
timestamp 1666464484
transform 1 0 25852 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_276
timestamp 1666464484
transform 1 0 26496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_281
timestamp 1666464484
transform 1 0 26956 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1666464484
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1666464484
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1666464484
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0537_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20608 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0539_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20884 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _0541_
timestamp 1666464484
transform -1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0542_
timestamp 1666464484
transform -1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0543_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21528 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0544_
timestamp 1666464484
transform -1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0545_
timestamp 1666464484
transform -1 0 20240 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19872 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1666464484
transform 1 0 17848 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0554_
timestamp 1666464484
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1666464484
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17664 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0558_
timestamp 1666464484
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0559_
timestamp 1666464484
transform 1 0 19044 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1666464484
transform -1 0 16376 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1666464484
transform -1 0 18584 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1666464484
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1666464484
transform -1 0 17664 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0565_
timestamp 1666464484
transform -1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0567_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21160 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1666464484
transform 1 0 16836 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1666464484
transform -1 0 15548 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1666464484
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13616 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1666464484
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1666464484
transform -1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0576_
timestamp 1666464484
transform -1 0 13524 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0577_
timestamp 1666464484
transform 1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 1666464484
transform 1 0 12512 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1666464484
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0580_
timestamp 1666464484
transform -1 0 13616 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1666464484
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1666464484
transform 1 0 11776 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0583_
timestamp 1666464484
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0584_
timestamp 1666464484
transform -1 0 13432 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1666464484
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1666464484
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1666464484
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0589_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14720 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0591_
timestamp 1666464484
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0592_
timestamp 1666464484
transform 1 0 21896 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24012 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1666464484
transform -1 0 15732 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1666464484
transform -1 0 16468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1666464484
transform 1 0 17296 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1666464484
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1666464484
transform 1 0 17388 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1666464484
transform -1 0 17848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1666464484
transform 1 0 16100 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0601_
timestamp 1666464484
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1666464484
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0603_
timestamp 1666464484
transform -1 0 21528 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17940 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17388 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1666464484
transform -1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0607_
timestamp 1666464484
transform -1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1666464484
transform 1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7912 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0610_
timestamp 1666464484
transform -1 0 7820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1666464484
transform -1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1666464484
transform -1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1666464484
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1666464484
transform -1 0 8280 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _0615_
timestamp 1666464484
transform -1 0 9752 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1666464484
transform -1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0618_
timestamp 1666464484
transform -1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0619_
timestamp 1666464484
transform -1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0620_
timestamp 1666464484
transform -1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19872 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0622_
timestamp 1666464484
transform -1 0 25668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0623_
timestamp 1666464484
transform -1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0624_
timestamp 1666464484
transform 1 0 18308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0625_
timestamp 1666464484
transform -1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0626_
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0627_
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0628_
timestamp 1666464484
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1666464484
transform 1 0 21160 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19044 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1666464484
transform 1 0 19412 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0632_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0633_
timestamp 1666464484
transform 1 0 20056 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0634_
timestamp 1666464484
transform 1 0 18676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17296 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0636_
timestamp 1666464484
transform 1 0 18032 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1666464484
transform -1 0 18032 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1666464484
transform 1 0 20608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0639_
timestamp 1666464484
transform -1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0640_
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20240 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_2  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19136 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0646_
timestamp 1666464484
transform 1 0 20884 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0647_
timestamp 1666464484
transform 1 0 18400 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1666464484
transform -1 0 19044 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 1666464484
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1666464484
transform -1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0652_
timestamp 1666464484
transform 1 0 22816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0655_
timestamp 1666464484
transform -1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1666464484
transform -1 0 22448 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22080 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22724 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1666464484
transform 1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0660_
timestamp 1666464484
transform 1 0 21712 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_2  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23552 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0664_
timestamp 1666464484
transform -1 0 23184 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23092 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0667_
timestamp 1666464484
transform -1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0668_
timestamp 1666464484
transform 1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0669_
timestamp 1666464484
transform -1 0 24840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0670_
timestamp 1666464484
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1666464484
transform -1 0 21528 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0672_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23920 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0674_
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0675_
timestamp 1666464484
transform -1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0677_
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0678_
timestamp 1666464484
transform 1 0 22816 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1666464484
transform -1 0 25852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0680_
timestamp 1666464484
transform 1 0 25024 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1666464484
transform 1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0682_
timestamp 1666464484
transform -1 0 24104 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0683_
timestamp 1666464484
transform 1 0 23552 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0684_
timestamp 1666464484
transform -1 0 24104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0685_
timestamp 1666464484
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1666464484
transform 1 0 21712 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0687_
timestamp 1666464484
transform -1 0 23736 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0688_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0689_
timestamp 1666464484
transform 1 0 24288 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0690_
timestamp 1666464484
transform 1 0 25208 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 1666464484
transform 1 0 26312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0692_
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0694_
timestamp 1666464484
transform -1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1666464484
transform 1 0 24932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0696_
timestamp 1666464484
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23276 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24932 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26864 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1666464484
transform 1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1666464484
transform 1 0 25668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0702_
timestamp 1666464484
transform -1 0 23460 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0703_
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0704_
timestamp 1666464484
transform 1 0 25944 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1666464484
transform -1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26956 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0708_
timestamp 1666464484
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1666464484
transform -1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 1666464484
transform -1 0 27232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0711_
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0712_
timestamp 1666464484
transform -1 0 27508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25760 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0714_
timestamp 1666464484
transform -1 0 26680 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0715_
timestamp 1666464484
transform 1 0 26404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0716_
timestamp 1666464484
transform 1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1666464484
transform 1 0 25300 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23828 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0720_
timestamp 1666464484
transform 1 0 24472 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _0721_
timestamp 1666464484
transform -1 0 26220 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0722_
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0723_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0724_
timestamp 1666464484
transform 1 0 27876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0725_
timestamp 1666464484
transform -1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1666464484
transform -1 0 28060 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0727_
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _0728_
timestamp 1666464484
transform 1 0 26680 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0729_
timestamp 1666464484
transform -1 0 21436 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0730_
timestamp 1666464484
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0731_
timestamp 1666464484
transform 1 0 20240 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0732_
timestamp 1666464484
transform -1 0 20608 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1666464484
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0734_
timestamp 1666464484
transform 1 0 23460 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23368 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0736_
timestamp 1666464484
transform 1 0 22448 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0737_
timestamp 1666464484
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0738_
timestamp 1666464484
transform -1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0739_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0740_
timestamp 1666464484
transform 1 0 25668 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0741_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0742_
timestamp 1666464484
transform -1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0743_
timestamp 1666464484
transform 1 0 24748 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1666464484
transform 1 0 27876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1666464484
transform 1 0 28060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 1666464484
transform 1 0 27048 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0749_
timestamp 1666464484
transform 1 0 23276 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0750_
timestamp 1666464484
transform -1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 1666464484
transform -1 0 24196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0752_
timestamp 1666464484
transform 1 0 23092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22172 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0754_
timestamp 1666464484
transform -1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0755_
timestamp 1666464484
transform -1 0 23828 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1666464484
transform 1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14536 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0758_
timestamp 1666464484
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1666464484
transform 1 0 20976 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0760_
timestamp 1666464484
transform 1 0 11684 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0761_
timestamp 1666464484
transform -1 0 11224 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0762_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10672 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0763_
timestamp 1666464484
transform 1 0 11868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1666464484
transform -1 0 9568 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8924 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 1666464484
transform 1 0 9108 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0767_
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0768_
timestamp 1666464484
transform 1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1666464484
transform -1 0 8648 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0770_
timestamp 1666464484
transform 1 0 9384 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0771_
timestamp 1666464484
transform -1 0 8464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1666464484
transform 1 0 11684 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 1666464484
transform 1 0 11868 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0774_
timestamp 1666464484
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0775_
timestamp 1666464484
transform 1 0 8924 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1666464484
transform 1 0 10120 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0777_
timestamp 1666464484
transform -1 0 11224 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1666464484
transform 1 0 14260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 1666464484
transform 1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0780_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15272 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14168 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0782_
timestamp 1666464484
transform -1 0 12604 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0783_
timestamp 1666464484
transform 1 0 17664 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 1666464484
transform -1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0785_
timestamp 1666464484
transform -1 0 13616 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1666464484
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0787_
timestamp 1666464484
transform -1 0 12328 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0788_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0789_
timestamp 1666464484
transform -1 0 10488 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0790_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6164 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0791_
timestamp 1666464484
transform 1 0 9108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0792_
timestamp 1666464484
transform -1 0 20148 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0793_
timestamp 1666464484
transform -1 0 12972 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0794_
timestamp 1666464484
transform 1 0 20516 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0795_
timestamp 1666464484
transform -1 0 2024 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0796_
timestamp 1666464484
transform -1 0 5704 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0797_
timestamp 1666464484
transform 1 0 4784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1666464484
transform -1 0 16744 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0799_
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1666464484
transform -1 0 13800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1666464484
transform -1 0 20792 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1666464484
transform -1 0 9384 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0804_
timestamp 1666464484
transform 1 0 13156 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0805_
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0806_
timestamp 1666464484
transform 1 0 11684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0807_
timestamp 1666464484
transform -1 0 13340 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0808_
timestamp 1666464484
transform -1 0 13984 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0809_
timestamp 1666464484
transform 1 0 9292 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _0810_
timestamp 1666464484
transform -1 0 11040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0811_
timestamp 1666464484
transform -1 0 11224 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0812_
timestamp 1666464484
transform -1 0 10672 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1666464484
transform 1 0 11684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1666464484
transform 1 0 12328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1666464484
transform 1 0 12052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0816_
timestamp 1666464484
transform -1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1666464484
transform -1 0 11040 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0818_
timestamp 1666464484
transform 1 0 11040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0819_
timestamp 1666464484
transform 1 0 12328 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0820_
timestamp 1666464484
transform 1 0 8832 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0821_
timestamp 1666464484
transform -1 0 10212 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12512 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1666464484
transform 1 0 12604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0824_
timestamp 1666464484
transform 1 0 12788 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0825_
timestamp 1666464484
transform 1 0 13248 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0826_
timestamp 1666464484
transform -1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0827_
timestamp 1666464484
transform 1 0 14628 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0828_
timestamp 1666464484
transform -1 0 12512 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1666464484
transform 1 0 13156 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 1666464484
transform -1 0 13800 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _0831_
timestamp 1666464484
transform -1 0 13616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0832_
timestamp 1666464484
transform -1 0 13800 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0833_
timestamp 1666464484
transform -1 0 13432 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1666464484
transform -1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0836_
timestamp 1666464484
transform -1 0 14812 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0837_
timestamp 1666464484
transform 1 0 13984 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0838_
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0840_
timestamp 1666464484
transform 1 0 24564 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1666464484
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1666464484
transform 1 0 20608 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0843_
timestamp 1666464484
transform -1 0 22632 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0844_
timestamp 1666464484
transform 1 0 21528 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0845_
timestamp 1666464484
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0846_
timestamp 1666464484
transform -1 0 14260 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1666464484
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0848_
timestamp 1666464484
transform -1 0 9752 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0849_
timestamp 1666464484
transform 1 0 6624 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0850_
timestamp 1666464484
transform 1 0 9936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0851_
timestamp 1666464484
transform 1 0 17112 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1666464484
transform 1 0 3956 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0853_
timestamp 1666464484
transform 1 0 11868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0854_
timestamp 1666464484
transform 1 0 13432 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0855_
timestamp 1666464484
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0856_
timestamp 1666464484
transform -1 0 12328 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0857_
timestamp 1666464484
transform 1 0 12604 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0858_
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1666464484
transform 1 0 18216 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0860_
timestamp 1666464484
transform 1 0 23460 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0861_
timestamp 1666464484
transform -1 0 25024 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1666464484
transform -1 0 19688 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1666464484
transform 1 0 21068 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1666464484
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1666464484
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0866_
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0867_
timestamp 1666464484
transform 1 0 19596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0868_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0869_
timestamp 1666464484
transform 1 0 6532 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0870_
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1666464484
transform -1 0 10212 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0872_
timestamp 1666464484
transform 1 0 9108 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1666464484
transform 1 0 6532 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1666464484
transform -1 0 9936 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0876_
timestamp 1666464484
transform 1 0 10120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0877_
timestamp 1666464484
transform 1 0 14260 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0878_
timestamp 1666464484
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0879_
timestamp 1666464484
transform 1 0 12328 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0880_
timestamp 1666464484
transform -1 0 18952 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0881_
timestamp 1666464484
transform -1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1666464484
transform -1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0883_
timestamp 1666464484
transform 1 0 18124 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0884_
timestamp 1666464484
transform 1 0 23000 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1666464484
transform -1 0 25760 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0886_
timestamp 1666464484
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1666464484
transform -1 0 19964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0889_
timestamp 1666464484
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0891_
timestamp 1666464484
transform -1 0 14628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0892_
timestamp 1666464484
transform 1 0 19872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0893_
timestamp 1666464484
transform -1 0 8280 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0894_
timestamp 1666464484
transform -1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0895_
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0896_
timestamp 1666464484
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0897_
timestamp 1666464484
transform -1 0 8464 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0898_
timestamp 1666464484
transform 1 0 9108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0899_
timestamp 1666464484
transform 1 0 18676 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0900_
timestamp 1666464484
transform 1 0 18032 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1666464484
transform -1 0 25484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0903_
timestamp 1666464484
transform -1 0 18676 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1666464484
transform -1 0 20056 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0905_
timestamp 1666464484
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1666464484
transform -1 0 21804 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0907_
timestamp 1666464484
transform -1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0908_
timestamp 1666464484
transform 1 0 19780 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1666464484
transform 1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 1666464484
transform -1 0 21528 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1666464484
transform -1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1666464484
transform -1 0 21068 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0913_
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1666464484
transform -1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1666464484
transform 1 0 25576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0916_
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0917_
timestamp 1666464484
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0918_
timestamp 1666464484
transform -1 0 25300 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0919_
timestamp 1666464484
transform -1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _0920_
timestamp 1666464484
transform 1 0 19596 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1666464484
transform 1 0 23368 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0922_
timestamp 1666464484
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1666464484
transform -1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0924_
timestamp 1666464484
transform 1 0 18676 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1666464484
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0926_
timestamp 1666464484
transform 1 0 19412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0927_
timestamp 1666464484
transform 1 0 20516 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0928_
timestamp 1666464484
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 1666464484
transform -1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0930_
timestamp 1666464484
transform -1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1666464484
transform 1 0 25576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1666464484
transform -1 0 22540 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0933_
timestamp 1666464484
transform 1 0 24564 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0934_
timestamp 1666464484
transform -1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1666464484
transform -1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0936_
timestamp 1666464484
transform 1 0 23184 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0937_
timestamp 1666464484
transform -1 0 24932 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1666464484
transform 1 0 22724 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0939_
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0940_
timestamp 1666464484
transform 1 0 25300 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0941_
timestamp 1666464484
transform -1 0 24012 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0942_
timestamp 1666464484
transform -1 0 25300 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1666464484
transform -1 0 23000 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0944_
timestamp 1666464484
transform -1 0 23092 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0945_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23828 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0946_
timestamp 1666464484
transform 1 0 24196 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0947_
timestamp 1666464484
transform 1 0 23184 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1666464484
transform 1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1666464484
transform -1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1666464484
transform -1 0 18952 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1666464484
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0952_
timestamp 1666464484
transform 1 0 15180 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1666464484
transform -1 0 12604 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0954_
timestamp 1666464484
transform -1 0 7820 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1666464484
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0956_
timestamp 1666464484
transform -1 0 20332 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1666464484
transform 1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1666464484
transform 1 0 8372 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1666464484
transform -1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1666464484
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1666464484
transform -1 0 13800 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1666464484
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 1666464484
transform -1 0 17848 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0965_
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 1666464484
transform 1 0 18308 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0967_
timestamp 1666464484
transform 1 0 18032 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 1666464484
transform 1 0 17848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0969_
timestamp 1666464484
transform -1 0 15272 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1666464484
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1666464484
transform 1 0 16652 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0972_
timestamp 1666464484
transform -1 0 16376 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1666464484
transform 1 0 21252 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1666464484
transform -1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0975_
timestamp 1666464484
transform -1 0 22632 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0976_
timestamp 1666464484
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12236 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0978_
timestamp 1666464484
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1666464484
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0980_
timestamp 1666464484
transform 1 0 1656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1666464484
transform -1 0 7728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0982_
timestamp 1666464484
transform 1 0 4324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1666464484
transform -1 0 8740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0984_
timestamp 1666464484
transform -1 0 3680 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1666464484
transform -1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0986_
timestamp 1666464484
transform -1 0 14720 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0987_
timestamp 1666464484
transform -1 0 12972 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0988_
timestamp 1666464484
transform -1 0 14720 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0989_
timestamp 1666464484
transform 1 0 13064 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1666464484
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0991_
timestamp 1666464484
transform 1 0 14720 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0992_
timestamp 1666464484
transform -1 0 6072 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0993_
timestamp 1666464484
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0994_
timestamp 1666464484
transform -1 0 6072 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1666464484
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0996_
timestamp 1666464484
transform 1 0 1656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1666464484
transform -1 0 4324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0998_
timestamp 1666464484
transform -1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1666464484
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1000_
timestamp 1666464484
transform -1 0 2760 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1002_
timestamp 1666464484
transform -1 0 11040 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1003_
timestamp 1666464484
transform 1 0 7452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1004_
timestamp 1666464484
transform 1 0 10672 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1005_
timestamp 1666464484
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1006_
timestamp 1666464484
transform -1 0 16376 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1007_
timestamp 1666464484
transform -1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1666464484
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1009_
timestamp 1666464484
transform 1 0 15088 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1010_
timestamp 1666464484
transform 1 0 10212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1011_
timestamp 1666464484
transform 1 0 4600 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1013_
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1014_
timestamp 1666464484
transform 1 0 10764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1015_
timestamp 1666464484
transform 1 0 5520 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1016_
timestamp 1666464484
transform -1 0 17296 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1017_
timestamp 1666464484
transform 1 0 9108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1018_
timestamp 1666464484
transform 1 0 6624 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1666464484
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1020_
timestamp 1666464484
transform 1 0 15364 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1021_
timestamp 1666464484
transform -1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1022_
timestamp 1666464484
transform 1 0 8372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1023_
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1024_
timestamp 1666464484
transform 1 0 5520 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1025_
timestamp 1666464484
transform -1 0 2208 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1026_
timestamp 1666464484
transform 1 0 4232 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1027_
timestamp 1666464484
transform -1 0 2208 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1028_
timestamp 1666464484
transform -1 0 2208 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1029_
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1030_
timestamp 1666464484
transform 1 0 2944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1031_
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1032_
timestamp 1666464484
transform -1 0 3496 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1033_
timestamp 1666464484
transform 1 0 3956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1666464484
transform 1 0 3128 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1035_
timestamp 1666464484
transform 1 0 2760 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1036_
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1037_
timestamp 1666464484
transform 1 0 2944 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1038_
timestamp 1666464484
transform -1 0 12236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1039_
timestamp 1666464484
transform -1 0 7084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1040_
timestamp 1666464484
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1041_
timestamp 1666464484
transform 1 0 10028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1042_
timestamp 1666464484
transform 1 0 8096 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1043_
timestamp 1666464484
transform -1 0 9660 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1044_
timestamp 1666464484
transform 1 0 10028 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1666464484
transform 1 0 12604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1046_
timestamp 1666464484
transform 1 0 12788 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1047_
timestamp 1666464484
transform 1 0 20424 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1048_
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1049_
timestamp 1666464484
transform -1 0 14812 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1050_
timestamp 1666464484
transform -1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1051_
timestamp 1666464484
transform 1 0 17664 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1052_
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1053_
timestamp 1666464484
transform 1 0 17664 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1054_
timestamp 1666464484
transform -1 0 17296 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1055_
timestamp 1666464484
transform -1 0 12972 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1056_
timestamp 1666464484
transform 1 0 20240 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1057_
timestamp 1666464484
transform -1 0 19504 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1058_
timestamp 1666464484
transform -1 0 18308 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1059_
timestamp 1666464484
transform -1 0 19872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1060_
timestamp 1666464484
transform -1 0 12144 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1061_
timestamp 1666464484
transform -1 0 9384 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1062_
timestamp 1666464484
transform 1 0 10672 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1063_
timestamp 1666464484
transform -1 0 12144 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1064_
timestamp 1666464484
transform 1 0 18216 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1065_
timestamp 1666464484
transform 1 0 14812 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1066__1
timestamp 1666464484
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067__2
timestamp 1666464484
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068__3
timestamp 1666464484
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069__4
timestamp 1666464484
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070__5
timestamp 1666464484
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071__6
timestamp 1666464484
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072__7
timestamp 1666464484
transform -1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073__8
timestamp 1666464484
transform -1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1074_
timestamp 1666464484
transform -1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1075_
timestamp 1666464484
transform 1 0 9752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1076_
timestamp 1666464484
transform -1 0 14812 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1077_
timestamp 1666464484
transform 1 0 11868 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1666464484
transform 1 0 21988 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1666464484
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1080_
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1666464484
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1082_
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 1666464484
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1084_
timestamp 1666464484
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1086_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1087_
timestamp 1666464484
transform 1 0 4692 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1088_
timestamp 1666464484
transform -1 0 3496 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 1666464484
transform 1 0 2024 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1090_
timestamp 1666464484
transform 1 0 2208 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1091_
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1092_
timestamp 1666464484
transform -1 0 4692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1093_
timestamp 1666464484
transform 1 0 6992 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1094_
timestamp 1666464484
transform -1 0 4876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1095_
timestamp 1666464484
transform -1 0 6716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1096_
timestamp 1666464484
transform -1 0 6072 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1097_
timestamp 1666464484
transform -1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1098_
timestamp 1666464484
transform 1 0 9016 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1099_
timestamp 1666464484
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1100_
timestamp 1666464484
transform -1 0 8648 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1101_
timestamp 1666464484
transform 1 0 8096 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1666464484
transform 1 0 10304 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1103_
timestamp 1666464484
transform -1 0 12236 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1104_
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1105_
timestamp 1666464484
transform -1 0 16192 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1106_
timestamp 1666464484
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1107_
timestamp 1666464484
transform -1 0 16192 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1108_
timestamp 1666464484
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1109_
timestamp 1666464484
transform 1 0 15548 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1110_
timestamp 1666464484
transform -1 0 14536 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1111_
timestamp 1666464484
transform 1 0 17020 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1112_
timestamp 1666464484
transform 1 0 15732 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1113_
timestamp 1666464484
transform 1 0 17848 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1114_
timestamp 1666464484
transform -1 0 16100 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1115_
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1116_
timestamp 1666464484
transform 1 0 18032 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1117_
timestamp 1666464484
transform 1 0 7452 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1118_
timestamp 1666464484
transform -1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4232 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1666464484
transform 1 0 4692 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1666464484
transform 1 0 6072 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1666464484
transform 1 0 6532 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1666464484
transform 1 0 4324 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1666464484
transform 1 0 4600 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1666464484
transform 1 0 2392 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1666464484
transform 1 0 2024 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1666464484
transform 1 0 2024 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1666464484
transform 1 0 2024 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1666464484
transform 1 0 2576 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1666464484
transform -1 0 3496 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1666464484
transform 1 0 4416 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1666464484
transform 1 0 2024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1666464484
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1666464484
transform 1 0 2116 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1666464484
transform 1 0 2024 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1666464484
transform 1 0 2024 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1666464484
transform -1 0 9016 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1666464484
transform 1 0 9476 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1666464484
transform -1 0 8648 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1666464484
transform -1 0 8924 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1666464484
transform 1 0 9292 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1666464484
transform 1 0 11684 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1666464484
transform 1 0 11684 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _1145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13156 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21528 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 1666464484
transform 1 0 15916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1149_
timestamp 1666464484
transform 1 0 15916 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1666464484
transform 1 0 14260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1666464484
transform 1 0 9292 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1666464484
transform 1 0 9752 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1666464484
transform 1 0 9660 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1666464484
transform 1 0 18032 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1666464484
transform 1 0 17480 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1666464484
transform 1 0 14260 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1666464484
transform 1 0 14168 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1666464484
transform 1 0 9384 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1666464484
transform 1 0 9476 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1666464484
transform 1 0 11500 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1666464484
transform 1 0 9752 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1666464484
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1666464484
transform 1 0 16836 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1666464484
transform 1 0 14260 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1666464484
transform 1 0 13984 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1666464484
transform 1 0 9384 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1666464484
transform 1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1666464484
transform 1 0 11684 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1666464484
transform 1 0 11040 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23368 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1174_
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1666464484
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1666464484
transform -1 0 21528 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _1177_
timestamp 1666464484
transform 1 0 22724 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1178_
timestamp 1666464484
transform 1 0 14352 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1666464484
transform 1 0 9752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1666464484
transform 1 0 10488 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1666464484
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1666464484
transform 1 0 12420 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1666464484
transform 1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1666464484
transform 1 0 15916 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1666464484
transform -1 0 19228 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1666464484
transform -1 0 19872 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1666464484
transform 1 0 9476 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1666464484
transform 1 0 9568 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1666464484
transform -1 0 12788 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1666464484
transform 1 0 11684 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1666464484
transform -1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1666464484
transform -1 0 22908 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1666464484
transform 1 0 21988 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1666464484
transform 1 0 4048 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1666464484
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1666464484
transform 1 0 6716 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp 1666464484
transform 1 0 4600 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp 1666464484
transform 1 0 6624 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1666464484
transform 1 0 4692 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1666464484
transform 1 0 6532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp 1666464484
transform 1 0 6440 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1666464484
transform 1 0 6992 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1666464484
transform -1 0 10580 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp 1666464484
transform 1 0 7912 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp 1666464484
transform 1 0 9752 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp 1666464484
transform 1 0 11684 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp 1666464484
transform 1 0 17112 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp 1666464484
transform 1 0 16836 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1666464484
transform 1 0 15272 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1666464484
transform 1 0 16836 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1666464484
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 1666464484
transform 1 0 14996 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1666464484
transform 1 0 14904 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp 1666464484
transform 1 0 16836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1220_
timestamp 1666464484
transform 1 0 15916 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1221_
timestamp 1666464484
transform 1 0 17020 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp 1666464484
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp 1666464484
transform 1 0 6532 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1224_
timestamp 1666464484
transform 1 0 4600 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10304 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform -1 0 5888 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform -1 0 8372 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 6808 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform -1 0 12236 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 15272 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 15088 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 6072 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 6164 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform -1 0 4140 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 1656 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 10580 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform -1 0 12512 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0142_
timestamp 1666464484
transform 1 0 13248 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0143_
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0498_
timestamp 1666464484
transform 1 0 7820 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0502_
timestamp 1666464484
transform 1 0 14444 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0526_
timestamp 1666464484
transform 1 0 16836 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 13340 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 11224 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform -1 0 4416 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 5244 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform -1 0 7084 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform -1 0 17480 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform -1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform -1 0 3404 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform -1 0 3404 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 1564 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform -1 0 9660 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform -1 0 9660 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0142_
timestamp 1666464484
transform -1 0 14812 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0143_
timestamp 1666464484
transform -1 0 14812 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0498_
timestamp 1666464484
transform -1 0 7084 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0502_
timestamp 1666464484
transform -1 0 12236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0526_
timestamp 1666464484
transform -1 0 17480 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1666464484
transform -1 0 11592 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 9660 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform -1 0 4416 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 5244 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 5244 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 12972 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 12972 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform -1 0 6072 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform -1 0 4416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform -1 0 3404 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 1564 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 12972 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0142_
timestamp 1666464484
transform -1 0 13800 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0143_
timestamp 1666464484
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0498_
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0502_
timestamp 1666464484
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0526_
timestamp 1666464484
transform -1 0 17480 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1666464484
transform 1 0 12972 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 9384 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 14536 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 16836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform 1 0 21252 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform 1 0 23736 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform 1 0 26220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform 1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1666464484
transform 1 0 3956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform -1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1666464484
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1666464484
transform -1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1666464484
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1666464484
transform -1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_29
timestamp 1666464484
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_30
timestamp 1666464484
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_31
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_32
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_33
timestamp 1666464484
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_34
timestamp 1666464484
transform -1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_35
timestamp 1666464484
transform -1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_36
timestamp 1666464484
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_37
timestamp 1666464484
transform -1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_38
timestamp 1666464484
transform -1 0 28428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_39
timestamp 1666464484
transform -1 0 28428 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 1306 29200 1362 30000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 6274 29200 6330 30000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 8758 29200 8814 30000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 11242 29200 11298 30000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 13726 29200 13782 30000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 16210 29200 16266 30000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 18694 29200 18750 30000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 21178 29200 21234 30000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 23662 29200 23718 30000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 26146 29200 26202 30000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 28630 29200 28686 30000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 29200 14832 30000 14952 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 3790 29200 3846 30000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 7890 2128 8210 27792 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 27792 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 27792 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 27792 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel via1 15076 27200 15076 27200 0 vssd1
rlabel metal1 16376 14314 16376 14314 0 CIRCUIT_1957.D0
rlabel metal1 16415 13498 16415 13498 0 CIRCUIT_1957.D1
rlabel metal2 18630 14484 18630 14484 0 CIRCUIT_1957.D2
rlabel metal2 15732 24276 15732 24276 0 CIRCUIT_1957.D3
rlabel metal1 22126 9452 22126 9452 0 CIRCUIT_1957.GATES_10.result
rlabel metal1 14812 7310 14812 7310 0 CIRCUIT_1957.GATES_27.result
rlabel metal1 14053 11322 14053 11322 0 CIRCUIT_1957.GATES_28.result
rlabel metal1 16964 4590 16964 4590 0 CIRCUIT_1957.GATES_30.result
rlabel metal2 6670 8704 6670 8704 0 CIRCUIT_1957.GATES_33.input2
rlabel metal1 9977 4522 9977 4522 0 CIRCUIT_1957.GATES_35.result
rlabel metal2 11086 10064 11086 10064 0 CIRCUIT_1957.GATES_38.result
rlabel metal1 9706 7310 9706 7310 0 CIRCUIT_1957.GATES_39.result
rlabel metal2 14214 4624 14214 4624 0 CIRCUIT_1957.GATES_40.result
rlabel metal1 16882 7242 16882 7242 0 CIRCUIT_1957.GATES_41.result
rlabel metal1 9108 6766 9108 6766 0 CIRCUIT_1957.GATES_42.result
rlabel metal2 13570 7922 13570 7922 0 CIRCUIT_1957.GATES_53.result
rlabel metal1 15180 8534 15180 8534 0 CIRCUIT_1957.GATES_60.result
rlabel metal1 22218 12784 22218 12784 0 CIRCUIT_1957.GATES_9.result
rlabel metal1 16100 8602 16100 8602 0 CIRCUIT_1957.MEMORY_62.d
rlabel metal1 17572 9690 17572 9690 0 CIRCUIT_1957.MEMORY_62.s_currentState
rlabel metal1 23133 8534 23133 8534 0 CIRCUIT_1957.MEMORY_63.d
rlabel metal1 13386 5066 13386 5066 0 CIRCUIT_1957.MEMORY_63.s_currentState
rlabel metal2 22678 9928 22678 9928 0 CIRCUIT_1957.MEMORY_64.d
rlabel metal2 21114 10064 21114 10064 0 CIRCUIT_1957.MEMORY_64.s_currentState
rlabel metal1 20934 12818 20934 12818 0 CIRCUIT_1957.MEMORY_65.d
rlabel metal1 20378 12954 20378 12954 0 CIRCUIT_1957.MEMORY_65.s_currentState
rlabel metal2 23230 13090 23230 13090 0 CIRCUIT_1957.MEMORY_66.d
rlabel metal1 15088 13362 15088 13362 0 CIRCUIT_1957.MEMORY_66.s_currentState
rlabel metal1 24467 11798 24467 11798 0 CIRCUIT_1957.MEMORY_67.d
rlabel metal1 18952 9690 18952 9690 0 CIRCUIT_1957.MEMORY_67.s_currentState
rlabel metal1 13110 15436 13110 15436 0 CIRCUIT_1957.MEMORY_68.s_currentState
rlabel metal1 14536 13226 14536 13226 0 CIRCUIT_1957.MEMORY_69.s_currentState
rlabel metal1 15778 15470 15778 15470 0 CIRCUIT_1957.MEMORY_70.s_currentState
rlabel viali 15133 15470 15133 15470 0 CIRCUIT_1957.MEMORY_71.s_currentState
rlabel metal1 16836 6222 16836 6222 0 CIRCUIT_1957.MEMORY_72.s_currentState
rlabel metal1 16560 6290 16560 6290 0 CIRCUIT_1957.MEMORY_73.s_currentState
rlabel metal1 18630 6290 18630 6290 0 CIRCUIT_1957.MEMORY_74.s_currentState
rlabel metal2 18906 6154 18906 6154 0 CIRCUIT_1957.MEMORY_75.s_currentState
rlabel metal2 12650 7718 12650 7718 0 CIRCUIT_1957.MEMORY_76.s_currentState
rlabel metal1 12788 6970 12788 6970 0 CIRCUIT_1957.MEMORY_77.s_currentState
rlabel metal1 10902 5780 10902 5780 0 CIRCUIT_1957.MEMORY_78.s_currentState
rlabel metal2 12650 4964 12650 4964 0 CIRCUIT_1957.MEMORY_79.s_currentState
rlabel metal1 16376 5338 16376 5338 0 CIRCUIT_1957.MEMORY_80.s_currentState
rlabel metal2 15686 4828 15686 4828 0 CIRCUIT_1957.MEMORY_81.s_currentState
rlabel metal1 19228 4726 19228 4726 0 CIRCUIT_1957.MEMORY_82.s_currentState
rlabel metal1 19688 5338 19688 5338 0 CIRCUIT_1957.MEMORY_83.s_currentState
rlabel metal1 11500 6970 11500 6970 0 CIRCUIT_1957.MEMORY_84.s_currentState
rlabel metal2 12466 6868 12466 6868 0 CIRCUIT_1957.MEMORY_85.s_currentState
rlabel via1 12466 5661 12466 5661 0 CIRCUIT_1957.MEMORY_86.s_currentState
rlabel via1 12466 5117 12466 5117 0 CIRCUIT_1957.MEMORY_87.s_currentState
rlabel metal1 15456 8466 15456 8466 0 CIRCUIT_1957.MEMORY_88.s_currentState
rlabel metal1 15870 13294 15870 13294 0 CIRCUIT_1957.clock_gen_2_1.CLK1
rlabel metal1 21298 7310 21298 7310 0 CIRCUIT_1957.clock_gen_2_1.GATES_1.input2
rlabel metal1 19872 6766 19872 6766 0 CIRCUIT_1957.clock_gen_2_1.GATES_3.result
rlabel metal2 20470 6324 20470 6324 0 CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
rlabel metal1 17112 4046 17112 4046 0 CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState
rlabel metal1 13478 11832 13478 11832 0 CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d
rlabel metal1 16238 6766 16238 6766 0 CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState
rlabel metal1 16790 6766 16790 6766 0 CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState
rlabel metal2 7406 7752 7406 7752 0 CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1
rlabel metal1 6992 8466 6992 8466 0 CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2
rlabel metal2 7590 7242 7590 7242 0 CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result
rlabel metal1 18446 13294 18446 13294 0 CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState
rlabel metal1 19872 13294 19872 13294 0 CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState
rlabel metal1 20838 9010 20838 9010 0 CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState
rlabel metal1 17848 9554 17848 9554 0 CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState
rlabel metal2 5474 21318 5474 21318 0 CIRCUIT_1957.int_memory_1.GATES_1.input2\[0\]
rlabel metal1 5658 20230 5658 20230 0 CIRCUIT_1957.int_memory_1.GATES_1.input2\[1\]
rlabel metal1 5612 22406 5612 22406 0 CIRCUIT_1957.int_memory_1.GATES_1.input2\[2\]
rlabel metal1 2622 22576 2622 22576 0 CIRCUIT_1957.int_memory_1.GATES_1.input2\[3\]
rlabel metal1 7912 18394 7912 18394 0 CIRCUIT_1957.int_memory_1.GATES_2.input2\[0\]
rlabel metal2 6026 18258 6026 18258 0 CIRCUIT_1957.int_memory_1.GATES_2.input2\[1\]
rlabel metal1 8418 20536 8418 20536 0 CIRCUIT_1957.int_memory_1.GATES_2.input2\[2\]
rlabel metal1 5750 18938 5750 18938 0 CIRCUIT_1957.int_memory_1.GATES_2.input2\[3\]
rlabel metal2 8510 9826 8510 9826 0 CIRCUIT_1957.int_memory_1.GATES_21.result
rlabel metal1 7314 21114 7314 21114 0 CIRCUIT_1957.int_memory_1.GATES_22.result
rlabel metal1 8418 18734 8418 18734 0 CIRCUIT_1957.int_memory_1.GATES_23.result
rlabel metal2 7498 23494 7498 23494 0 CIRCUIT_1957.int_memory_1.GATES_24.result
rlabel metal2 12558 20910 12558 20910 0 CIRCUIT_1957.int_memory_1.GATES_25.result
rlabel metal1 14950 16422 14950 16422 0 CIRCUIT_1957.int_memory_1.GATES_26.result
rlabel metal1 14168 22202 14168 22202 0 CIRCUIT_1957.int_memory_1.GATES_27.result
rlabel metal1 16790 20502 16790 20502 0 CIRCUIT_1957.int_memory_1.GATES_28.result
rlabel metal1 5750 14382 5750 14382 0 CIRCUIT_1957.int_memory_1.GATES_29.result
rlabel metal1 6854 16048 6854 16048 0 CIRCUIT_1957.int_memory_1.GATES_3.input2\[0\]
rlabel metal1 5750 15130 5750 15130 0 CIRCUIT_1957.int_memory_1.GATES_3.input2\[1\]
rlabel metal1 7682 14518 7682 14518 0 CIRCUIT_1957.int_memory_1.GATES_3.input2\[2\]
rlabel metal1 7820 13158 7820 13158 0 CIRCUIT_1957.int_memory_1.GATES_3.input2\[3\]
rlabel metal1 6118 7514 6118 7514 0 CIRCUIT_1957.int_memory_1.GATES_30.result
rlabel metal2 4094 16830 4094 16830 0 CIRCUIT_1957.int_memory_1.GATES_31.result
rlabel metal2 4002 10608 4002 10608 0 CIRCUIT_1957.int_memory_1.GATES_32.result
rlabel metal1 1656 18734 1656 18734 0 CIRCUIT_1957.int_memory_1.GATES_33.result
rlabel via1 7313 12818 7313 12818 0 CIRCUIT_1957.int_memory_1.GATES_4.input2\[0\]
rlabel metal2 9522 13911 9522 13911 0 CIRCUIT_1957.int_memory_1.GATES_4.input2\[1\]
rlabel metal1 5750 8874 5750 8874 0 CIRCUIT_1957.int_memory_1.GATES_4.input2\[2\]
rlabel metal1 7774 13226 7774 13226 0 CIRCUIT_1957.int_memory_1.GATES_4.input2\[3\]
rlabel metal2 9246 13821 9246 13821 0 CIRCUIT_1957.int_memory_1.GATES_49.input2\[0\]
rlabel metal2 10718 15980 10718 15980 0 CIRCUIT_1957.int_memory_1.GATES_49.input2\[1\]
rlabel via1 12650 15130 12650 15130 0 CIRCUIT_1957.int_memory_1.GATES_49.input2\[2\]
rlabel metal1 13156 14382 13156 14382 0 CIRCUIT_1957.int_memory_1.GATES_49.input2\[3\]
rlabel metal2 3818 14926 3818 14926 0 CIRCUIT_1957.int_memory_1.GATES_5.input2\[0\]
rlabel metal1 4048 16558 4048 16558 0 CIRCUIT_1957.int_memory_1.GATES_5.input2\[1\]
rlabel metal1 3726 13498 3726 13498 0 CIRCUIT_1957.int_memory_1.GATES_5.input2\[2\]
rlabel metal1 1794 18224 1794 18224 0 CIRCUIT_1957.int_memory_1.GATES_5.input2\[3\]
rlabel metal1 10120 14314 10120 14314 0 CIRCUIT_1957.int_memory_1.GATES_50.result
rlabel metal1 9798 18394 9798 18394 0 CIRCUIT_1957.int_memory_1.GATES_51.input2\[0\]
rlabel metal1 10258 17578 10258 17578 0 CIRCUIT_1957.int_memory_1.GATES_51.input2\[1\]
rlabel metal1 12696 16762 12696 16762 0 CIRCUIT_1957.int_memory_1.GATES_51.input2\[2\]
rlabel metal1 13294 18598 13294 18598 0 CIRCUIT_1957.int_memory_1.GATES_51.input2\[3\]
rlabel metal2 11914 18394 11914 18394 0 CIRCUIT_1957.int_memory_1.GATES_53.result
rlabel metal1 3450 8806 3450 8806 0 CIRCUIT_1957.int_memory_1.GATES_6.input2\[0\]
rlabel metal1 3266 8840 3266 8840 0 CIRCUIT_1957.int_memory_1.GATES_6.input2\[1\]
rlabel metal1 4462 13702 4462 13702 0 CIRCUIT_1957.int_memory_1.GATES_6.input2\[2\]
rlabel metal1 3772 9418 3772 9418 0 CIRCUIT_1957.int_memory_1.GATES_6.input2\[3\]
rlabel metal1 3450 19924 3450 19924 0 CIRCUIT_1957.int_memory_1.GATES_7.input2\[0\]
rlabel metal2 3542 19312 3542 19312 0 CIRCUIT_1957.int_memory_1.GATES_7.input2\[1\]
rlabel metal2 3450 19754 3450 19754 0 CIRCUIT_1957.int_memory_1.GATES_7.input2\[2\]
rlabel metal1 3358 19482 3358 19482 0 CIRCUIT_1957.int_memory_1.GATES_7.input2\[3\]
rlabel metal1 7498 10778 7498 10778 0 CIRCUIT_1957.int_memory_1.GATES_8.input2\[0\]
rlabel metal1 10856 11254 10856 11254 0 CIRCUIT_1957.int_memory_1.GATES_8.input2\[1\]
rlabel via1 10442 12835 10442 12835 0 CIRCUIT_1957.int_memory_1.GATES_8.input2\[2\]
rlabel metal1 7544 11526 7544 11526 0 CIRCUIT_1957.int_memory_1.GATES_8.input2\[3\]
rlabel metal1 15870 17238 15870 17238 0 CIRCUIT_1957.int_memory_1.div_1.A0
rlabel metal2 21206 16728 21206 16728 0 CIRCUIT_1957.int_memory_1.div_1.A1
rlabel metal1 17112 16422 17112 16422 0 CIRCUIT_1957.int_memory_1.div_1.A2
rlabel metal2 21206 18224 21206 18224 0 CIRCUIT_1957.int_memory_1.div_1.A3
rlabel metal1 16146 21658 16146 21658 0 CIRCUIT_1957.int_memory_1.div_1.A4
rlabel metal2 16422 22440 16422 22440 0 CIRCUIT_1957.int_memory_1.div_1.A5
rlabel metal1 18078 21522 18078 21522 0 CIRCUIT_1957.int_memory_1.div_1.A6
rlabel metal1 20102 21930 20102 21930 0 CIRCUIT_1957.int_memory_1.div_1.A7
rlabel metal1 18676 21658 18676 21658 0 CIRCUIT_1957.int_memory_1.div_1.B0
rlabel metal2 19228 21692 19228 21692 0 CIRCUIT_1957.int_memory_1.div_1.B1
rlabel metal2 19320 20434 19320 20434 0 CIRCUIT_1957.int_memory_1.div_1.B2
rlabel metal1 21206 20468 21206 20468 0 CIRCUIT_1957.int_memory_1.div_1.B3
rlabel metal1 7130 22746 7130 22746 0 CIRCUIT_1957.int_memory_1.mul2_1.A0
rlabel metal1 8648 21930 8648 21930 0 CIRCUIT_1957.int_memory_1.mul2_1.A1
rlabel metal1 8970 23766 8970 23766 0 CIRCUIT_1957.int_memory_1.mul2_1.A2
rlabel metal2 9430 24463 9430 24463 0 CIRCUIT_1957.int_memory_1.mul2_1.A3
rlabel metal1 10028 24786 10028 24786 0 CIRCUIT_1957.int_memory_1.mul2_1.B0
rlabel metal2 9338 21828 9338 21828 0 CIRCUIT_1957.int_memory_1.mul2_1.B1
rlabel metal1 10948 22950 10948 22950 0 CIRCUIT_1957.int_memory_1.mul2_1.B2
rlabel metal2 11822 22134 11822 22134 0 CIRCUIT_1957.int_memory_1.mul2_1.B3
rlabel metal2 20838 6528 20838 6528 0 _0000_
rlabel metal1 14306 12138 14306 12138 0 _0001_
rlabel metal2 22310 7616 22310 7616 0 _0002_
rlabel metal1 21758 7310 21758 7310 0 _0003_
rlabel metal1 17763 14314 17763 14314 0 _0004_
rlabel metal2 16330 13056 16330 13056 0 _0005_
rlabel metal2 18170 11968 18170 11968 0 _0006_
rlabel metal1 16836 12750 16836 12750 0 _0007_
rlabel metal1 13938 9418 13938 9418 0 _0008_
rlabel metal1 19005 6698 19005 6698 0 _0009_
rlabel metal2 19090 7922 19090 7922 0 _0010_
rlabel metal1 16291 6698 16291 6698 0 _0011_
rlabel metal2 19458 7650 19458 7650 0 _0012_
rlabel metal2 11730 7990 11730 7990 0 _0013_
rlabel metal1 9476 7242 9476 7242 0 _0014_
rlabel metal1 12098 11016 12098 11016 0 _0015_
rlabel metal2 12006 9112 12006 9112 0 _0016_
rlabel metal1 18814 8534 18814 8534 0 _0017_
rlabel metal1 14858 5882 14858 5882 0 _0018_
rlabel metal1 4733 14314 4733 14314 0 _0027_
rlabel metal1 5423 13226 5423 13226 0 _0028_
rlabel metal1 6578 8942 6578 8942 0 _0029_
rlabel metal1 7217 9554 7217 9554 0 _0030_
rlabel metal2 4922 9962 4922 9962 0 _0031_
rlabel metal2 5566 9299 5566 9299 0 _0032_
rlabel metal1 2208 11866 2208 11866 0 _0033_
rlabel metal2 2714 13362 2714 13362 0 _0034_
rlabel metal2 2162 12002 2162 12002 0 _0035_
rlabel metal1 2208 18054 2208 18054 0 _0036_
rlabel metal1 2944 9146 2944 9146 0 _0037_
rlabel metal1 3864 8942 3864 8942 0 _0038_
rlabel metal1 4002 13838 4002 13838 0 _0039_
rlabel metal1 3680 8058 3680 8058 0 _0040_
rlabel metal1 2755 19822 2755 19822 0 _0041_
rlabel metal2 2806 19278 2806 19278 0 _0042_
rlabel via1 2341 17646 2341 17646 0 _0043_
rlabel metal2 2898 20213 2898 20213 0 _0044_
rlabel via2 10994 10693 10994 10693 0 _0045_
rlabel metal1 9230 11050 9230 11050 0 _0046_
rlabel metal1 9568 12614 9568 12614 0 _0047_
rlabel metal1 8234 10166 8234 10166 0 _0048_
rlabel viali 9609 11730 9609 11730 0 _0049_
rlabel metal2 10074 15266 10074 15266 0 _0050_
rlabel metal1 12604 13498 12604 13498 0 _0051_
rlabel metal2 12834 14110 12834 14110 0 _0052_
rlabel metal1 10018 3094 10018 3094 0 _0053_
rlabel metal1 9154 2618 9154 2618 0 _0054_
rlabel metal1 9798 2312 9798 2312 0 _0055_
rlabel metal2 12006 4012 12006 4012 0 _0056_
rlabel viali 15221 2346 15221 2346 0 _0057_
rlabel metal1 16417 3502 16417 3502 0 _0058_
rlabel metal1 18630 2618 18630 2618 0 _0059_
rlabel metal1 19836 4114 19836 4114 0 _0060_
rlabel metal1 9414 18326 9414 18326 0 _0061_
rlabel metal1 9844 17782 9844 17782 0 _0062_
rlabel metal1 12895 16490 12895 16490 0 _0063_
rlabel metal1 11960 18394 11960 18394 0 _0064_
rlabel via1 22305 4182 22305 4182 0 _0065_
rlabel metal1 22550 3502 22550 3502 0 _0066_
rlabel metal1 24564 2890 24564 2890 0 _0067_
rlabel metal1 23455 3094 23455 3094 0 _0068_
rlabel metal1 4595 21998 4595 21998 0 _0069_
rlabel metal1 4641 20434 4641 20434 0 _0070_
rlabel metal2 2070 22814 2070 22814 0 _0071_
rlabel metal1 2387 21930 2387 21930 0 _0072_
rlabel metal1 7079 18326 7079 18326 0 _0073_
rlabel via1 4917 17170 4917 17170 0 _0074_
rlabel metal1 6987 19414 6987 19414 0 _0075_
rlabel via1 5009 18734 5009 18734 0 _0076_
rlabel metal1 6746 22678 6746 22678 0 _0077_
rlabel via1 6757 21998 6757 21998 0 _0078_
rlabel metal2 9062 23970 9062 23970 0 _0079_
rlabel metal1 9016 23290 9016 23290 0 _0080_
rlabel via1 10262 20502 10262 20502 0 _0081_
rlabel metal2 7912 21556 7912 21556 0 _0082_
rlabel metal1 10207 21590 10207 21590 0 _0083_
rlabel metal1 12093 21590 12093 21590 0 _0084_
rlabel metal1 17332 16558 17332 16558 0 _0085_
rlabel metal1 16468 16218 16468 16218 0 _0086_
rlabel metal1 16095 16558 16095 16558 0 _0087_
rlabel metal1 16636 18326 16636 18326 0 _0088_
rlabel metal1 15405 22610 15405 22610 0 _0089_
rlabel via1 15313 21998 15313 21998 0 _0090_
rlabel metal2 17066 24310 17066 24310 0 _0091_
rlabel metal2 15778 23970 15778 23970 0 _0092_
rlabel metal2 17894 20978 17894 20978 0 _0093_
rlabel metal1 16136 19822 16136 19822 0 _0094_
rlabel metal1 18395 19414 18395 19414 0 _0095_
rlabel metal1 18032 18938 18032 18938 0 _0096_
rlabel metal1 7033 13294 7033 13294 0 _0097_
rlabel metal1 5096 14994 5096 14994 0 _0098_
rlabel metal1 19044 12614 19044 12614 0 _0099_
rlabel metal1 21344 10234 21344 10234 0 _0100_
rlabel metal1 20838 10064 20838 10064 0 _0101_
rlabel metal2 19918 14144 19918 14144 0 _0102_
rlabel metal1 20240 8942 20240 8942 0 _0103_
rlabel metal1 16238 5134 16238 5134 0 _0104_
rlabel metal2 19458 6052 19458 6052 0 _0105_
rlabel metal1 19780 3502 19780 3502 0 _0106_
rlabel metal1 20608 3026 20608 3026 0 _0107_
rlabel metal1 18998 2414 18998 2414 0 _0108_
rlabel metal2 20194 4692 20194 4692 0 _0109_
rlabel metal1 20562 4250 20562 4250 0 _0110_
rlabel metal2 20562 4318 20562 4318 0 _0111_
rlabel metal1 18538 2482 18538 2482 0 _0112_
rlabel metal1 16928 5882 16928 5882 0 _0113_
rlabel metal1 17940 6086 17940 6086 0 _0114_
rlabel metal1 20148 14994 20148 14994 0 _0115_
rlabel metal2 11178 13430 11178 13430 0 _0116_
rlabel metal1 14996 14314 14996 14314 0 _0117_
rlabel metal2 21114 14620 21114 14620 0 _0118_
rlabel metal2 2530 22406 2530 22406 0 _0119_
rlabel metal2 15870 9316 15870 9316 0 _0120_
rlabel metal1 18538 10778 18538 10778 0 _0121_
rlabel metal2 15870 6018 15870 6018 0 _0122_
rlabel metal2 18170 4964 18170 4964 0 _0123_
rlabel metal1 19458 3706 19458 3706 0 _0124_
rlabel metal2 17250 4624 17250 4624 0 _0125_
rlabel metal1 20746 9962 20746 9962 0 _0126_
rlabel metal1 18722 9384 18722 9384 0 _0127_
rlabel metal1 14950 9554 14950 9554 0 _0128_
rlabel metal1 16882 4114 16882 4114 0 _0129_
rlabel metal1 15226 3502 15226 3502 0 _0130_
rlabel metal1 15916 3706 15916 3706 0 _0131_
rlabel metal1 9200 4114 9200 4114 0 _0132_
rlabel metal2 11822 3638 11822 3638 0 _0133_
rlabel metal1 8878 5236 8878 5236 0 _0134_
rlabel metal1 9614 2448 9614 2448 0 _0135_
rlabel metal2 9430 5508 9430 5508 0 _0136_
rlabel metal2 8418 2244 8418 2244 0 _0137_
rlabel metal1 9292 3026 9292 3026 0 _0138_
rlabel metal1 9614 4556 9614 4556 0 _0139_
rlabel metal2 15042 6052 15042 6052 0 _0140_
rlabel metal1 16146 12750 16146 12750 0 _0141_
rlabel metal2 11362 11016 11362 11016 0 _0142_
rlabel metal1 15226 4488 15226 4488 0 _0143_
rlabel via2 18722 25653 18722 25653 0 _0144_
rlabel metal1 15962 25262 15962 25262 0 _0145_
rlabel metal2 17158 25738 17158 25738 0 _0146_
rlabel metal2 17618 25466 17618 25466 0 _0147_
rlabel metal2 16238 26044 16238 26044 0 _0148_
rlabel metal1 20930 7922 20930 7922 0 _0149_
rlabel metal2 17342 9180 17342 9180 0 _0150_
rlabel metal2 15686 8449 15686 8449 0 _0151_
rlabel metal1 6578 8398 6578 8398 0 _0152_
rlabel metal2 7314 7820 7314 7820 0 _0153_
rlabel metal1 7682 7854 7682 7854 0 _0154_
rlabel metal2 7774 8364 7774 8364 0 _0155_
rlabel metal1 8096 6970 8096 6970 0 _0156_
rlabel metal2 9338 8058 9338 8058 0 _0157_
rlabel metal1 8188 7990 8188 7990 0 _0158_
rlabel metal1 16606 6868 16606 6868 0 _0159_
rlabel metal1 20286 10982 20286 10982 0 _0160_
rlabel metal1 24610 9486 24610 9486 0 _0161_
rlabel metal1 16652 18734 16652 18734 0 _0162_
rlabel metal1 18400 20774 18400 20774 0 _0163_
rlabel metal2 19642 17442 19642 17442 0 _0164_
rlabel metal2 20378 17340 20378 17340 0 _0165_
rlabel metal2 20562 20366 20562 20366 0 _0166_
rlabel metal2 19826 19788 19826 19788 0 _0167_
rlabel metal1 20930 23052 20930 23052 0 _0168_
rlabel metal1 19550 20434 19550 20434 0 _0169_
rlabel metal1 19918 23120 19918 23120 0 _0170_
rlabel metal1 19136 24038 19136 24038 0 _0171_
rlabel metal1 18676 24174 18676 24174 0 _0172_
rlabel metal1 18446 22712 18446 22712 0 _0173_
rlabel metal1 18078 23086 18078 23086 0 _0174_
rlabel metal1 18032 23290 18032 23290 0 _0175_
rlabel metal2 18906 24412 18906 24412 0 _0176_
rlabel metal1 20470 21590 20470 21590 0 _0177_
rlabel metal1 20700 22202 20700 22202 0 _0178_
rlabel metal1 19550 21658 19550 21658 0 _0179_
rlabel metal2 19918 21828 19918 21828 0 _0180_
rlabel metal1 19688 21522 19688 21522 0 _0181_
rlabel metal1 19642 21590 19642 21590 0 _0182_
rlabel metal1 20286 22610 20286 22610 0 _0183_
rlabel metal1 21068 23086 21068 23086 0 _0184_
rlabel metal1 21620 23086 21620 23086 0 _0185_
rlabel metal2 18538 23936 18538 23936 0 _0186_
rlabel metal1 16514 20910 16514 20910 0 _0187_
rlabel metal2 18998 24072 18998 24072 0 _0188_
rlabel metal1 22034 23052 22034 23052 0 _0189_
rlabel metal2 22218 22406 22218 22406 0 _0190_
rlabel metal1 21735 23698 21735 23698 0 _0191_
rlabel metal1 20102 24378 20102 24378 0 _0192_
rlabel metal1 21390 24208 21390 24208 0 _0193_
rlabel metal1 21482 24752 21482 24752 0 _0194_
rlabel metal2 21298 23120 21298 23120 0 _0195_
rlabel metal1 23598 24344 23598 24344 0 _0196_
rlabel metal2 22770 24412 22770 24412 0 _0197_
rlabel metal1 22264 23086 22264 23086 0 _0198_
rlabel metal2 21666 20604 21666 20604 0 _0199_
rlabel metal2 23874 20570 23874 20570 0 _0200_
rlabel metal1 20286 20434 20286 20434 0 _0201_
rlabel metal1 24380 24174 24380 24174 0 _0202_
rlabel metal2 23138 24548 23138 24548 0 _0203_
rlabel metal1 24196 24582 24196 24582 0 _0204_
rlabel via1 25072 21998 25072 21998 0 _0205_
rlabel metal1 24794 19788 24794 19788 0 _0206_
rlabel metal1 23184 20910 23184 20910 0 _0207_
rlabel via1 23414 20995 23414 20995 0 _0208_
rlabel metal1 25116 20910 25116 20910 0 _0209_
rlabel metal2 21482 24174 21482 24174 0 _0210_
rlabel metal2 23874 23290 23874 23290 0 _0211_
rlabel metal1 24058 23052 24058 23052 0 _0212_
rlabel metal1 24380 21862 24380 21862 0 _0213_
rlabel metal1 24334 22406 24334 22406 0 _0214_
rlabel metal1 24610 21658 24610 21658 0 _0215_
rlabel metal1 25254 23018 25254 23018 0 _0216_
rlabel metal1 25162 23188 25162 23188 0 _0217_
rlabel metal1 25760 21998 25760 21998 0 _0218_
rlabel metal1 24380 21522 24380 21522 0 _0219_
rlabel metal1 23598 19856 23598 19856 0 _0220_
rlabel metal2 24058 20230 24058 20230 0 _0221_
rlabel metal1 26266 20400 26266 20400 0 _0222_
rlabel metal1 25300 21522 25300 21522 0 _0223_
rlabel metal1 23000 20570 23000 20570 0 _0224_
rlabel metal1 22770 20026 22770 20026 0 _0225_
rlabel metal1 25070 21386 25070 21386 0 _0226_
rlabel metal1 24840 21114 24840 21114 0 _0227_
rlabel metal1 25070 21454 25070 21454 0 _0228_
rlabel metal2 26358 21114 26358 21114 0 _0229_
rlabel metal2 27278 20230 27278 20230 0 _0230_
rlabel metal1 20194 19686 20194 19686 0 _0231_
rlabel via1 27186 19669 27186 19669 0 _0232_
rlabel metal1 25116 18734 25116 18734 0 _0233_
rlabel metal2 25898 18190 25898 18190 0 _0234_
rlabel metal1 23141 19686 23141 19686 0 _0235_
rlabel metal2 25990 18972 25990 18972 0 _0236_
rlabel metal1 26082 19380 26082 19380 0 _0237_
rlabel via1 27378 19414 27378 19414 0 _0238_
rlabel metal1 26312 21998 26312 21998 0 _0239_
rlabel metal1 26220 21862 26220 21862 0 _0240_
rlabel metal1 26542 21556 26542 21556 0 _0241_
rlabel metal1 26174 22542 26174 22542 0 _0242_
rlabel metal1 26496 22134 26496 22134 0 _0243_
rlabel metal2 27186 21318 27186 21318 0 _0244_
rlabel metal1 27324 19822 27324 19822 0 _0245_
rlabel metal1 26542 19754 26542 19754 0 _0246_
rlabel metal1 26266 17850 26266 17850 0 _0247_
rlabel metal2 27186 18122 27186 18122 0 _0248_
rlabel metal1 27186 17850 27186 17850 0 _0249_
rlabel metal2 27922 17646 27922 17646 0 _0250_
rlabel metal2 27094 16694 27094 16694 0 _0251_
rlabel metal2 26266 18666 26266 18666 0 _0252_
rlabel metal2 25622 17408 25622 17408 0 _0253_
rlabel metal1 26772 15674 26772 15674 0 _0254_
rlabel metal1 23736 17238 23736 17238 0 _0255_
rlabel metal1 25438 16660 25438 16660 0 _0256_
rlabel metal2 23230 18428 23230 18428 0 _0257_
rlabel metal2 23598 17952 23598 17952 0 _0258_
rlabel metal2 23782 17340 23782 17340 0 _0259_
rlabel metal1 26910 16592 26910 16592 0 _0260_
rlabel metal1 27646 20570 27646 20570 0 _0261_
rlabel metal2 27554 20196 27554 20196 0 _0262_
rlabel metal2 28106 20468 28106 20468 0 _0263_
rlabel metal1 27462 20332 27462 20332 0 _0264_
rlabel metal2 28014 18428 28014 18428 0 _0265_
rlabel metal1 27278 16592 27278 16592 0 _0266_
rlabel metal2 21666 16388 21666 16388 0 _0267_
rlabel metal1 21252 17034 21252 17034 0 _0268_
rlabel metal2 21390 16932 21390 16932 0 _0269_
rlabel metal2 20102 17408 20102 17408 0 _0270_
rlabel metal1 20700 16966 20700 16966 0 _0271_
rlabel metal1 24242 17714 24242 17714 0 _0272_
rlabel metal2 22862 17408 22862 17408 0 _0273_
rlabel metal1 22954 17680 22954 17680 0 _0274_
rlabel metal1 22126 16592 22126 16592 0 _0275_
rlabel metal2 22402 16762 22402 16762 0 _0276_
rlabel metal2 22770 16286 22770 16286 0 _0277_
rlabel metal2 24978 15674 24978 15674 0 _0278_
rlabel metal2 25806 15674 25806 15674 0 _0279_
rlabel metal2 25622 15300 25622 15300 0 _0280_
rlabel metal2 23966 15164 23966 15164 0 _0281_
rlabel metal2 23506 16048 23506 16048 0 _0282_
rlabel metal1 27600 16218 27600 16218 0 _0283_
rlabel metal2 28106 15810 28106 15810 0 _0284_
rlabel metal2 27370 15334 27370 15334 0 _0285_
rlabel metal1 27646 15674 27646 15674 0 _0286_
rlabel metal1 24196 16014 24196 16014 0 _0287_
rlabel metal1 22816 15606 22816 15606 0 _0288_
rlabel metal2 21574 15708 21574 15708 0 _0289_
rlabel metal1 22862 15096 22862 15096 0 _0290_
rlabel metal1 22908 16218 22908 16218 0 _0291_
rlabel metal1 21666 17578 21666 17578 0 _0292_
rlabel metal2 22862 15436 22862 15436 0 _0293_
rlabel metal2 21666 15708 21666 15708 0 _0294_
rlabel metal1 20516 18258 20516 18258 0 _0295_
rlabel metal2 14582 15674 14582 15674 0 _0296_
rlabel metal2 21206 15878 21206 15878 0 _0297_
rlabel metal2 13754 19924 13754 19924 0 _0298_
rlabel metal1 12742 25330 12742 25330 0 _0299_
rlabel metal1 10994 23664 10994 23664 0 _0300_
rlabel metal1 11914 23698 11914 23698 0 _0301_
rlabel metal2 12098 23290 12098 23290 0 _0302_
rlabel metal1 8802 25194 8802 25194 0 _0303_
rlabel metal2 9614 23460 9614 23460 0 _0304_
rlabel metal1 9154 24072 9154 24072 0 _0305_
rlabel metal2 8418 26656 8418 26656 0 _0306_
rlabel metal1 9246 24650 9246 24650 0 _0307_
rlabel metal1 9062 26282 9062 26282 0 _0308_
rlabel metal1 10856 25670 10856 25670 0 _0309_
rlabel metal1 10994 25806 10994 25806 0 _0310_
rlabel metal1 12144 24174 12144 24174 0 _0311_
rlabel metal1 13478 23222 13478 23222 0 _0312_
rlabel metal1 10764 23834 10764 23834 0 _0313_
rlabel metal1 9982 24174 9982 24174 0 _0314_
rlabel metal1 10672 23698 10672 23698 0 _0315_
rlabel metal2 11270 23290 11270 23290 0 _0316_
rlabel metal1 14398 22032 14398 22032 0 _0317_
rlabel viali 13017 20445 13017 20445 0 _0318_
rlabel metal2 9338 17408 9338 17408 0 _0319_
rlabel metal2 13938 15470 13938 15470 0 _0320_
rlabel metal2 12190 17068 12190 17068 0 _0321_
rlabel metal1 14444 5882 14444 5882 0 _0322_
rlabel metal1 5750 12886 5750 12886 0 _0323_
rlabel metal1 8602 17612 8602 17612 0 _0324_
rlabel metal1 6164 9554 6164 9554 0 _0325_
rlabel metal2 1794 10710 1794 10710 0 _0326_
rlabel metal2 16974 14314 16974 14314 0 _0327_
rlabel metal1 4784 8602 4784 8602 0 _0328_
rlabel metal1 7958 12410 7958 12410 0 _0329_
rlabel metal1 10856 13158 10856 13158 0 _0330_
rlabel metal1 16606 18394 16606 18394 0 _0331_
rlabel metal1 1886 12920 1886 12920 0 _0332_
rlabel metal1 16514 15640 16514 15640 0 _0333_
rlabel metal1 1840 14042 1840 14042 0 _0334_
rlabel metal1 4830 18292 4830 18292 0 _0335_
rlabel metal1 6532 18394 6532 18394 0 _0336_
rlabel metal1 15594 18870 15594 18870 0 _0337_
rlabel metal1 14858 21556 14858 21556 0 _0338_
rlabel metal1 14812 19822 14812 19822 0 _0339_
rlabel metal2 14950 20128 14950 20128 0 _0340_
rlabel metal2 13570 17408 13570 17408 0 _0341_
rlabel metal1 9430 15368 9430 15368 0 _0342_
rlabel metal2 13754 18836 13754 18836 0 _0343_
rlabel metal1 11730 19788 11730 19788 0 _0344_
rlabel metal1 12420 20026 12420 20026 0 _0345_
rlabel metal2 13386 20128 13386 20128 0 _0346_
rlabel metal1 13110 19822 13110 19822 0 _0347_
rlabel metal2 9982 26316 9982 26316 0 _0348_
rlabel metal1 10672 26554 10672 26554 0 _0349_
rlabel metal1 10810 26350 10810 26350 0 _0350_
rlabel metal2 12834 27200 12834 27200 0 _0351_
rlabel metal1 11960 26350 11960 26350 0 _0352_
rlabel metal2 12742 26418 12742 26418 0 _0353_
rlabel metal1 14122 26894 14122 26894 0 _0354_
rlabel metal1 13432 27030 13432 27030 0 _0355_
rlabel metal2 11178 26656 11178 26656 0 _0356_
rlabel metal1 12742 26350 12742 26350 0 _0357_
rlabel metal1 13248 25874 13248 25874 0 _0358_
rlabel metal1 9476 25806 9476 25806 0 _0359_
rlabel metal1 13248 25942 13248 25942 0 _0360_
rlabel metal2 13202 26180 13202 26180 0 _0361_
rlabel metal2 13018 27132 13018 27132 0 _0362_
rlabel metal2 13662 26010 13662 26010 0 _0363_
rlabel metal1 13892 24786 13892 24786 0 _0364_
rlabel metal1 14536 25942 14536 25942 0 _0365_
rlabel metal2 13386 24378 13386 24378 0 _0366_
rlabel metal1 13110 23154 13110 23154 0 _0367_
rlabel metal1 14030 21998 14030 21998 0 _0368_
rlabel metal1 13708 21590 13708 21590 0 _0369_
rlabel metal2 13570 24004 13570 24004 0 _0370_
rlabel metal1 13156 25466 13156 25466 0 _0371_
rlabel metal1 13662 26418 13662 26418 0 _0372_
rlabel metal1 14214 26758 14214 26758 0 _0373_
rlabel metal1 14674 20536 14674 20536 0 _0374_
rlabel metal1 14490 20366 14490 20366 0 _0375_
rlabel metal1 13386 19856 13386 19856 0 _0376_
rlabel via2 15870 13923 15870 13923 0 _0377_
rlabel metal1 16706 13974 16706 13974 0 _0378_
rlabel metal1 25484 8806 25484 8806 0 _0379_
rlabel metal1 25668 9146 25668 9146 0 _0380_
rlabel metal2 21574 18122 21574 18122 0 _0381_
rlabel metal1 21758 18258 21758 18258 0 _0382_
rlabel metal2 21298 18054 21298 18054 0 _0383_
rlabel metal1 20378 18394 20378 18394 0 _0384_
rlabel metal1 11178 20468 11178 20468 0 _0385_
rlabel metal2 12466 21182 12466 21182 0 _0386_
rlabel metal1 6578 13906 6578 13906 0 _0387_
rlabel via3 12765 22100 12765 22100 0 _0388_
rlabel metal1 11684 22202 11684 22202 0 _0389_
rlabel metal1 16974 22406 16974 22406 0 _0390_
rlabel metal1 11132 17170 11132 17170 0 _0391_
rlabel metal1 13248 17306 13248 17306 0 _0392_
rlabel metal1 13340 19482 13340 19482 0 _0393_
rlabel metal1 11224 20366 11224 20366 0 _0394_
rlabel metal2 12650 21284 12650 21284 0 _0395_
rlabel metal2 13018 21590 13018 21590 0 _0396_
rlabel metal2 18446 14450 18446 14450 0 _0397_
rlabel metal2 18814 14025 18814 14025 0 _0398_
rlabel via1 24786 9962 24786 9962 0 _0399_
rlabel metal1 24656 10234 24656 10234 0 _0400_
rlabel metal3 18975 15164 18975 15164 0 _0401_
rlabel metal1 18676 14858 18676 14858 0 _0402_
rlabel metal1 20148 16082 20148 16082 0 _0403_
rlabel metal1 20424 16014 20424 16014 0 _0404_
rlabel metal2 19458 15980 19458 15980 0 _0405_
rlabel metal2 19734 15742 19734 15742 0 _0406_
rlabel metal2 19550 15164 19550 15164 0 _0407_
rlabel metal1 8142 14858 8142 14858 0 _0408_
rlabel metal2 12558 17306 12558 17306 0 _0409_
rlabel metal1 9798 23494 9798 23494 0 _0410_
rlabel metal2 9706 20876 9706 20876 0 _0411_
rlabel metal1 5566 16422 5566 16422 0 _0412_
rlabel metal1 7268 17034 7268 17034 0 _0413_
rlabel metal1 10028 19686 10028 19686 0 _0414_
rlabel metal2 12466 17680 12466 17680 0 _0415_
rlabel metal2 14582 21495 14582 21495 0 _0416_
rlabel metal2 13478 20060 13478 20060 0 _0417_
rlabel via2 18722 16099 18722 16099 0 _0418_
rlabel metal1 19412 14926 19412 14926 0 _0419_
rlabel metal1 18630 15028 18630 15028 0 _0420_
rlabel metal2 18814 15198 18814 15198 0 _0421_
rlabel metal2 18170 14620 18170 14620 0 _0422_
rlabel metal1 24426 13906 24426 13906 0 _0423_
rlabel metal1 25208 12614 25208 12614 0 _0424_
rlabel metal2 24518 13532 24518 13532 0 _0425_
rlabel metal1 19458 19482 19458 19482 0 _0426_
rlabel metal1 19320 17306 19320 17306 0 _0427_
rlabel metal1 18262 17680 18262 17680 0 _0428_
rlabel metal2 14122 21794 14122 21794 0 _0429_
rlabel metal2 18354 17697 18354 17697 0 _0430_
rlabel metal1 19182 18292 19182 18292 0 _0431_
rlabel metal1 7498 12818 7498 12818 0 _0432_
rlabel metal1 7130 12682 7130 12682 0 _0433_
rlabel metal1 7498 15470 7498 15470 0 _0434_
rlabel metal2 8510 16082 8510 16082 0 _0435_
rlabel metal1 8602 16762 8602 16762 0 _0436_
rlabel metal1 19458 18190 19458 18190 0 _0437_
rlabel metal1 18676 17646 18676 17646 0 _0438_
rlabel metal2 18722 14722 18722 14722 0 _0439_
rlabel metal1 20286 15538 20286 15538 0 _0440_
rlabel metal2 20102 15334 20102 15334 0 _0441_
rlabel metal2 18906 14620 18906 14620 0 _0442_
rlabel metal1 21666 14382 21666 14382 0 _0443_
rlabel metal1 20194 14314 20194 14314 0 _0444_
rlabel metal1 21942 14314 21942 14314 0 _0445_
rlabel metal1 20608 13770 20608 13770 0 _0446_
rlabel metal1 21444 8874 21444 8874 0 _0447_
rlabel metal1 20930 10540 20930 10540 0 _0448_
rlabel metal1 20792 13158 20792 13158 0 _0449_
rlabel metal1 20838 13260 20838 13260 0 _0450_
rlabel metal2 25070 13668 25070 13668 0 _0451_
rlabel metal1 25438 13906 25438 13906 0 _0452_
rlabel metal1 24610 12716 24610 12716 0 _0453_
rlabel metal1 24886 11220 24886 11220 0 _0454_
rlabel metal1 25162 12750 25162 12750 0 _0455_
rlabel metal2 24978 9928 24978 9928 0 _0456_
rlabel metal2 24610 10064 24610 10064 0 _0457_
rlabel metal2 24886 9656 24886 9656 0 _0458_
rlabel metal2 24702 9350 24702 9350 0 _0459_
rlabel metal1 20286 12104 20286 12104 0 _0460_
rlabel metal1 20976 14518 20976 14518 0 _0461_
rlabel metal2 19734 13600 19734 13600 0 _0462_
rlabel metal1 20838 14790 20838 14790 0 _0463_
rlabel metal2 20010 12682 20010 12682 0 _0464_
rlabel metal1 21758 12818 21758 12818 0 _0465_
rlabel metal1 21436 12206 21436 12206 0 _0466_
rlabel metal1 20700 12206 20700 12206 0 _0467_
rlabel metal1 23414 12852 23414 12852 0 _0468_
rlabel metal1 19228 11118 19228 11118 0 _0469_
rlabel metal1 24518 13498 24518 13498 0 _0470_
rlabel via1 23703 12818 23703 12818 0 _0471_
rlabel metal1 23736 12410 23736 12410 0 _0472_
rlabel metal1 24932 12614 24932 12614 0 _0473_
rlabel metal2 23690 11322 23690 11322 0 _0474_
rlabel metal1 24472 10778 24472 10778 0 _0475_
rlabel metal1 24196 11118 24196 11118 0 _0476_
rlabel metal2 24702 11730 24702 11730 0 _0477_
rlabel metal1 23184 8058 23184 8058 0 _0478_
rlabel metal2 23138 9860 23138 9860 0 _0479_
rlabel metal2 23506 9146 23506 9146 0 _0480_
rlabel metal2 23874 9180 23874 9180 0 _0481_
rlabel metal1 19458 6800 19458 6800 0 _0482_
rlabel metal1 18400 12070 18400 12070 0 _0483_
rlabel viali 8426 6630 8426 6630 0 _0484_
rlabel metal1 7268 6970 7268 6970 0 _0485_
rlabel metal1 19596 7378 19596 7378 0 _0486_
rlabel metal2 16054 5644 16054 5644 0 _0487_
rlabel metal1 8510 5678 8510 5678 0 _0488_
rlabel metal2 12926 8704 12926 8704 0 _0489_
rlabel metal2 17802 8772 17802 8772 0 _0490_
rlabel metal1 18216 9690 18216 9690 0 _0491_
rlabel metal1 16560 11118 16560 11118 0 _0492_
rlabel metal1 17940 9962 17940 9962 0 _0493_
rlabel metal2 16698 10404 16698 10404 0 _0494_
rlabel metal1 21850 8466 21850 8466 0 _0495_
rlabel metal1 2254 6834 2254 6834 0 _0496_
rlabel metal1 8326 7412 8326 7412 0 _0497_
rlabel metal2 2530 9299 2530 9299 0 _0498_
rlabel metal1 2162 23664 2162 23664 0 _0499_
rlabel metal1 8096 19346 8096 19346 0 _0500_
rlabel metal1 5474 20570 5474 20570 0 _0501_
rlabel metal1 14536 13498 14536 13498 0 _0502_
rlabel metal2 13478 21556 13478 21556 0 _0503_
rlabel metal2 5658 14960 5658 14960 0 _0504_
rlabel metal1 5474 7378 5474 7378 0 _0505_
rlabel metal2 4186 15776 4186 15776 0 _0506_
rlabel metal2 1702 8772 1702 8772 0 _0507_
rlabel metal1 2024 20434 2024 20434 0 _0508_
rlabel metal2 10626 12444 10626 12444 0 _0509_
rlabel metal1 11408 17306 11408 17306 0 _0510_
rlabel metal1 20424 11866 20424 11866 0 _0511_
rlabel metal2 1702 13430 1702 13430 0 _0512_
rlabel metal2 14766 13906 14766 13906 0 _0513_
rlabel metal2 19642 19924 19642 19924 0 _0514_
rlabel metal2 2622 26010 2622 26010 0 _0515_
rlabel metal1 13386 12172 13386 12172 0 _0516_
rlabel metal1 15962 18224 15962 18224 0 _0517_
rlabel metal1 2346 22610 2346 22610 0 _0518_
rlabel metal2 15778 21284 15778 21284 0 _0519_
rlabel metal2 2714 6256 2714 6256 0 _0520_
rlabel metal1 13754 13498 13754 13498 0 _0521_
rlabel metal1 16767 22066 16767 22066 0 _0522_
rlabel metal1 7360 14382 7360 14382 0 _0523_
rlabel metal1 2346 21488 2346 21488 0 _0524_
rlabel metal3 7038 12444 7038 12444 0 _0525_
rlabel metal1 16882 10744 16882 10744 0 _0526_
rlabel metal1 22954 5202 22954 5202 0 _0527_
rlabel metal2 22954 4250 22954 4250 0 _0528_
rlabel metal1 23644 2278 23644 2278 0 _0529_
rlabel metal1 21942 2278 21942 2278 0 _0530_
rlabel metal1 2622 23086 2622 23086 0 _0531_
rlabel metal1 15548 18258 15548 18258 0 _0532_
rlabel metal1 18630 18734 18630 18734 0 _0533_
rlabel metal2 683 29308 683 29308 0 clk
rlabel metal1 10442 13974 10442 13974 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result
rlabel metal2 4370 19822 4370 19822 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result
rlabel metal2 7038 17034 7038 17034 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result
rlabel metal2 5290 23324 5290 23324 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result
rlabel metal1 10994 21862 10994 21862 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result
rlabel metal1 13110 17238 13110 17238 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result
rlabel metal1 14122 18258 14122 18258 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result
rlabel metal1 18124 20230 18124 20230 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result
rlabel metal2 7406 13600 7406 13600 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result
rlabel metal1 4370 10676 4370 10676 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result
rlabel metal1 3082 14790 3082 14790 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result
rlabel metal2 5290 11050 5290 11050 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result
rlabel metal2 2990 17374 2990 17374 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result
rlabel metal2 10442 13770 10442 13770 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result
rlabel metal2 11178 16252 11178 16252 0 clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result
rlabel metal1 13846 10030 13846 10030 0 clknet_0__0142_
rlabel metal2 16514 3774 16514 3774 0 clknet_0__0143_
rlabel metal1 7820 17170 7820 17170 0 clknet_0__0498_
rlabel metal1 13662 18666 13662 18666 0 clknet_0__0502_
rlabel metal1 17710 11050 17710 11050 0 clknet_0__0526_
rlabel metal2 13846 9826 13846 9826 0 clknet_0_clk
rlabel metal1 9016 10642 9016 10642 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result
rlabel metal1 3588 20366 3588 20366 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result
rlabel metal1 4692 17170 4692 17170 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result
rlabel metal1 6532 21998 6532 21998 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result
rlabel metal1 7866 21454 7866 21454 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result
rlabel metal1 16928 16626 16928 16626 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result
rlabel metal1 14904 21998 14904 21998 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result
rlabel metal2 15962 17748 15962 17748 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result
rlabel metal2 4738 13124 4738 13124 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result
rlabel metal2 6118 8500 6118 8500 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result
rlabel metal1 1978 13294 1978 13294 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result
rlabel metal2 2070 11492 2070 11492 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result
rlabel metal1 2116 17646 2116 17646 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result
rlabel metal1 8832 12954 8832 12954 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result
rlabel metal1 9384 18190 9384 18190 0 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result
rlabel metal1 15824 8330 15824 8330 0 clknet_1_0__leaf__0142_
rlabel metal1 10534 2414 10534 2414 0 clknet_1_0__leaf__0143_
rlabel metal1 2714 20468 2714 20468 0 clknet_1_0__leaf__0498_
rlabel metal2 12650 17748 12650 17748 0 clknet_1_0__leaf__0502_
rlabel metal1 18170 7786 18170 7786 0 clknet_1_0__leaf__0526_
rlabel metal1 2484 5338 2484 5338 0 clknet_1_0__leaf_clk
rlabel metal2 8602 12954 8602 12954 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result
rlabel metal1 2714 21896 2714 21896 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result
rlabel metal2 6762 18020 6762 18020 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result
rlabel metal1 7084 24174 7084 24174 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result
rlabel metal1 11132 20774 11132 20774 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result
rlabel metal1 15410 17102 15410 17102 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result
rlabel metal2 15226 23970 15226 23970 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result
rlabel metal2 16882 21284 16882 21284 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result
rlabel metal1 4692 14994 4692 14994 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result
rlabel metal2 4370 10948 4370 10948 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result
rlabel metal2 2070 16116 2070 16116 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result
rlabel metal1 5014 13974 5014 13974 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result
rlabel metal2 2070 20332 2070 20332 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result
rlabel metal2 11730 13668 11730 13668 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result
rlabel metal2 12742 16422 12742 16422 0 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result
rlabel metal1 13662 13260 13662 13260 0 clknet_1_1__leaf__0142_
rlabel metal1 14996 2414 14996 2414 0 clknet_1_1__leaf__0143_
rlabel metal2 13110 19346 13110 19346 0 clknet_1_1__leaf__0498_
rlabel metal1 15318 21522 15318 21522 0 clknet_1_1__leaf__0502_
rlabel metal1 15640 12818 15640 12818 0 clknet_1_1__leaf__0526_
rlabel via1 22034 4131 22034 4131 0 clknet_1_1__leaf_clk
rlabel metal2 6578 28373 6578 28373 0 io_in[0]
rlabel metal2 8602 28441 8602 28441 0 io_in[1]
rlabel metal1 11500 27438 11500 27438 0 io_in[2]
rlabel metal1 14076 27438 14076 27438 0 io_in[3]
rlabel metal1 16652 27438 16652 27438 0 io_in[4]
rlabel metal1 19182 27438 19182 27438 0 io_in[5]
rlabel metal1 21022 27574 21022 27574 0 io_in[6]
rlabel metal1 23506 27574 23506 27574 0 io_in[7]
rlabel metal1 25990 27574 25990 27574 0 io_in[8]
rlabel metal2 28382 28373 28382 28373 0 io_in[9]
rlabel metal2 598 1792 598 1792 0 io_out[0]
rlabel metal2 11638 1520 11638 1520 0 io_out[10]
rlabel metal1 12604 2822 12604 2822 0 io_out[11]
rlabel metal2 13846 1554 13846 1554 0 io_out[12]
rlabel metal1 17802 2312 17802 2312 0 io_out[13]
rlabel metal2 16054 823 16054 823 0 io_out[14]
rlabel metal2 17158 1792 17158 1792 0 io_out[15]
rlabel metal2 18262 1554 18262 1554 0 io_out[16]
rlabel metal2 19366 1656 19366 1656 0 io_out[17]
rlabel metal2 20470 1622 20470 1622 0 io_out[18]
rlabel metal2 21574 1690 21574 1690 0 io_out[19]
rlabel metal2 1702 1520 1702 1520 0 io_out[1]
rlabel metal1 22816 2822 22816 2822 0 io_out[20]
rlabel metal2 23782 1656 23782 1656 0 io_out[21]
rlabel metal2 2806 1520 2806 1520 0 io_out[2]
rlabel metal2 3910 1520 3910 1520 0 io_out[3]
rlabel metal1 14628 26282 14628 26282 0 net1
rlabel metal1 20861 26350 20861 26350 0 net10
rlabel metal1 20884 2414 20884 2414 0 net11
rlabel metal2 13386 4080 13386 4080 0 net12
rlabel metal2 11178 3842 11178 3842 0 net13
rlabel metal1 12098 3706 12098 3706 0 net14
rlabel metal1 12558 2414 12558 2414 0 net15
rlabel metal1 17618 2482 17618 2482 0 net16
rlabel metal2 16330 2516 16330 2516 0 net17
rlabel metal1 17710 3366 17710 3366 0 net18
rlabel metal1 18446 2278 18446 2278 0 net19
rlabel metal2 17802 26962 17802 26962 0 net2
rlabel metal1 19918 2414 19918 2414 0 net20
rlabel metal2 21390 3400 21390 3400 0 net21
rlabel metal1 23552 2414 23552 2414 0 net22
rlabel metal1 2070 2380 2070 2380 0 net23
rlabel metal1 21436 2550 21436 2550 0 net24
rlabel metal1 24242 2414 24242 2414 0 net25
rlabel metal1 3174 2482 3174 2482 0 net26
rlabel metal1 4278 2448 4278 2448 0 net27
rlabel metal2 5014 1588 5014 1588 0 net28
rlabel metal1 6348 2822 6348 2822 0 net29
rlabel metal2 17894 26758 17894 26758 0 net3
rlabel metal2 7222 1792 7222 1792 0 net30
rlabel metal1 8188 2822 8188 2822 0 net31
rlabel metal2 9430 1622 9430 1622 0 net32
rlabel metal2 10534 1656 10534 1656 0 net33
rlabel metal2 24886 1588 24886 1588 0 net34
rlabel metal2 25990 1588 25990 1588 0 net35
rlabel metal2 27094 1588 27094 1588 0 net36
rlabel metal2 28198 1588 28198 1588 0 net37
rlabel via2 28382 14909 28382 14909 0 net38
rlabel metal1 28842 2958 28842 2958 0 net39
rlabel metal1 15916 26418 15916 26418 0 net4
rlabel metal1 9200 2958 9200 2958 0 net40
rlabel metal1 9522 3570 9522 3570 0 net41
rlabel metal1 11040 2618 11040 2618 0 net42
rlabel metal2 10442 4250 10442 4250 0 net43
rlabel metal1 14950 2516 14950 2516 0 net44
rlabel metal1 15180 2618 15180 2618 0 net45
rlabel metal1 19274 3026 19274 3026 0 net46
rlabel metal1 20378 4046 20378 4046 0 net47
rlabel metal2 15318 26826 15318 26826 0 net5
rlabel metal2 17710 26826 17710 26826 0 net6
rlabel metal1 17894 26010 17894 26010 0 net7
rlabel metal1 16514 26316 16514 26316 0 net8
rlabel metal1 25852 26350 25852 26350 0 net9
rlabel metal1 3634 27574 3634 27574 0 rst
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
