module alu_mask_rom_32(
	input [4:0] op_size,
	
	output [31:0] mask_val
);

reg [31:0] rom_val;

assign mask_val = rom_val;

always @(*) begin
	case(op_size)
		0:  rom_val = 32'b00000000_00000000_00000000_00000001;
		1:  rom_val = 32'b00000000_00000000_00000000_00000011;
		2:  rom_val = 32'b00000000_00000000_00000000_00000111;
		3:  rom_val = 32'b00000000_00000000_00000000_00001111;
		4:  rom_val = 32'b00000000_00000000_00000000_00011111;
		5:  rom_val = 32'b00000000_00000000_00000000_00111111;
		6:  rom_val = 32'b00000000_00000000_00000000_01111111;
		7:  rom_val = 32'b00000000_00000000_00000000_11111111;
		8:  rom_val = 32'b00000000_00000000_00000001_11111111;
		9:  rom_val = 32'b00000000_00000000_00000011_11111111;
		10: rom_val = 32'b00000000_00000000_00000111_11111111;
		11: rom_val = 32'b00000000_00000000_00001111_11111111;
		12: rom_val = 32'b00000000_00000000_00011111_11111111;
		13: rom_val = 32'b00000000_00000000_00111111_11111111;
		14: rom_val = 32'b00000000_00000000_01111111_11111111;
		15: rom_val = 32'b00000000_00000000_11111111_11111111;
		16: rom_val = 32'b00000000_00000001_11111111_11111111;
		17: rom_val = 32'b00000000_00000011_11111111_11111111;
		18: rom_val = 32'b00000000_00000111_11111111_11111111;
		19: rom_val = 32'b00000000_00001111_11111111_11111111;
		20: rom_val = 32'b00000000_00011111_11111111_11111111;
		21: rom_val = 32'b00000000_00111111_11111111_11111111;
		22: rom_val = 32'b00000000_01111111_11111111_11111111;
		23: rom_val = 32'b00000000_11111111_11111111_11111111;
		24: rom_val = 32'b00000001_11111111_11111111_11111111;
		25: rom_val = 32'b00000011_11111111_11111111_11111111;
		26: rom_val = 32'b00000111_11111111_11111111_11111111;
		27: rom_val = 32'b00001111_11111111_11111111_11111111;
		28: rom_val = 32'b00011111_11111111_11111111_11111111;
		29: rom_val = 32'b00111111_11111111_11111111_11111111;
		30: rom_val = 32'b01111111_11111111_11111111_11111111;
		31: rom_val = 32'b11111111_11111111_11111111_11111111;
	endcase
end

endmodule

module alu_mask_rom_16(
	input [3:0] op_size,
	
	output [15:0] mask_val
);

reg [15:0] rom_val;

assign mask_val = rom_val;

always @(*) begin
	case(op_size)
		0:  rom_val = 16'b00000000_00000001;
		1:  rom_val = 16'b00000000_00000011;
		2:  rom_val = 16'b00000000_00000111;
		3:  rom_val = 16'b00000000_00001111;
		4:  rom_val = 16'b00000000_00011111;
		5:  rom_val = 32'b00000000_00111111;
		6:  rom_val = 16'b00000000_01111111;
		7:  rom_val = 16'b00000000_11111111;
		8:  rom_val = 16'b00000001_11111111;
		9:  rom_val = 16'b00000011_11111111;
		10: rom_val = 16'b00000111_11111111;
		11: rom_val = 16'b00001111_11111111;
		12: rom_val = 16'b00011111_11111111;
		13: rom_val = 16'b00111111_11111111;
		14: rom_val = 16'b01111111_11111111;
		15: rom_val = 16'b11111111_11111111;
	endcase
end

endmodule
