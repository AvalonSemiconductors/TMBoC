* NGSPICE file created from tt2_tholin_namebadge.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

.subckt tt2_tholin_namebadge clk io_in[0] io_in[1] io_in[2] io_oeb[0] io_oeb[10] io_oeb[11]
+ io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19]
+ io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ rst vccd1 vssd1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _429_/B _429_/D _655_/A _429_/C vssd1 vssd1 vccd1 vccd1 _638_/B sky130_fd_sc_hd__o31a_1
X_501_ _752_/Q _501_/B vssd1 vssd1 vccd1 vccd1 _501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__568__A1 _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_415_ _429_/D _426_/C _656_/B vssd1 vssd1 vccd1 vccd1 _417_/C sky130_fd_sc_hd__or3_2
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_680_ _680_/A _680_/B vssd1 vssd1 vccd1 vccd1 _683_/B sky130_fd_sc_hd__and2_1
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__622__B1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_732_ _728_/X _731_/A _769_/Q vssd1 vssd1 vccd1 vccd1 _769_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_663_ _382_/C _426_/D _434_/A vssd1 vssd1 vccd1 vccd1 _664_/C sky130_fd_sc_hd__a21o_2
X_594_ _474_/A _567_/X _625_/A vssd1 vssd1 vccd1 vccd1 _595_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__598__C1 _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout20_A _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput7 _798_/X vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_4
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_715_ _684_/A _754_/D _714_/Y _737_/A vssd1 vssd1 vccd1 vccd1 _763_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_646_ _644_/X _645_/X _657_/B vssd1 vssd1 vccd1 vccd1 _646_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_577_ _750_/D _577_/B _585_/B _577_/D vssd1 vssd1 vccd1 vccd1 _577_/X sky130_fd_sc_hd__and4_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_500_ _474_/Y _625_/B _496_/X vssd1 vssd1 vccd1 vccd1 _500_/X sky130_fd_sc_hd__a21o_1
X_431_ _434_/A _434_/B vssd1 vssd1 vccd1 vccd1 _431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_629_ _751_/D _626_/X _628_/X vssd1 vssd1 vccd1 vccd1 _629_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_414_ _685_/A _656_/B vssd1 vssd1 vccd1 vccd1 _655_/B sky130_fd_sc_hd__nor2_1
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__405__A _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__503__A _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_662_ _760_/Q _756_/Q _678_/A vssd1 vssd1 vccd1 vccd1 _662_/X sky130_fd_sc_hd__mux2_4
X_731_ _731_/A _731_/B vssd1 vssd1 vccd1 vccd1 _768_/D sky130_fd_sc_hd__and2_1
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_593_ _751_/D _593_/B _593_/C vssd1 vssd1 vccd1 vccd1 _593_/Y sky130_fd_sc_hd__nor3_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput8 _739_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_4
Xoutput10 _741_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_4
X_645_ _408_/Y _636_/X _638_/A vssd1 vssd1 vccd1 vccd1 _645_/X sky130_fd_sc_hd__a21bo_1
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_714_ _723_/A _714_/B vssd1 vssd1 vccd1 vccd1 _714_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_576_ _510_/A _589_/A _551_/Y _584_/B vssd1 vssd1 vccd1 vccd1 _576_/X sky130_fd_sc_hd__a31o_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_430_ _430_/A _655_/C vssd1 vssd1 vccd1 vccd1 _430_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__662__S _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_628_ _589_/Y _614_/X _627_/X _610_/B vssd1 vssd1 vccd1 vccd1 _628_/X sky130_fd_sc_hd__o211a_1
X_559_ _555_/X _556_/X _558_/X _547_/A vssd1 vssd1 vccd1 vccd1 _559_/X sky130_fd_sc_hd__o211a_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_413_ _744_/Q _745_/Q vssd1 vssd1 vccd1 vccd1 _418_/B sky130_fd_sc_hd__xor2_4
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__707__B1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__722__A3 _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__622__A2 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_661_ _652_/X _659_/X _660_/Y _453_/A _798_/A vssd1 vssd1 vccd1 vccd1 _738_/D sky130_fd_sc_hd__a32o_1
X_730_ _737_/A _728_/C _768_/Q vssd1 vssd1 vccd1 vccd1 _731_/B sky130_fd_sc_hd__a21o_1
X_592_ _510_/A _596_/B _577_/B _585_/B _558_/A vssd1 vssd1 vccd1 vccd1 _593_/C sky130_fd_sc_hd__o2111a_1
XFILLER_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__513__A1 _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput9 _740_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_4
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput11 _748_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_4
X_575_ _533_/A _574_/X _533_/X vssd1 vssd1 vccd1 vccd1 _575_/Y sky130_fd_sc_hd__a21boi_1
X_644_ _426_/C _656_/B _664_/A _643_/X _426_/D vssd1 vssd1 vccd1 vccd1 _644_/X sky130_fd_sc_hd__o221a_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_713_ _712_/B _754_/D _723_/A _712_/Y vssd1 vssd1 vccd1 vccd1 _762_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_627_ _596_/A _545_/B _545_/A vssd1 vssd1 vccd1 vccd1 _627_/X sky130_fd_sc_hd__a21o_1
X_558_ _558_/A _558_/B _558_/C vssd1 vssd1 vccd1 vccd1 _558_/X sky130_fd_sc_hd__or3_1
X_489_ _749_/Q _750_/Q _751_/Q _489_/D vssd1 vssd1 vccd1 vccd1 _501_/B sky130_fd_sc_hd__or4_2
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_412_ _745_/Q _744_/Q vssd1 vssd1 vccd1 vccd1 _412_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__517__A _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_660_ _712_/A _660_/B vssd1 vssd1 vccd1 vccd1 _660_/Y sky130_fd_sc_hd__nor2_2
X_591_ _749_/D _589_/B _590_/X _750_/D vssd1 vssd1 vccd1 vccd1 _593_/B sky130_fd_sc_hd__o211a_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput12 _798_/A vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_4
XANTENNA__514__B _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_712_ _712_/A _712_/B vssd1 vssd1 vccd1 vccd1 _712_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_643_ _684_/A _743_/Q _742_/Q _685_/A vssd1 vssd1 vccd1 vccd1 _643_/X sky130_fd_sc_hd__o22a_1
X_574_ _610_/A _514_/D _567_/X _584_/B vssd1 vssd1 vccd1 vccd1 _574_/X sky130_fd_sc_hd__a31o_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_626_ _545_/A _605_/X _625_/Y _624_/X _483_/Y vssd1 vssd1 vccd1 vccd1 _626_/X sky130_fd_sc_hd__a32o_1
XANTENNA__435__A _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_557_ _541_/B _514_/D _480_/A _480_/B vssd1 vssd1 vccd1 vccd1 _558_/C sky130_fd_sc_hd__a211oi_2
X_488_ _589_/A _530_/B _625_/A _483_/Y vssd1 vssd1 vccd1 vccd1 _488_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__661__B2 _798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_411_ _745_/Q _744_/Q vssd1 vssd1 vccd1 vccd1 _430_/A sky130_fd_sc_hd__and2b_4
X_609_ _610_/B _609_/B vssd1 vssd1 vccd1 vccd1 _609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__641__A1_N _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__540__A3 _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_590_ _462_/A _544_/A _573_/C _514_/A _584_/A vssd1 vssd1 vccd1 vccd1 _590_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_642_ _428_/Y _636_/X _641_/X _421_/X _412_/Y vssd1 vssd1 vccd1 vccd1 _642_/X sky130_fd_sc_hd__a221o_1
X_711_ _418_/B _706_/X _709_/X _745_/Q vssd1 vssd1 vccd1 vccd1 _745_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_573_ _746_/D _748_/D _573_/C vssd1 vssd1 vccd1 vccd1 _584_/B sky130_fd_sc_hd__and3_2
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__541__A _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_625_ _625_/A _625_/B vssd1 vssd1 vccd1 vccd1 _625_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__422__A2 _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_487_ _551_/A _544_/A vssd1 vssd1 vccd1 vccd1 _530_/B sky130_fd_sc_hd__nand2_4
X_556_ _618_/A _498_/Y _585_/A vssd1 vssd1 vccd1 vccd1 _556_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__716__A3 _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_410_ _664_/B vssd1 vssd1 vccd1 vccd1 _410_/Y sky130_fd_sc_hd__inv_2
X_608_ _561_/X _607_/X _606_/X _750_/D vssd1 vssd1 vccd1 vccd1 _609_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA__446__A _748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_539_ _749_/D _577_/B _530_/B _750_/D vssd1 vssd1 vccd1 vccd1 _539_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_572_ _616_/B _571_/X _560_/X vssd1 vssd1 vccd1 vccd1 _757_/D sky130_fd_sc_hd__o21a_1
X_641_ _678_/A _435_/B _639_/X _640_/X vssd1 vssd1 vccd1 vccd1 _641_/X sky130_fd_sc_hd__a2bb2o_1
X_710_ _706_/X _709_/X _744_/Q vssd1 vssd1 vccd1 vccd1 _744_/D sky130_fd_sc_hd__mux2_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__541__B _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_624_ _746_/D _585_/B _749_/D vssd1 vssd1 vccd1 vccd1 _624_/X sky130_fd_sc_hd__a21o_1
X_555_ _552_/C _618_/B _610_/A _552_/B vssd1 vssd1 vccd1 vccd1 _555_/X sky130_fd_sc_hd__o211a_1
XANTENNA__591__C1 _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_486_ _747_/Q _577_/B vssd1 vssd1 vccd1 vccd1 _625_/A sky130_fd_sc_hd__or2_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_538_ _616_/B _532_/Y _533_/X _537_/X vssd1 vssd1 vccd1 vccd1 _538_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_607_ _589_/A _618_/C _618_/B _533_/A vssd1 vssd1 vccd1 vccd1 _607_/X sky130_fd_sc_hd__a211o_1
X_469_ _443_/X _470_/B _495_/B _445_/X _493_/C vssd1 vssd1 vccd1 vccd1 _520_/A sky130_fd_sc_hd__a2111o_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__372__A _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__546__C1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__537__C1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_640_ _636_/X _637_/Y _638_/Y vssd1 vssd1 vccd1 vccd1 _640_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_571_ _492_/Y _562_/X _563_/X _570_/X vssd1 vssd1 vccd1 vccd1 _571_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__673__A1 _739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_769_ _769_/CLK _769_/D vssd1 vssd1 vccd1 vccd1 _769_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__375__A _748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_554_ _558_/A _549_/X _550_/X _552_/Y _553_/X vssd1 vssd1 vccd1 vccd1 _554_/X sky130_fd_sc_hd__o32a_1
X_485_ _564_/A _493_/B _493_/C _493_/D vssd1 vssd1 vccd1 vccd1 _577_/B sky130_fd_sc_hd__or4_4
X_623_ _547_/A _620_/X _621_/X _622_/X vssd1 vssd1 vccd1 vccd1 _623_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_537_ _533_/A _536_/B _534_/X _752_/D vssd1 vssd1 vccd1 vccd1 _537_/X sky130_fd_sc_hd__o211a_1
X_606_ _747_/D _530_/A _484_/Y _597_/A vssd1 vssd1 vccd1 vccd1 _606_/X sky130_fd_sc_hd__a31o_1
X_468_ _470_/A _493_/D _471_/C vssd1 vssd1 vccd1 vccd1 _610_/A sky130_fd_sc_hd__or3_4
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_399_ _680_/A _678_/B vssd1 vssd1 vccd1 vccd1 _399_/X sky130_fd_sc_hd__and2_1
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__555__B1 _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_570_ _496_/X _565_/X _569_/X _547_/A vssd1 vssd1 vccd1 vccd1 _570_/X sky130_fd_sc_hd__o211a_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_768_ _769_/CLK _768_/D vssd1 vssd1 vccd1 vccd1 _768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_699_ _678_/B _449_/Y _692_/B _678_/Y vssd1 vssd1 vccd1 vccd1 _699_/X sky130_fd_sc_hd__a31o_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__391__A _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_622_ _545_/A _480_/B _751_/D vssd1 vssd1 vccd1 vccd1 _622_/X sky130_fd_sc_hd__a21o_1
XANTENNA__566__A _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_553_ _552_/B _541_/B _551_/Y _585_/A vssd1 vssd1 vccd1 vccd1 _553_/X sky130_fd_sc_hd__a31o_1
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_484_ _746_/D _544_/A vssd1 vssd1 vccd1 vccd1 _484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__591__A1 _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__386__A _769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_605_ _747_/D _484_/Y _749_/D vssd1 vssd1 vccd1 vccd1 _605_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_536_ _536_/A _536_/B vssd1 vssd1 vccd1 vccd1 _536_/Y sky130_fd_sc_hd__nor2_1
X_398_ _394_/Y _704_/A _396_/Y _383_/X _397_/X vssd1 vssd1 vccd1 vccd1 _678_/B sky130_fd_sc_hd__a221o_4
X_467_ _470_/A _746_/D vssd1 vssd1 vccd1 vccd1 _552_/A sky130_fd_sc_hd__nor2_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout40 _764_/Q vssd1 vssd1 vccd1 vccd1 _426_/C sky130_fd_sc_hd__buf_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_519_ _520_/A _566_/B vssd1 vssd1 vccd1 vccd1 _618_/B sky130_fd_sc_hd__and2_2
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__700__A1 _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__484__A _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__437__B1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ _769_/CLK _767_/D vssd1 vssd1 vccd1 vccd1 _767_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_698_ _412_/Y _695_/X _697_/X _406_/S vssd1 vssd1 vccd1 vccd1 _698_/X sky130_fd_sc_hd__o211a_1
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_621_ _509_/Y _558_/B _533_/A vssd1 vssd1 vccd1 vccd1 _621_/X sky130_fd_sc_hd__o21a_1
X_483_ _474_/Y _596_/B _545_/A vssd1 vssd1 vccd1 vccd1 _483_/Y sky130_fd_sc_hd__a21oi_2
X_552_ _552_/A _552_/B _552_/C _618_/B vssd1 vssd1 vccd1 vccd1 _552_/Y sky130_fd_sc_hd__nor4_1
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_604_ _616_/B _599_/X _601_/X _603_/X vssd1 vssd1 vccd1 vccd1 _759_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__577__A _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _770_/CLK sky130_fd_sc_hd__clkbuf_16
X_535_ _474_/Y _748_/D _530_/A _577_/B _480_/B vssd1 vssd1 vccd1 vccd1 _536_/B sky130_fd_sc_hd__o32a_1
X_466_ _584_/A vssd1 vssd1 vccd1 vccd1 _747_/D sky130_fd_sc_hd__inv_2
X_397_ _433_/A _403_/B _429_/B vssd1 vssd1 vccd1 vccd1 _397_/X sky130_fd_sc_hd__or3b_1
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout30 _433_/A vssd1 vssd1 vccd1 vccd1 _434_/A sky130_fd_sc_hd__buf_4
Xfanout41 _764_/Q vssd1 vssd1 vccd1 vccd1 _685_/A sky130_fd_sc_hd__buf_4
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_518_ _520_/A _566_/B vssd1 vssd1 vccd1 vccd1 _552_/C sky130_fd_sc_hd__nor2_2
X_449_ _403_/B _648_/B _769_/Q vssd1 vssd1 vccd1 vccd1 _449_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__680__A _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__667__A1 _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_766_ _769_/CLK _766_/D vssd1 vssd1 vccd1 vccd1 _766_/Q sky130_fd_sc_hd__dfxtp_1
X_697_ _692_/B _696_/X _647_/X vssd1 vssd1 vccd1 vccd1 _697_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_551_ _551_/A _566_/B vssd1 vssd1 vccd1 vccd1 _551_/Y sky130_fd_sc_hd__nand2_2
X_620_ _533_/A _585_/C _597_/Y _618_/X _619_/X vssd1 vssd1 vccd1 vccd1 _620_/X sky130_fd_sc_hd__a32o_1
XFILLER_8_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_482_ _749_/Q _489_/D _475_/X _493_/C vssd1 vssd1 vccd1 vccd1 _596_/B sky130_fd_sc_hd__a31o_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__567__B1 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_749_ _762_/CLK _749_/D vssd1 vssd1 vccd1 vccd1 _749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_603_ _547_/A _602_/X _752_/D vssd1 vssd1 vccd1 vccd1 _603_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_465_ _495_/B _495_/C vssd1 vssd1 vccd1 vccd1 _584_/A sky130_fd_sc_hd__nor2_8
XANTENNA__593__A _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_534_ _618_/A _589_/B _499_/X _514_/X _558_/A vssd1 vssd1 vccd1 vccd1 _534_/X sky130_fd_sc_hd__a311o_1
X_396_ _429_/D _656_/B vssd1 vssd1 vccd1 vccd1 _396_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__678__A _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout20 _750_/D vssd1 vssd1 vccd1 vccd1 _533_/A sky130_fd_sc_hd__buf_4
Xfanout31 _769_/Q vssd1 vssd1 vccd1 vccd1 _433_/A sky130_fd_sc_hd__buf_4
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout42 _763_/Q vssd1 vssd1 vccd1 vccd1 _656_/B sky130_fd_sc_hd__buf_4
X_448_ _656_/C _426_/D _417_/C _434_/A vssd1 vssd1 vccd1 vccd1 _448_/X sky130_fd_sc_hd__a31o_2
X_517_ _751_/D _517_/B vssd1 vssd1 vccd1 vccd1 _517_/X sky130_fd_sc_hd__and2_1
X_379_ _434_/A _429_/C vssd1 vssd1 vccd1 vccd1 _657_/B sky130_fd_sc_hd__or2_4
XANTENNA__498__A _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__630__S _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__751__D _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__667__A2 _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_765_ _769_/CLK _765_/D vssd1 vssd1 vccd1 vccd1 _765_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_696_ _403_/B _664_/B _648_/Y vssd1 vssd1 vccd1 vccd1 _696_/X sky130_fd_sc_hd__a21o_1
XANTENNA__746__D _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_550_ _552_/C _618_/B _552_/B vssd1 vssd1 vccd1 vccd1 _550_/X sky130_fd_sc_hd__o21a_1
X_481_ _552_/B vssd1 vssd1 vccd1 vccd1 _481_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_679_ _678_/B _449_/Y _675_/X _678_/Y vssd1 vssd1 vccd1 vccd1 _680_/B sky130_fd_sc_hd__a31o_1
X_748_ _762_/CLK _748_/D vssd1 vssd1 vccd1 vccd1 _748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_602_ _750_/D _596_/B _584_/B _589_/Y _610_/C vssd1 vssd1 vccd1 vccd1 _602_/X sky130_fd_sc_hd__o32a_1
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_533_ _533_/A _573_/C _589_/B vssd1 vssd1 vccd1 vccd1 _533_/X sky130_fd_sc_hd__or3_1
X_464_ _445_/C _452_/C _452_/A _452_/B vssd1 vssd1 vccd1 vccd1 _495_/C sky130_fd_sc_hd__o211a_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_395_ _655_/A _426_/C vssd1 vssd1 vccd1 vccd1 _704_/A sky130_fd_sc_hd__nand2_2
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__678__B _678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout21 _536_/A vssd1 vssd1 vccd1 vccd1 _750_/D sky130_fd_sc_hd__buf_4
Xfanout32 _403_/B vssd1 vssd1 vccd1 vccd1 _429_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__703__B2 _741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout43 _763_/Q vssd1 vssd1 vccd1 vccd1 _684_/A sky130_fd_sc_hd__clkbuf_4
X_378_ _433_/A _403_/B vssd1 vssd1 vccd1 vccd1 _653_/B sky130_fd_sc_hd__nor2_2
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_447_ _749_/Q _750_/Q _489_/D vssd1 vssd1 vccd1 vccd1 _455_/A sky130_fd_sc_hd__nor3_2
X_516_ _510_/A _558_/B _514_/X _585_/A vssd1 vssd1 vccd1 vccd1 _517_/B sky130_fd_sc_hd__a211o_1
XANTENNA__498__B _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__449__B1 _769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__749__D _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__603__B1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__521__C1 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_764_ _770_/CLK _764_/D vssd1 vssd1 vccd1 vccd1 _764_/Q sky130_fd_sc_hd__dfxtp_1
X_695_ _428_/Y _692_/B _694_/X _421_/X vssd1 vssd1 vccd1 vccd1 _695_/X sky130_fd_sc_hd__a22o_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_480_ _480_/A _480_/B vssd1 vssd1 vccd1 vccd1 _480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_747_ _758_/CLK _747_/D vssd1 vssd1 vccd1 vccd1 _747_/Q sky130_fd_sc_hd__dfxtp_4
X_678_ _678_/A _678_/B vssd1 vssd1 vccd1 vccd1 _678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_601_ _533_/A _600_/X _536_/Y _751_/D vssd1 vssd1 vccd1 vccd1 _601_/X sky130_fd_sc_hd__a211o_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_394_ _656_/B _429_/D vssd1 vssd1 vccd1 vccd1 _394_/Y sky130_fd_sc_hd__nand2b_1
X_463_ _393_/X _453_/B _444_/B _747_/Q vssd1 vssd1 vccd1 vccd1 _495_/B sky130_fd_sc_hd__o31a_4
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_532_ _530_/X _531_/X _505_/X vssd1 vssd1 vccd1 vccd1 _532_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout22 _480_/Y vssd1 vssd1 vccd1 vccd1 _552_/B sky130_fd_sc_hd__buf_4
Xfanout33 _768_/Q vssd1 vssd1 vccd1 vccd1 _403_/B sky130_fd_sc_hd__buf_4
Xfanout44 _712_/B vssd1 vssd1 vccd1 vccd1 _678_/A sky130_fd_sc_hd__buf_6
Xtt2_tholin_namebadge_70 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_70/HI io_oeb[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_515_ _493_/C _480_/B _514_/D vssd1 vssd1 vccd1 vccd1 _558_/B sky130_fd_sc_hd__o21a_4
X_377_ _429_/D _655_/A vssd1 vssd1 vccd1 vccd1 _656_/C sky130_fd_sc_hd__or2_4
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_446_ _748_/Q _453_/A _453_/B _445_/C vssd1 vssd1 vccd1 vccd1 _489_/D sky130_fd_sc_hd__or4b_4
XANTENNA__458__A1 _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__612__B2 _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_429_ _434_/A _429_/B _429_/C _429_/D vssd1 vssd1 vccd1 vccd1 _655_/C sky130_fd_sc_hd__or4_2
XANTENNA__679__A1 _678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 _632_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__521__B1 _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_694_ _689_/Y _692_/X _693_/X vssd1 vssd1 vccd1 vccd1 _694_/X sky130_fd_sc_hd__a21bo_1
X_763_ _770_/CLK _763_/D vssd1 vssd1 vccd1 vccd1 _763_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_677_ _431_/Y _674_/Y _675_/X _676_/X vssd1 vssd1 vccd1 vccd1 _677_/X sky130_fd_sc_hd__a2bb2o_1
X_746_ _762_/CLK _746_/D vssd1 vssd1 vccd1 vccd1 _746_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_output11_A _748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__798__A _798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_600_ _618_/A _524_/Y _551_/Y _561_/X _498_/Y vssd1 vssd1 vccd1 vccd1 _600_/X sky130_fd_sc_hd__a32o_1
XFILLER_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_531_ _589_/A _618_/C _455_/Y vssd1 vssd1 vccd1 vccd1 _531_/X sky130_fd_sc_hd__a21o_1
X_462_ _462_/A vssd1 vssd1 vccd1 vccd1 _746_/D sky130_fd_sc_hd__clkinv_4
X_393_ _754_/D _660_/B vssd1 vssd1 vccd1 vccd1 _393_/X sky130_fd_sc_hd__or2_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_729_ _712_/A _737_/B _728_/X vssd1 vssd1 vccd1 vccd1 _731_/A sky130_fd_sc_hd__a21oi_1
Xfanout34 _656_/A vssd1 vssd1 vccd1 vccd1 _429_/B sky130_fd_sc_hd__buf_4
Xfanout45 _762_/Q vssd1 vssd1 vccd1 vccd1 _712_/B sky130_fd_sc_hd__clkbuf_8
Xfanout23 _480_/Y vssd1 vssd1 vccd1 vccd1 _530_/A sky130_fd_sc_hd__buf_2
Xtt2_tholin_namebadge_60 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_60/HI io_oeb[13]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_71 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_71/HI io_oeb[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_514_ _514_/A _746_/D _573_/C _514_/D vssd1 vssd1 vccd1 vccd1 _514_/X sky130_fd_sc_hd__and4_2
X_445_ _452_/A _452_/B _445_/C vssd1 vssd1 vccd1 vccd1 _445_/X sky130_fd_sc_hd__and3_1
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_376_ _754_/Q _737_/B vssd1 vssd1 vccd1 vccd1 _754_/D sky130_fd_sc_hd__nor2_8
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_428_ _429_/B _429_/D _657_/B vssd1 vssd1 vccd1 vccd1 _428_/Y sky130_fd_sc_hd__nor3_4
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 _634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__579__A1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_693_ _678_/A _424_/Y _431_/Y _433_/Y _435_/B vssd1 vssd1 vccd1 vccd1 _693_/X sky130_fd_sc_hd__o41a_1
X_762_ _762_/CLK _762_/D vssd1 vssd1 vccd1 vccd1 _762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__497__B1 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_676_ _637_/A _435_/B _692_/A _637_/B _428_/Y vssd1 vssd1 vccd1 vccd1 _676_/X sky130_fd_sc_hd__a41o_1
X_745_ _770_/CLK _745_/D vssd1 vssd1 vccd1 vccd1 _745_/Q sky130_fd_sc_hd__dfxtp_4
X_461_ _493_/D _471_/C vssd1 vssd1 vccd1 vccd1 _462_/A sky130_fd_sc_hd__nor2_4
X_530_ _530_/A _530_/B _530_/C vssd1 vssd1 vccd1 vccd1 _530_/X sky130_fd_sc_hd__and3_1
X_392_ _754_/D _660_/B vssd1 vssd1 vccd1 vccd1 _452_/A sky130_fd_sc_hd__nor2_4
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_659_ _658_/B _684_/A _659_/S vssd1 vssd1 vccd1 vccd1 _659_/X sky130_fd_sc_hd__mux2_1
X_728_ _737_/A _768_/Q _728_/C vssd1 vssd1 vccd1 vccd1 _728_/X sky130_fd_sc_hd__and3_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 _492_/Y vssd1 vssd1 vccd1 vccd1 _751_/D sky130_fd_sc_hd__buf_4
Xfanout24 _748_/D vssd1 vssd1 vccd1 vccd1 _566_/B sky130_fd_sc_hd__buf_4
Xfanout35 _705_/A vssd1 vssd1 vccd1 vccd1 _656_/A sky130_fd_sc_hd__buf_4
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout46 _754_/Q vssd1 vssd1 vccd1 vccd1 _737_/A sky130_fd_sc_hd__clkbuf_4
Xtt2_tholin_namebadge_50 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_50/HI io_oeb[3]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_72 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_72/HI io_oeb[25]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_61 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_61/HI io_oeb[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__624__B1 _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_444_ _747_/Q _444_/B vssd1 vssd1 vccd1 vccd1 _445_/C sky130_fd_sc_hd__nor2_2
X_513_ _541_/B _625_/B _509_/Y _530_/B _545_/A vssd1 vssd1 vccd1 vccd1 _513_/X sky130_fd_sc_hd__a221o_1
X_375_ _748_/Q vssd1 vssd1 vccd1 vccd1 _564_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__560__C1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_427_ _439_/A _439_/B _426_/X _430_/A _421_/X vssd1 vssd1 vccd1 vccd1 _427_/Y sky130_fd_sc_hd__o311ai_4
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 _632_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__610__A _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_761_ _762_/CLK _761_/D vssd1 vssd1 vccd1 vccd1 _761_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_692_ _692_/A _692_/B vssd1 vssd1 vccd1 vccd1 _692_/X sky130_fd_sc_hd__and2_1
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__430__A _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout16_A _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__497__A1 _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_744_ _769_/CLK _744_/D vssd1 vssd1 vccd1 vccd1 _744_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_675_ _761_/Q _757_/Q _678_/A vssd1 vssd1 vccd1 vccd1 _675_/X sky130_fd_sc_hd__mux2_2
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_460_ _442_/C _452_/C _452_/A _452_/B vssd1 vssd1 vccd1 vccd1 _471_/C sky130_fd_sc_hd__o211a_4
X_391_ _712_/A _683_/A _723_/A vssd1 vssd1 vccd1 vccd1 _660_/B sky130_fd_sc_hd__nor3_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_727_ _705_/A _754_/D _726_/Y _737_/A vssd1 vssd1 vccd1 vccd1 _767_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_658_ _659_/S _658_/B _658_/C vssd1 vssd1 vccd1 vccd1 _658_/Y sky130_fd_sc_hd__nand3b_1
X_589_ _589_/A _589_/B vssd1 vssd1 vccd1 vccd1 _589_/Y sky130_fd_sc_hd__nor2_2
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtt2_tholin_namebadge_73 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_73/HI io_oeb[26]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_51 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_51/HI io_oeb[4]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_62 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_62/HI io_oeb[15]
+ sky130_fd_sc_hd__conb_1
Xfanout25 _477_/Y vssd1 vssd1 vccd1 vccd1 _748_/D sky130_fd_sc_hd__buf_4
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout36 _767_/Q vssd1 vssd1 vccd1 vccd1 _705_/A sky130_fd_sc_hd__buf_2
Xfanout14 _491_/X vssd1 vssd1 vccd1 vccd1 _547_/A sky130_fd_sc_hd__buf_4
XANTENNA__624__A1 _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_374_ _747_/Q vssd1 vssd1 vccd1 vccd1 _470_/A sky130_fd_sc_hd__inv_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_443_ _453_/A _453_/B _444_/B vssd1 vssd1 vccd1 vccd1 _443_/X sky130_fd_sc_hd__or3_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_512_ _488_/Y _492_/Y _500_/X _511_/X vssd1 vssd1 vccd1 vccd1 _512_/X sky130_fd_sc_hd__a31o_1
XANTENNA__523__A _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_426_ _656_/C _433_/A _426_/C _426_/D vssd1 vssd1 vccd1 vccd1 _426_/X sky130_fd_sc_hd__and4bb_2
Xinput4 rst vssd1 vssd1 vccd1 vccd1 _737_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _769_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_409_ _429_/C _405_/A _426_/D _434_/A vssd1 vssd1 vccd1 vccd1 _664_/B sky130_fd_sc_hd__a211oi_4
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_760_ _762_/CLK _760_/D vssd1 vssd1 vccd1 vccd1 _760_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__681__C1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_691_ _691_/A vssd1 vssd1 vccd1 vccd1 _692_/B sky130_fd_sc_hd__inv_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__497__A2 _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_743_ _758_/CLK _743_/D vssd1 vssd1 vccd1 vccd1 _743_/Q sky130_fd_sc_hd__dfxtp_1
X_674_ _678_/A _439_/A _638_/Y vssd1 vssd1 vccd1 vccd1 _674_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__441__A _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_390_ _385_/X _706_/B _680_/A _390_/D vssd1 vssd1 vccd1 vccd1 _723_/A sky130_fd_sc_hd__nand4b_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_657_ _664_/A _657_/B _657_/C vssd1 vssd1 vccd1 vccd1 _658_/C sky130_fd_sc_hd__or3_1
X_726_ _728_/C _725_/Y _723_/A vssd1 vssd1 vccd1 vccd1 _726_/Y sky130_fd_sc_hd__o21ai_1
X_588_ _616_/B _579_/Y _583_/X _587_/X vssd1 vssd1 vccd1 vccd1 _758_/D sky130_fd_sc_hd__o22a_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout15 _491_/X vssd1 vssd1 vccd1 vccd1 _610_/B sky130_fd_sc_hd__buf_2
Xfanout26 _455_/Y vssd1 vssd1 vccd1 vccd1 _545_/A sky130_fd_sc_hd__buf_4
Xfanout37 _721_/A vssd1 vssd1 vccd1 vccd1 _429_/D sky130_fd_sc_hd__buf_4
Xtt2_tholin_namebadge_63 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_63/HI io_oeb[16]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_52 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_52/HI io_oeb[5]
+ sky130_fd_sc_hd__conb_1
X_511_ _558_/A _508_/Y _510_/X _547_/A _507_/X vssd1 vssd1 vccd1 vccd1 _511_/X sky130_fd_sc_hd__o311a_1
X_373_ _746_/Q vssd1 vssd1 vccd1 vccd1 _441_/B sky130_fd_sc_hd__inv_2
X_442_ _452_/A _452_/B _442_/C vssd1 vssd1 vccd1 vccd1 _493_/B sky130_fd_sc_hd__and3_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__560__A1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_709_ _706_/X _709_/B vssd1 vssd1 vccd1 vccd1 _709_/X sky130_fd_sc_hd__and2b_1
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_425_ _429_/D _655_/A _426_/C _429_/C _429_/B vssd1 vssd1 vccd1 vccd1 _434_/B sky130_fd_sc_hd__o311a_1
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__451__B1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_408_ _656_/A _405_/A _403_/B vssd1 vssd1 vccd1 vccd1 _408_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__444__A _747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_690_ _712_/B _758_/Q vssd1 vssd1 vccd1 vccd1 _691_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_742_ _758_/CLK _742_/D vssd1 vssd1 vccd1 vccd1 _742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__406__A0 _678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_673_ _739_/Q _453_/A _671_/X _672_/X vssd1 vssd1 vccd1 vccd1 _739_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__590__C1 _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_656_ _656_/A _656_/B _656_/C _426_/C vssd1 vssd1 vccd1 vccd1 _657_/C sky130_fd_sc_hd__or4b_1
X_725_ _721_/A _721_/B _705_/A vssd1 vssd1 vccd1 vccd1 _725_/Y sky130_fd_sc_hd__a21oi_1
X_587_ _547_/A _585_/Y _586_/X _752_/D vssd1 vssd1 vccd1 vccd1 _587_/X sky130_fd_sc_hd__a31o_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout27 _455_/Y vssd1 vssd1 vccd1 vccd1 _558_/A sky130_fd_sc_hd__buf_4
Xfanout16 _749_/D vssd1 vssd1 vccd1 vccd1 _618_/A sky130_fd_sc_hd__buf_4
Xfanout38 _766_/Q vssd1 vssd1 vccd1 vccd1 _721_/A sky130_fd_sc_hd__clkbuf_4
Xtt2_tholin_namebadge_64 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_64/HI io_oeb[17]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_53 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_53/HI io_oeb[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_441_ _678_/A _441_/B vssd1 vssd1 vccd1 vccd1 _444_/B sky130_fd_sc_hd__nand2_2
X_510_ _510_/A _552_/B _541_/B _514_/D vssd1 vssd1 vccd1 vccd1 _510_/X sky130_fd_sc_hd__and4_1
X_372_ _678_/A vssd1 vssd1 vccd1 vccd1 _664_/A sky130_fd_sc_hd__inv_2
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_639_ _664_/A _439_/A _435_/B _637_/A vssd1 vssd1 vccd1 vccd1 _639_/X sky130_fd_sc_hd__a22o_1
X_708_ _737_/A _382_/X _707_/Y _754_/D vssd1 vssd1 vccd1 vccd1 _709_/B sky130_fd_sc_hd__a211o_1
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_424_ _439_/A _638_/A vssd1 vssd1 vccd1 vccd1 _424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__515__A2 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__451__A1 _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_407_ _429_/B _429_/C vssd1 vssd1 vccd1 vccd1 _426_/D sky130_fd_sc_hd__and2_4
XANTENNA__506__A2 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__672__A1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_741_ _758_/CLK _741_/D vssd1 vssd1 vccd1 vccd1 _741_/Q sky130_fd_sc_hd__dfxtp_1
X_672_ _430_/A _658_/C _660_/Y _658_/B vssd1 vssd1 vccd1 vccd1 _672_/X sky130_fd_sc_hd__o211a_1
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_724_ _721_/A _754_/D _723_/Y _737_/A vssd1 vssd1 vccd1 vccd1 _766_/D sky130_fd_sc_hd__a22o_1
X_655_ _655_/A _655_/B _655_/C _655_/D vssd1 vssd1 vccd1 vccd1 _658_/B sky130_fd_sc_hd__or4_2
X_586_ _596_/A _545_/B _555_/X _508_/Y _533_/A vssd1 vssd1 vccd1 vccd1 _586_/X sky130_fd_sc_hd__a2111o_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 _765_/Q vssd1 vssd1 vccd1 vccd1 _655_/A sky130_fd_sc_hd__buf_4
Xfanout28 _480_/A vssd1 vssd1 vccd1 vccd1 _493_/C sky130_fd_sc_hd__buf_6
Xfanout17 _749_/D vssd1 vssd1 vccd1 vccd1 _589_/A sky130_fd_sc_hd__clkbuf_4
Xtt2_tholin_namebadge_65 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_65/HI io_oeb[18]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_54 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_54/HI io_oeb[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_371_ _429_/C vssd1 vssd1 vccd1 vccd1 _404_/C sky130_fd_sc_hd__inv_2
X_440_ _664_/A _746_/Q vssd1 vssd1 vccd1 vccd1 _442_/C sky130_fd_sc_hd__nor2_1
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_707_ _744_/Q _745_/Q _712_/A vssd1 vssd1 vccd1 vccd1 _707_/Y sky130_fd_sc_hd__a21oi_1
X_638_ _638_/A _638_/B vssd1 vssd1 vccd1 vccd1 _638_/Y sky130_fd_sc_hd__nand2_1
X_569_ _552_/B _566_/Y _567_/X _558_/A vssd1 vssd1 vccd1 vccd1 _569_/X sky130_fd_sc_hd__a211o_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_423_ _656_/C _426_/D _433_/A vssd1 vssd1 vccd1 vccd1 _638_/A sky130_fd_sc_hd__a21oi_4
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_406_ _678_/B _405_/X _406_/S vssd1 vssd1 vccd1 vccd1 _406_/X sky130_fd_sc_hd__mux2_2
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__471__A _747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_740_ _770_/CLK _740_/D vssd1 vssd1 vccd1 vccd1 _740_/Q sky130_fd_sc_hd__dfxtp_1
X_671_ _683_/A _671_/B _671_/C _671_/D vssd1 vssd1 vccd1 vccd1 _671_/X sky130_fd_sc_hd__or4_1
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__466__A _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_654_ _685_/A _656_/B _712_/B vssd1 vssd1 vccd1 vccd1 _655_/D sky130_fd_sc_hd__a21o_1
X_723_ _723_/A _723_/B vssd1 vssd1 vccd1 vccd1 _723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_585_ _585_/A _585_/B _585_/C vssd1 vssd1 vccd1 vccd1 _585_/Y sky130_fd_sc_hd__nand3_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtt2_tholin_namebadge_55 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_55/HI io_oeb[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_13_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout29 _393_/X vssd1 vssd1 vccd1 vccd1 _453_/A sky130_fd_sc_hd__buf_4
Xfanout18 _481_/Y vssd1 vssd1 vccd1 vccd1 _749_/D sky130_fd_sc_hd__clkbuf_4
Xtt2_tholin_namebadge_66 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_66/HI io_oeb[19]
+ sky130_fd_sc_hd__conb_1
X_370_ _656_/A vssd1 vssd1 vccd1 vccd1 _404_/B sky130_fd_sc_hd__inv_2
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_637_ _637_/A _637_/B vssd1 vssd1 vccd1 vccd1 _637_/Y sky130_fd_sc_hd__nand2_1
X_706_ _737_/A _706_/B _728_/C vssd1 vssd1 vccd1 vccd1 _706_/X sky130_fd_sc_hd__and3_1
X_499_ _551_/A _510_/A _544_/A vssd1 vssd1 vccd1 vccd1 _499_/X sky130_fd_sc_hd__a21o_1
X_568_ _746_/D _544_/A _573_/C _514_/A vssd1 vssd1 vccd1 vccd1 _577_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__463__B1 _747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_422_ _706_/B _405_/A _401_/Y _394_/Y _402_/X vssd1 vssd1 vccd1 vccd1 _439_/B sky130_fd_sc_hd__o221a_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_405_ _405_/A _637_/A vssd1 vssd1 vccd1 vccd1 _405_/X sky130_fd_sc_hd__or2_1
XANTENNA__427__B1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_670_ _448_/X _662_/X _399_/X vssd1 vssd1 vccd1 vccd1 _671_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__557__C1 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_722_ _656_/B _712_/B _405_/A _721_/Y vssd1 vssd1 vccd1 vccd1 _723_/B sky130_fd_sc_hd__a31o_1
X_653_ _712_/B _653_/B _653_/C vssd1 vssd1 vccd1 vccd1 _659_/S sky130_fd_sc_hd__and3_1
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_584_ _584_/A _584_/B vssd1 vssd1 vccd1 vccd1 _585_/C sky130_fd_sc_hd__nand2_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout19 _533_/A vssd1 vssd1 vccd1 vccd1 _585_/A sky130_fd_sc_hd__buf_4
Xtt2_tholin_namebadge_67 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_67/HI io_oeb[20]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_56 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_56/HI io_oeb[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_567_ _462_/A _566_/B _480_/B _480_/A vssd1 vssd1 vccd1 vccd1 _567_/X sky130_fd_sc_hd__o22a_1
X_705_ _705_/A _721_/A _721_/B vssd1 vssd1 vccd1 vccd1 _728_/C sky130_fd_sc_hd__and3_1
X_636_ _759_/Q _755_/Q _762_/Q vssd1 vssd1 vccd1 vccd1 _636_/X sky130_fd_sc_hd__mux2_4
X_498_ _610_/A _748_/D vssd1 vssd1 vccd1 vccd1 _498_/Y sky130_fd_sc_hd__nand2_2
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_421_ _429_/B _655_/A _426_/C _435_/B vssd1 vssd1 vccd1 vccd1 _421_/X sky130_fd_sc_hd__a31o_4
XANTENNA__564__B _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_619_ _530_/A _625_/A _545_/A vssd1 vssd1 vccd1 vccd1 _619_/X sky130_fd_sc_hd__o21a_1
XANTENNA__693__A1 _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output8_A _739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_404_ _434_/A _404_/B _404_/C _405_/A vssd1 vssd1 vccd1 vccd1 _439_/A sky130_fd_sc_hd__and4_4
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_798_ _798_/A vssd1 vssd1 vccd1 vccd1 _798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_721_ _721_/A _721_/B vssd1 vssd1 vccd1 vccd1 _721_/Y sky130_fd_sc_hd__nor2_1
X_583_ _751_/D _583_/B _583_/C vssd1 vssd1 vccd1 vccd1 _583_/X sky130_fd_sc_hd__and3_1
X_652_ _683_/A _652_/B vssd1 vssd1 vccd1 vccd1 _652_/X sky130_fd_sc_hd__or2_1
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__583__A _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__539__B1 _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__493__A _748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtt2_tholin_namebadge_68 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_68/HI io_oeb[21]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_57 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_57/HI io_oeb[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_704_ _704_/A _704_/B vssd1 vssd1 vccd1 vccd1 _721_/B sky130_fd_sc_hd__nor2_2
X_635_ _634_/A _633_/A _633_/B vssd1 vssd1 vccd1 vccd1 _743_/D sky130_fd_sc_hd__a21bo_1
X_566_ _584_/A _566_/B vssd1 vssd1 vccd1 vccd1 _566_/Y sky130_fd_sc_hd__xnor2_1
X_497_ _584_/A _748_/D _480_/B _493_/C vssd1 vssd1 vccd1 vccd1 _625_/B sky130_fd_sc_hd__o22a_4
XFILLER_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_420_ _656_/A _429_/D _429_/C _433_/A vssd1 vssd1 vccd1 vccd1 _435_/B sky130_fd_sc_hd__a211o_4
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ _474_/Y _566_/B _558_/B vssd1 vssd1 vccd1 vccd1 _549_/X sky130_fd_sc_hd__o21a_1
X_618_ _618_/A _618_/B _618_/C vssd1 vssd1 vccd1 vccd1 _618_/X sky130_fd_sc_hd__or3_1
XANTENNA__669__C1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_403_ _656_/A _403_/B _433_/A vssd1 vssd1 vccd1 vccd1 _637_/A sky130_fd_sc_hd__or3b_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__409__A2 _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _762_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__557__A1 _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_720_ _765_/Q _754_/D _719_/Y _737_/A vssd1 vssd1 vccd1 vccd1 _765_/D sky130_fd_sc_hd__a22o_1
X_651_ _406_/S _642_/X _649_/X _650_/X vssd1 vssd1 vccd1 vccd1 _652_/B sky130_fd_sc_hd__a31o_1
X_582_ _462_/A _558_/B _514_/X _585_/A vssd1 vssd1 vccd1 vccd1 _583_/C sky130_fd_sc_hd__a211o_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__539__A1 _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtt2_tholin_namebadge_69 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_69/HI io_oeb[22]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_47 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_47/HI io_oeb[0]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_58 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_58/HI io_oeb[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__702__A1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_634_ _634_/A _634_/B vssd1 vssd1 vccd1 vccd1 _742_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_703_ _660_/Y _700_/X _702_/X _453_/A _741_/Q vssd1 vssd1 vccd1 vccd1 _741_/D sky130_fd_sc_hd__a32o_1
X_496_ _552_/B _589_/B _514_/D _585_/A vssd1 vssd1 vccd1 vccd1 _496_/X sky130_fd_sc_hd__a31o_1
X_565_ _610_/A _618_/A _585_/B vssd1 vssd1 vccd1 vccd1 _565_/X sky130_fd_sc_hd__and3_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_617_ _752_/D _609_/Y _610_/X _616_/X vssd1 vssd1 vccd1 vccd1 _760_/D sky130_fd_sc_hd__a31o_1
X_548_ _547_/A _538_/X _542_/Y _547_/Y vssd1 vssd1 vccd1 vccd1 _756_/D sky130_fd_sc_hd__a22oi_2
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_479_ _749_/Q _489_/D vssd1 vssd1 vccd1 vccd1 _480_/B sky130_fd_sc_hd__xnor2_4
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_402_ _429_/B _429_/C _434_/A vssd1 vssd1 vccd1 vccd1 _402_/X sky130_fd_sc_hd__o21a_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__752__D _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_650_ _448_/X _636_/X _399_/X vssd1 vssd1 vccd1 vccd1 _650_/X sky130_fd_sc_hd__o21a_1
X_581_ _618_/A _552_/C _580_/Y _558_/A vssd1 vssd1 vccd1 vccd1 _583_/B sky130_fd_sc_hd__a211o_1
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtt2_tholin_namebadge_48 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_48/HI io_oeb[1]
+ sky130_fd_sc_hd__conb_1
Xtt2_tholin_namebadge_59 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_59/HI io_oeb[12]
+ sky130_fd_sc_hd__conb_1
X_633_ _633_/A _633_/B vssd1 vssd1 vccd1 vccd1 _634_/B sky130_fd_sc_hd__nand2_1
X_702_ _430_/A _658_/Y _714_/B _686_/X vssd1 vssd1 vccd1 vccd1 _702_/X sky130_fd_sc_hd__a31o_1
X_495_ _564_/A _495_/B _495_/C vssd1 vssd1 vccd1 vccd1 _514_/D sky130_fd_sc_hd__or3_4
X_564_ _564_/A _584_/A vssd1 vssd1 vccd1 vccd1 _585_/B sky130_fd_sc_hd__nand2_2
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__687__A1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_616_ _615_/X _616_/B _616_/C vssd1 vssd1 vccd1 vccd1 _616_/X sky130_fd_sc_hd__and3b_1
X_547_ _547_/A _547_/B vssd1 vssd1 vccd1 vccd1 _547_/Y sky130_fd_sc_hd__nor2_1
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_478_ _749_/Q _489_/D vssd1 vssd1 vccd1 vccd1 _573_/C sky130_fd_sc_hd__xor2_4
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__602__A1 _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_401_ _429_/C _429_/B _434_/A vssd1 vssd1 vccd1 vccd1 _401_/Y sky130_fd_sc_hd__nand3b_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__587__B1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output6_A _753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__732__S _769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_580_ _589_/B _499_/X _618_/A vssd1 vssd1 vccd1 vccd1 _580_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtt2_tholin_namebadge_49 vssd1 vssd1 vccd1 vccd1 tt2_tholin_namebadge_49/HI io_oeb[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_632_ _632_/A _632_/B vssd1 vssd1 vccd1 vccd1 _633_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_563_ _618_/A _530_/B _558_/C _558_/A vssd1 vssd1 vccd1 vccd1 _563_/X sky130_fd_sc_hd__a211o_1
X_701_ _390_/D _704_/B vssd1 vssd1 vccd1 vccd1 _714_/B sky130_fd_sc_hd__nand2b_1
X_494_ _748_/Q _610_/A vssd1 vssd1 vccd1 vccd1 _589_/B sky130_fd_sc_hd__or2_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_615_ _545_/A _589_/Y _597_/A _614_/X _610_/B vssd1 vssd1 vccd1 vccd1 _615_/X sky130_fd_sc_hd__o311a_1
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_546_ _530_/X _610_/C _543_/X _752_/D vssd1 vssd1 vccd1 vccd1 _547_/B sky130_fd_sc_hd__o211a_1
X_477_ _544_/A vssd1 vssd1 vccd1 vccd1 _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_400_ _721_/A _655_/A _426_/C vssd1 vssd1 vccd1 vccd1 _405_/A sky130_fd_sc_hd__and3_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_529_ _512_/X _528_/X _752_/D vssd1 vssd1 vccd1 vccd1 _755_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_700_ _680_/A _699_/X _698_/X _683_/A vssd1 vssd1 vccd1 vccd1 _700_/X sky130_fd_sc_hd__a211o_1
X_631_ _632_/A _632_/B vssd1 vssd1 vccd1 vccd1 _633_/A sky130_fd_sc_hd__or2_1
X_493_ _748_/Q _493_/B _493_/C _493_/D vssd1 vssd1 vccd1 vccd1 _541_/B sky130_fd_sc_hd__or4_4
X_562_ _577_/B _625_/B _561_/X _625_/A _585_/A vssd1 vssd1 vccd1 vccd1 _562_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__605__B1 _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_545_ _545_/A _545_/B vssd1 vssd1 vccd1 vccd1 _610_/C sky130_fd_sc_hd__or2_2
X_614_ _552_/A _545_/B _536_/A vssd1 vssd1 vccd1 vccd1 _614_/X sky130_fd_sc_hd__a21o_1
X_476_ _489_/D _475_/X _493_/C vssd1 vssd1 vccd1 vccd1 _544_/A sky130_fd_sc_hd__a21o_4
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_459_ _444_/B _453_/C _453_/A _453_/B vssd1 vssd1 vccd1 vccd1 _470_/C sky130_fd_sc_hd__a211o_1
X_528_ _513_/X _517_/X _527_/X _547_/A vssd1 vssd1 vccd1 vccd1 _528_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__699__A1 _678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_630_ _623_/X _629_/Y _752_/D vssd1 vssd1 vccd1 vccd1 _761_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_492_ _610_/B vssd1 vssd1 vccd1 vccd1 _492_/Y sky130_fd_sc_hd__inv_2
X_561_ _520_/A _566_/B _573_/C _514_/A vssd1 vssd1 vccd1 vccd1 _561_/X sky130_fd_sc_hd__o211a_2
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_759_ _769_/CLK _759_/D vssd1 vssd1 vccd1 vccd1 _759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_613_ _611_/X _612_/X _610_/B vssd1 vssd1 vccd1 vccd1 _616_/C sky130_fd_sc_hd__a21o_1
X_475_ _452_/A _452_/B _445_/C _564_/A vssd1 vssd1 vccd1 vccd1 _475_/X sky130_fd_sc_hd__a31o_2
X_544_ _544_/A _573_/C vssd1 vssd1 vccd1 vccd1 _545_/B sky130_fd_sc_hd__nor2_2
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_527_ _521_/X _522_/X _525_/X _526_/X vssd1 vssd1 vccd1 vccd1 _527_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_458_ _678_/A _452_/A _452_/B _441_/B vssd1 vssd1 vccd1 vccd1 _470_/B sky130_fd_sc_hd__a31o_2
X_389_ _684_/A _712_/B vssd1 vssd1 vccd1 vccd1 _390_/D sky130_fd_sc_hd__nor2_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_560_ _751_/D _554_/X _559_/X _752_/D vssd1 vssd1 vccd1 vccd1 _560_/X sky130_fd_sc_hd__a211o_1
X_491_ _514_/A _501_/B _491_/C vssd1 vssd1 vccd1 vccd1 _491_/X sky130_fd_sc_hd__and3_1
X_758_ _758_/CLK _758_/D vssd1 vssd1 vccd1 vccd1 _758_/Q sky130_fd_sc_hd__dfxtp_1
X_689_ _638_/A _637_/Y _433_/Y vssd1 vssd1 vccd1 vccd1 _689_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_612_ _530_/A _625_/A _558_/B _610_/A _545_/A vssd1 vssd1 vccd1 vccd1 _612_/X sky130_fd_sc_hd__a221o_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__675__S _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_543_ _514_/D _504_/X _530_/C _589_/A _585_/A vssd1 vssd1 vccd1 vccd1 _543_/X sky130_fd_sc_hd__a221o_1
X_474_ _474_/A _596_/A vssd1 vssd1 vccd1 vccd1 _474_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__599__A1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__524__A _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__450__B1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_526_ _618_/A _541_/B _530_/C _558_/A vssd1 vssd1 vccd1 vccd1 _526_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_457_ _664_/A _453_/A _453_/B _746_/Q vssd1 vssd1 vccd1 vccd1 _493_/D sky130_fd_sc_hd__o31a_4
X_388_ _744_/Q _745_/Q vssd1 vssd1 vccd1 vccd1 _406_/S sky130_fd_sc_hd__nand2b_4
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__510__C _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__404__D _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_509_ _596_/A _589_/A vssd1 vssd1 vccd1 vccd1 _509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__712__A _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_490_ _455_/A _751_/Q vssd1 vssd1 vccd1 vccd1 _491_/C sky130_fd_sc_hd__nand2b_1
Xclkbuf_2_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _758_/CLK sky130_fd_sc_hd__clkbuf_16
X_688_ _660_/Y _683_/X _687_/X _453_/A _740_/Q vssd1 vssd1 vccd1 vccd1 _740_/D sky130_fd_sc_hd__a32o_1
X_757_ _762_/CLK _757_/D vssd1 vssd1 vccd1 vccd1 _757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_542_ _625_/B _541_/Y _540_/X _616_/B vssd1 vssd1 vccd1 vccd1 _542_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_473_ _495_/C _495_/B _470_/C _470_/B vssd1 vssd1 vccd1 vccd1 _510_/A sky130_fd_sc_hd__a2bb2o_4
X_611_ _510_/A _618_/A _596_/B _561_/X _536_/A vssd1 vssd1 vccd1 vccd1 _611_/X sky130_fd_sc_hd__a2111o_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_456_ _545_/A vssd1 vssd1 vccd1 vccd1 _536_/A sky130_fd_sc_hd__inv_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_525_ _510_/A _566_/B _552_/B _551_/A vssd1 vssd1 vccd1 vccd1 _525_/X sky130_fd_sc_hd__o211a_1
XANTENNA__450__A1 _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_387_ _744_/Q _745_/Q vssd1 vssd1 vccd1 vccd1 _680_/A sky130_fd_sc_hd__and2b_4
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ _439_/A _439_/B vssd1 vssd1 vccd1 vccd1 _637_/B sky130_fd_sc_hd__nor2_1
X_508_ _552_/B _589_/B vssd1 vssd1 vccd1 vccd1 _508_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__617__A1 _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__608__B2 _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout31_A _769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_756_ _758_/CLK _756_/D vssd1 vssd1 vccd1 vccd1 _756_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output12_A _798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_687_ _430_/A _658_/Y _685_/Y _686_/X vssd1 vssd1 vccd1 vccd1 _687_/X sky130_fd_sc_hd__a31o_1
X_610_ _610_/A _610_/B _610_/C vssd1 vssd1 vccd1 vccd1 _610_/X sky130_fd_sc_hd__or3_1
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_541_ _750_/D _541_/B vssd1 vssd1 vccd1 vccd1 _541_/Y sky130_fd_sc_hd__nand2_1
X_472_ _493_/D _471_/C _495_/B _495_/C vssd1 vssd1 vccd1 vccd1 _596_/A sky130_fd_sc_hd__o22a_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_739_ _762_/CLK _739_/D vssd1 vssd1 vccd1 vccd1 _739_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_386_ _769_/Q _403_/B vssd1 vssd1 vccd1 vccd1 _706_/B sky130_fd_sc_hd__and2_2
X_524_ _610_/A _544_/A vssd1 vssd1 vccd1 vccd1 _524_/Y sky130_fd_sc_hd__nand2_1
X_455_ _455_/A _493_/C _455_/C vssd1 vssd1 vccd1 vccd1 _455_/Y sky130_fd_sc_hd__nor3_2
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_438_ _406_/X _419_/X _427_/Y _436_/X _712_/A vssd1 vssd1 vccd1 vccd1 _452_/B sky130_fd_sc_hd__a41o_4
X_369_ _754_/Q vssd1 vssd1 vccd1 vccd1 _712_/A sky130_fd_sc_hd__inv_6
X_507_ _498_/Y _504_/X _506_/X _585_/A vssd1 vssd1 vccd1 vccd1 _507_/X sky130_fd_sc_hd__a211o_1
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout24_A _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_755_ _762_/CLK _755_/D vssd1 vssd1 vccd1 vccd1 _755_/Q sky130_fd_sc_hd__dfxtp_1
X_686_ _656_/B _412_/Y _659_/S _382_/X vssd1 vssd1 vccd1 vccd1 _686_/X sky130_fd_sc_hd__a31o_1
XANTENNA__535__B2 _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_540_ _747_/D _530_/A _541_/B _539_/X vssd1 vssd1 vccd1 vccd1 _540_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_471_ _747_/Q _493_/D _471_/C vssd1 vssd1 vccd1 vccd1 _551_/A sky130_fd_sc_hd__or3_4
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_738_ _758_/CLK _738_/D vssd1 vssd1 vccd1 vccd1 _798_/A sky130_fd_sc_hd__dfxtp_2
X_669_ _637_/Y _662_/X _668_/X _430_/A vssd1 vssd1 vccd1 vccd1 _671_/C sky130_fd_sc_hd__o211a_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__374__A _747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_523_ _610_/A _544_/A vssd1 vssd1 vccd1 vccd1 _618_/C sky130_fd_sc_hd__and2_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_385_ _705_/A _721_/A _765_/Q _685_/A vssd1 vssd1 vccd1 vccd1 _385_/X sky130_fd_sc_hd__or4_1
X_454_ _749_/Q _489_/D _750_/Q vssd1 vssd1 vccd1 vccd1 _455_/C sky130_fd_sc_hd__o21a_1
XANTENNA__729__A1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_506_ _493_/C _480_/B _577_/B _551_/A vssd1 vssd1 vccd1 vccd1 _506_/X sky130_fd_sc_hd__o211a_1
X_437_ _406_/X _419_/X _427_/Y _436_/X _712_/A vssd1 vssd1 vccd1 vccd1 _453_/B sky130_fd_sc_hd__a41oi_4
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__647__B1 _430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__553__A2 _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout17_A _749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_685_ _685_/A _704_/B vssd1 vssd1 vccd1 vccd1 _685_/Y sky130_fd_sc_hd__xnor2_1
X_754_ _770_/CLK _754_/D vssd1 vssd1 vccd1 vccd1 _754_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__535__A2 _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__526__A2 _541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__660__A _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_470_ _470_/A _470_/B _470_/C vssd1 vssd1 vccd1 vccd1 _474_/A sky130_fd_sc_hd__and3_1
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_668_ _435_/B _638_/Y _667_/X _662_/X _428_/Y vssd1 vssd1 vccd1 vccd1 _668_/X sky130_fd_sc_hd__a32o_1
X_737_ _737_/A _737_/B vssd1 vssd1 vccd1 vccd1 _753_/D sky130_fd_sc_hd__nor2_1
X_599_ _751_/D _595_/Y _598_/X _593_/Y vssd1 vssd1 vccd1 vccd1 _599_/X sky130_fd_sc_hd__a31o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_453_ _453_/A _453_/B _453_/C vssd1 vssd1 vccd1 vccd1 _514_/A sky130_fd_sc_hd__or3_4
X_522_ _499_/X _504_/X _585_/A vssd1 vssd1 vccd1 vccd1 _522_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__565__A _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_384_ _705_/A _685_/A _656_/C vssd1 vssd1 vccd1 vccd1 _653_/C sky130_fd_sc_hd__nor3_1
XANTENNA__674__A1 _678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_436_ _692_/A _435_/X _430_/Y vssd1 vssd1 vccd1 vccd1 _436_/X sky130_fd_sc_hd__a21o_2
X_505_ _498_/Y _504_/X _533_/A vssd1 vssd1 vccd1 vccd1 _505_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__629__A1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_419_ _664_/B _418_/B _418_/X _382_/X vssd1 vssd1 vccd1 vccd1 _419_/X sky130_fd_sc_hd__o211a_4
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_770_ _770_/CLK _770_/D vssd1 vssd1 vccd1 vccd1 _770_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__573__A _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__467__B _746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_753_ _769_/CLK _753_/D vssd1 vssd1 vccd1 vccd1 _753_/Q sky130_fd_sc_hd__dfxtp_1
X_684_ _684_/A _712_/B vssd1 vssd1 vccd1 vccd1 _704_/B sky130_fd_sc_hd__nand2_2
XFILLER_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_736_ _382_/X _660_/Y _735_/X _453_/A _770_/Q vssd1 vssd1 vccd1 vccd1 _770_/D sky130_fd_sc_hd__a32o_1
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output10_A _741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_667_ _678_/A _405_/A _637_/A vssd1 vssd1 vccd1 vccd1 _667_/X sky130_fd_sc_hd__a21o_1
X_598_ _573_/C _484_/Y _597_/A _750_/D vssd1 vssd1 vccd1 vccd1 _598_/X sky130_fd_sc_hd__a211o_1
XANTENNA__480__B _480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__601__C1 _751_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_383_ _655_/A _426_/C vssd1 vssd1 vccd1 vccd1 _383_/X sky130_fd_sc_hd__or2_1
X_452_ _452_/A _452_/B _452_/C vssd1 vssd1 vccd1 vccd1 _480_/A sky130_fd_sc_hd__and3_4
X_521_ _552_/C _618_/B _610_/A _480_/B vssd1 vssd1 vccd1 vccd1 _521_/X sky130_fd_sc_hd__o211a_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_719_ _721_/B _718_/Y _723_/A vssd1 vssd1 vccd1 vccd1 _719_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__408__A2 _405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_435_ _680_/A _435_/B vssd1 vssd1 vccd1 vccd1 _435_/X sky130_fd_sc_hd__or2_1
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_504_ _474_/A _596_/A _566_/B _573_/C _514_/A vssd1 vssd1 vccd1 vccd1 _504_/X sky130_fd_sc_hd__o311a_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__486__A _747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__574__A1 _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_418_ _657_/B _418_/B _418_/C _417_/C vssd1 vssd1 vccd1 vccd1 _418_/X sky130_fd_sc_hd__or4b_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__573__B _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_752_ _758_/CLK _752_/D vssd1 vssd1 vccd1 vccd1 _752_/Q sky130_fd_sc_hd__dfxtp_1
X_683_ _683_/A _683_/B _683_/C vssd1 vssd1 vccd1 vccd1 _683_/X sky130_fd_sc_hd__or3_1
XANTENNA__584__A _584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__494__A _748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__438__B1 _712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_735_ _406_/S _733_/X _734_/Y _399_/X _449_/Y vssd1 vssd1 vccd1 vccd1 _735_/X sky130_fd_sc_hd__a32o_1
X_666_ _410_/Y _662_/X _665_/X _412_/Y _406_/S vssd1 vssd1 vccd1 vccd1 _671_/B sky130_fd_sc_hd__o2111a_1
X_597_ _597_/A vssd1 vssd1 vccd1 vccd1 _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__399__A _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__390__C _680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_520_ _520_/A _566_/B vssd1 vssd1 vccd1 vccd1 _530_/C sky130_fd_sc_hd__nand2_2
X_382_ _429_/B _657_/B _382_/C vssd1 vssd1 vccd1 vccd1 _382_/X sky130_fd_sc_hd__or3_4
X_451_ _680_/A _448_/X _712_/A vssd1 vssd1 vccd1 vccd1 _452_/C sky130_fd_sc_hd__a21o_2
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_649_ _636_/X _648_/Y _647_/X _646_/X vssd1 vssd1 vccd1 vccd1 _649_/X sky130_fd_sc_hd__a211o_1
X_718_ _685_/A _684_/A _712_/B _765_/Q vssd1 vssd1 vccd1 vccd1 _718_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_503_ _752_/D vssd1 vssd1 vccd1 vccd1 _616_/B sky130_fd_sc_hd__inv_2
X_434_ _434_/A _434_/B _638_/B vssd1 vssd1 vccd1 vccd1 _692_/A sky130_fd_sc_hd__or3b_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_417_ _656_/A _656_/C _417_/C vssd1 vssd1 vccd1 vccd1 _648_/B sky130_fd_sc_hd__and3_4
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_751_ _758_/CLK _751_/D vssd1 vssd1 vccd1 vccd1 _751_/Q sky130_fd_sc_hd__dfxtp_1
X_682_ _412_/Y _677_/X _681_/X _406_/S vssd1 vssd1 vccd1 vccd1 _683_/C sky130_fd_sc_hd__o211a_1
XANTENNA__750__D _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__494__B _610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_734_ _657_/B _648_/B _664_/C _404_/C _412_/Y vssd1 vssd1 vccd1 vccd1 _734_/Y sky130_fd_sc_hd__o221ai_4
X_665_ _648_/Y _662_/X _664_/X _657_/B vssd1 vssd1 vccd1 vccd1 _665_/X sky130_fd_sc_hd__a22o_1
XANTENNA__595__A _750_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_596_ _596_/A _596_/B vssd1 vssd1 vccd1 vccd1 _597_/A sky130_fd_sc_hd__and2_2
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__399__B _678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_381_ _382_/C _404_/B _653_/B vssd1 vssd1 vccd1 vccd1 _683_/A sky130_fd_sc_hd__and3b_4
X_450_ _680_/A _448_/X _712_/A vssd1 vssd1 vccd1 vccd1 _453_/C sky130_fd_sc_hd__a21oi_1
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput5 _770_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_4
X_648_ _657_/B _648_/B vssd1 vssd1 vccd1 vccd1 _648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_717_ _685_/A _754_/D _716_/X _737_/A vssd1 vssd1 vccd1 vccd1 _764_/D sky130_fd_sc_hd__a22o_1
XANTENNA__529__S _752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_579_ _751_/D _575_/Y _578_/X vssd1 vssd1 vccd1 vccd1 _579_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _433_/A _638_/B vssd1 vssd1 vccd1 vccd1 _433_/Y sky130_fd_sc_hd__nor2_1
X_502_ _752_/Q _501_/B _501_/Y _493_/C vssd1 vssd1 vccd1 vccd1 _752_/D sky130_fd_sc_hd__a211o_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_416_ _721_/A _655_/A _656_/A vssd1 vssd1 vccd1 vccd1 _418_/C sky130_fd_sc_hd__o21ai_1
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__748__D _748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_750_ _758_/CLK _750_/D vssd1 vssd1 vccd1 vccd1 _750_/Q sky130_fd_sc_hd__dfxtp_1
X_681_ _653_/B _648_/B _675_/X _664_/B _430_/A vssd1 vssd1 vccd1 vccd1 _681_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_733_ _435_/B _689_/Y _430_/Y vssd1 vssd1 vccd1 vccd1 _733_/X sky130_fd_sc_hd__a21o_1
X_664_ _664_/A _664_/B _664_/C vssd1 vssd1 vccd1 vccd1 _664_/X sky130_fd_sc_hd__or3_1
X_595_ _750_/D _595_/B vssd1 vssd1 vccd1 vccd1 _595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_380_ _426_/C _656_/B _429_/D _655_/A vssd1 vssd1 vccd1 vccd1 _382_/C sky130_fd_sc_hd__a211o_1
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput6 _753_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_4
X_716_ _653_/C _706_/B _680_/A _390_/D _685_/Y vssd1 vssd1 vccd1 vccd1 _716_/X sky130_fd_sc_hd__a41o_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_647_ _664_/A _653_/B _648_/B _430_/A vssd1 vssd1 vccd1 vccd1 _647_/X sky130_fd_sc_hd__a31o_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_578_ _558_/A _576_/X _577_/X _547_/A vssd1 vssd1 vccd1 vccd1 _578_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

