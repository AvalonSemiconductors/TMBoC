VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_MC14500
  CLASS BLOCK ;
  FOREIGN wrapped_MC14500 ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 90.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 86.000 15.090 90.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 8.880 60.000 9.480 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 26.560 60.000 27.160 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 44.240 60.000 44.840 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 61.920 60.000 62.520 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 79.600 60.000 80.200 ;
    END
  END io_in[4]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_out[8]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 86.000 44.990 90.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 79.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.910 10.640 18.510 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.100 10.640 30.700 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.290 10.640 42.890 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.480 10.640 55.080 79.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 78.965 ;
      LAYER met1 ;
        RECT 2.830 10.640 56.970 79.120 ;
      LAYER met2 ;
        RECT 2.860 85.720 14.530 86.770 ;
        RECT 15.370 85.720 44.430 86.770 ;
        RECT 45.270 85.720 56.940 86.770 ;
        RECT 2.860 4.280 56.940 85.720 ;
        RECT 3.410 4.000 8.550 4.280 ;
        RECT 9.390 4.000 14.530 4.280 ;
        RECT 15.370 4.000 20.510 4.280 ;
        RECT 21.350 4.000 26.490 4.280 ;
        RECT 27.330 4.000 32.470 4.280 ;
        RECT 33.310 4.000 38.450 4.280 ;
        RECT 39.290 4.000 44.430 4.280 ;
        RECT 45.270 4.000 50.410 4.280 ;
        RECT 51.250 4.000 56.390 4.280 ;
      LAYER met3 ;
        RECT 10.825 79.200 55.600 80.065 ;
        RECT 10.825 62.920 56.730 79.200 ;
        RECT 10.825 61.520 55.600 62.920 ;
        RECT 10.825 45.240 56.730 61.520 ;
        RECT 10.825 43.840 55.600 45.240 ;
        RECT 10.825 27.560 56.730 43.840 ;
        RECT 10.825 26.160 55.600 27.560 ;
        RECT 10.825 9.880 56.730 26.160 ;
        RECT 10.825 9.015 55.600 9.880 ;
  END
END wrapped_MC14500
END LIBRARY

