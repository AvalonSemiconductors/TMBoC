magic
tech sky130B
magscale 1 2
timestamp 1687097464
<< viali >>
rect 11069 61353 11103 61387
rect 18061 61353 18095 61387
rect 33425 61353 33459 61387
rect 47961 61353 47995 61387
rect 51457 61353 51491 61387
rect 40233 61285 40267 61319
rect 44557 61285 44591 61319
rect 48789 61285 48823 61319
rect 2237 61217 2271 61251
rect 3065 61217 3099 61251
rect 21465 61217 21499 61251
rect 25513 61217 25547 61251
rect 32689 61217 32723 61251
rect 52285 61217 52319 61251
rect 56793 61217 56827 61251
rect 1685 61149 1719 61183
rect 2789 61149 2823 61183
rect 4721 61149 4755 61183
rect 5641 61149 5675 61183
rect 6653 61149 6687 61183
rect 7573 61149 7607 61183
rect 9229 61149 9263 61183
rect 10241 61149 10275 61183
rect 10977 61149 11011 61183
rect 12081 61149 12115 61183
rect 12817 61149 12851 61183
rect 14933 61149 14967 61183
rect 16129 61149 16163 61183
rect 17141 61149 17175 61183
rect 17969 61149 18003 61183
rect 18705 61149 18739 61183
rect 19809 61149 19843 61183
rect 20545 61149 20579 61183
rect 21281 61149 21315 61183
rect 22385 61149 22419 61183
rect 23857 61149 23891 61183
rect 25237 61149 25271 61183
rect 26249 61149 26283 61183
rect 27261 61149 27295 61183
rect 28181 61149 28215 61183
rect 29837 61149 29871 61183
rect 31217 61149 31251 61183
rect 32413 61149 32447 61183
rect 33333 61149 33367 61183
rect 34069 61149 34103 61183
rect 34989 61149 35023 61183
rect 36461 61149 36495 61183
rect 37565 61149 37599 61183
rect 38301 61149 38335 61183
rect 38945 61149 38979 61183
rect 40049 61149 40083 61183
rect 40877 61149 40911 61183
rect 41613 61149 41647 61183
rect 42625 61149 42659 61183
rect 43545 61149 43579 61183
rect 44373 61149 44407 61183
rect 45293 61149 45327 61183
rect 46029 61149 46063 61183
rect 46765 61149 46799 61183
rect 47869 61149 47903 61183
rect 48605 61149 48639 61183
rect 49341 61149 49375 61183
rect 50445 61149 50479 61183
rect 51365 61149 51399 61183
rect 52101 61149 52135 61183
rect 53205 61149 53239 61183
rect 54125 61149 54159 61183
rect 55505 61149 55539 61183
rect 56517 61149 56551 61183
rect 58173 61149 58207 61183
rect 4905 61081 4939 61115
rect 6929 61081 6963 61115
rect 7849 61081 7883 61115
rect 15209 61081 15243 61115
rect 16313 61081 16347 61115
rect 19993 61081 20027 61115
rect 26433 61081 26467 61115
rect 28457 61081 28491 61115
rect 31585 61081 31619 61115
rect 35725 61081 35759 61115
rect 38485 61081 38519 61115
rect 42901 61081 42935 61115
rect 49525 61081 49559 61115
rect 53481 61081 53515 61115
rect 55781 61081 55815 61115
rect 58357 61081 58391 61115
rect 5733 61013 5767 61047
rect 9321 61013 9355 61047
rect 10333 61013 10367 61047
rect 12173 61013 12207 61047
rect 12909 61013 12943 61047
rect 17325 61013 17359 61047
rect 18797 61013 18831 61047
rect 20637 61013 20671 61047
rect 22477 61013 22511 61047
rect 23949 61013 23983 61047
rect 27353 61013 27387 61047
rect 29929 61013 29963 61047
rect 34161 61013 34195 61047
rect 35081 61013 35115 61047
rect 35817 61013 35851 61047
rect 36553 61013 36587 61047
rect 37657 61013 37691 61047
rect 39129 61013 39163 61047
rect 40969 61013 41003 61047
rect 41705 61013 41739 61047
rect 43729 61013 43763 61047
rect 45385 61013 45419 61047
rect 46121 61013 46155 61047
rect 46857 61013 46891 61047
rect 50537 61013 50571 61047
rect 54309 61013 54343 61047
rect 3985 60741 4019 60775
rect 5457 60741 5491 60775
rect 8401 60741 8435 60775
rect 9873 60741 9907 60775
rect 13553 60741 13587 60775
rect 14289 60741 14323 60775
rect 15761 60741 15795 60775
rect 19441 60741 19475 60775
rect 23305 60741 23339 60775
rect 24593 60741 24627 60775
rect 27537 60741 27571 60775
rect 29009 60741 29043 60775
rect 30481 60741 30515 60775
rect 36369 60741 36403 60775
rect 41521 60741 41555 60775
rect 46673 60741 46707 60775
rect 50353 60741 50387 60775
rect 53021 60741 53055 60775
rect 1593 60673 1627 60707
rect 3157 60673 3191 60707
rect 14473 60673 14507 60707
rect 22109 60673 22143 60707
rect 54677 60673 54711 60707
rect 55413 60673 55447 60707
rect 56149 60673 56183 60707
rect 56885 60673 56919 60707
rect 58081 60673 58115 60707
rect 1869 60605 1903 60639
rect 8585 60605 8619 60639
rect 13737 60605 13771 60639
rect 22661 60605 22695 60639
rect 4169 60537 4203 60571
rect 5641 60537 5675 60571
rect 19625 60537 19659 60571
rect 23489 60537 23523 60571
rect 58265 60537 58299 60571
rect 3341 60469 3375 60503
rect 9965 60469 9999 60503
rect 15853 60469 15887 60503
rect 24685 60469 24719 60503
rect 27629 60469 27663 60503
rect 29101 60469 29135 60503
rect 30573 60469 30607 60503
rect 36461 60469 36495 60503
rect 41613 60469 41647 60503
rect 46765 60469 46799 60503
rect 50445 60469 50479 60503
rect 53113 60469 53147 60503
rect 54861 60469 54895 60503
rect 55597 60469 55631 60503
rect 56333 60469 56367 60503
rect 57069 60469 57103 60503
rect 6561 60197 6595 60231
rect 20545 60197 20579 60231
rect 27445 60197 27479 60231
rect 18061 60129 18095 60163
rect 33609 60129 33643 60163
rect 41705 60129 41739 60163
rect 41889 60129 41923 60163
rect 43545 60129 43579 60163
rect 57437 60129 57471 60163
rect 2605 60061 2639 60095
rect 6009 60061 6043 60095
rect 6285 60061 6319 60095
rect 6429 60061 6463 60095
rect 18245 60061 18279 60095
rect 18613 60061 18647 60095
rect 18797 60061 18831 60095
rect 19993 60061 20027 60095
rect 20269 60061 20303 60095
rect 20413 60061 20447 60095
rect 21189 60061 21223 60095
rect 22293 60061 22327 60095
rect 22666 60061 22700 60095
rect 23397 60061 23431 60095
rect 23817 60061 23851 60095
rect 23966 60061 24000 60095
rect 24685 60061 24719 60095
rect 25145 60061 25179 60095
rect 25237 60061 25271 60095
rect 25513 60061 25547 60095
rect 25789 60061 25823 60095
rect 25973 60061 26007 60095
rect 26801 60061 26835 60095
rect 26894 60061 26928 60095
rect 27169 60061 27203 60095
rect 27266 60061 27300 60095
rect 27997 60061 28031 60095
rect 28090 60061 28124 60095
rect 28373 60061 28407 60095
rect 28462 60061 28496 60095
rect 29193 60061 29227 60095
rect 29745 60061 29779 60095
rect 29838 60061 29872 60095
rect 30210 60061 30244 60095
rect 33793 60061 33827 60095
rect 34161 60061 34195 60095
rect 34345 60061 34379 60095
rect 41613 60061 41647 60095
rect 41981 60061 42015 60095
rect 43085 60061 43119 60095
rect 43269 60061 43303 60095
rect 43637 60061 43671 60095
rect 56517 60061 56551 60095
rect 57253 60061 57287 60095
rect 57989 60061 58023 60095
rect 1685 59993 1719 60027
rect 2053 59993 2087 60027
rect 6193 59993 6227 60027
rect 20177 59993 20211 60027
rect 21557 59993 21591 60027
rect 22477 59993 22511 60027
rect 22569 59993 22603 60027
rect 22862 59993 22896 60027
rect 23581 59993 23615 60027
rect 23673 59993 23707 60027
rect 27077 59993 27111 60027
rect 28273 59993 28307 60027
rect 30021 59993 30055 60027
rect 30113 59993 30147 60027
rect 42625 59993 42659 60027
rect 58357 59993 58391 60027
rect 2697 59925 2731 59959
rect 17693 59925 17727 59959
rect 26433 59925 26467 59959
rect 28641 59925 28675 59959
rect 30389 59925 30423 59959
rect 30665 59925 30699 59959
rect 32873 59925 32907 59959
rect 33241 59925 33275 59959
rect 34897 59925 34931 59959
rect 41061 59925 41095 59959
rect 56609 59925 56643 59959
rect 24869 59721 24903 59755
rect 57437 59721 57471 59755
rect 58265 59721 58299 59755
rect 2421 59653 2455 59687
rect 6745 59653 6779 59687
rect 19073 59653 19107 59687
rect 24593 59653 24627 59687
rect 25881 59653 25915 59687
rect 57345 59653 57379 59687
rect 1593 59585 1627 59619
rect 6561 59585 6595 59619
rect 6837 59585 6871 59619
rect 6929 59585 6963 59619
rect 18797 59585 18831 59619
rect 18981 59585 19015 59619
rect 19170 59585 19204 59619
rect 24317 59585 24351 59619
rect 24501 59585 24535 59619
rect 24685 59585 24719 59619
rect 25605 59585 25639 59619
rect 25789 59585 25823 59619
rect 25978 59585 26012 59619
rect 43269 59585 43303 59619
rect 43637 59585 43671 59619
rect 58173 59585 58207 59619
rect 42717 59517 42751 59551
rect 43085 59517 43119 59551
rect 43545 59517 43579 59551
rect 1777 59381 1811 59415
rect 2513 59381 2547 59415
rect 7113 59381 7147 59415
rect 18521 59381 18555 59415
rect 19349 59381 19383 59415
rect 26157 59381 26191 59415
rect 29009 59381 29043 59415
rect 1869 59109 1903 59143
rect 40601 59041 40635 59075
rect 41061 59041 41095 59075
rect 1685 58973 1719 59007
rect 37197 58973 37231 59007
rect 37289 58973 37323 59007
rect 37565 58973 37599 59007
rect 37841 58973 37875 59007
rect 38117 58973 38151 59007
rect 40785 58973 40819 59007
rect 41153 58973 41187 59007
rect 57161 58973 57195 59007
rect 57897 58973 57931 59007
rect 36737 58905 36771 58939
rect 58173 58905 58207 58939
rect 40417 58837 40451 58871
rect 57345 58837 57379 58871
rect 58173 58565 58207 58599
rect 1593 58497 1627 58531
rect 40601 58497 40635 58531
rect 40785 58497 40819 58531
rect 41153 58497 41187 58531
rect 41337 58497 41371 58531
rect 1777 58429 1811 58463
rect 40417 58293 40451 58327
rect 58265 58293 58299 58327
rect 58265 57953 58299 57987
rect 1593 57885 1627 57919
rect 1869 57817 1903 57851
rect 57989 57817 58023 57851
rect 1593 57409 1627 57443
rect 1777 57205 1811 57239
rect 35265 56933 35299 56967
rect 33977 56865 34011 56899
rect 1593 56797 1627 56831
rect 33517 56797 33551 56831
rect 33701 56797 33735 56831
rect 34069 56797 34103 56831
rect 35633 56797 35667 56831
rect 35909 56797 35943 56831
rect 36001 56797 36035 56831
rect 36277 56797 36311 56831
rect 36553 56797 36587 56831
rect 57897 56797 57931 56831
rect 58173 56729 58207 56763
rect 1777 56661 1811 56695
rect 33333 56661 33367 56695
rect 58173 56389 58207 56423
rect 29285 56321 29319 56355
rect 29653 56321 29687 56355
rect 29837 56321 29871 56355
rect 35633 56321 35667 56355
rect 36461 56321 36495 56355
rect 40969 56321 41003 56355
rect 41153 56321 41187 56355
rect 41521 56321 41555 56355
rect 29193 56253 29227 56287
rect 41429 56253 41463 56287
rect 28733 56117 28767 56151
rect 40785 56117 40819 56151
rect 58265 56117 58299 56151
rect 58357 55913 58391 55947
rect 27261 55709 27295 55743
rect 27353 55709 27387 55743
rect 27629 55709 27663 55743
rect 27813 55709 27847 55743
rect 1685 55641 1719 55675
rect 26617 55641 26651 55675
rect 1777 55573 1811 55607
rect 1777 55369 1811 55403
rect 1593 55233 1627 55267
rect 40417 55233 40451 55267
rect 40601 55233 40635 55267
rect 40969 55233 41003 55267
rect 40049 55165 40083 55199
rect 40877 55165 40911 55199
rect 23581 54689 23615 54723
rect 23489 54621 23523 54655
rect 23857 54621 23891 54655
rect 24041 54621 24075 54655
rect 58357 54621 58391 54655
rect 1685 54553 1719 54587
rect 22845 54553 22879 54587
rect 1777 54485 1811 54519
rect 1593 54145 1627 54179
rect 1777 53941 1811 53975
rect 40509 53601 40543 53635
rect 40693 53533 40727 53567
rect 41061 53533 41095 53567
rect 41245 53533 41279 53567
rect 40325 53397 40359 53431
rect 23305 53125 23339 53159
rect 23397 53125 23431 53159
rect 1685 53057 1719 53091
rect 23121 53057 23155 53091
rect 23541 53057 23575 53091
rect 24317 53057 24351 53091
rect 24593 52989 24627 53023
rect 1777 52853 1811 52887
rect 23673 52853 23707 52887
rect 58357 52853 58391 52887
rect 1869 52513 1903 52547
rect 1593 52445 1627 52479
rect 1869 52037 1903 52071
rect 7021 52037 7055 52071
rect 1685 51969 1719 52003
rect 6837 51969 6871 52003
rect 7113 51969 7147 52003
rect 6653 51765 6687 51799
rect 58357 51357 58391 51391
rect 1685 51289 1719 51323
rect 1869 51289 1903 51323
rect 3985 50949 4019 50983
rect 3709 50881 3743 50915
rect 3893 50881 3927 50915
rect 4129 50881 4163 50915
rect 4261 50677 4295 50711
rect 57897 50269 57931 50303
rect 1685 50201 1719 50235
rect 1869 50201 1903 50235
rect 58173 50201 58207 50235
rect 1593 49793 1627 49827
rect 1777 49657 1811 49691
rect 1685 49113 1719 49147
rect 57989 49113 58023 49147
rect 1777 49045 1811 49079
rect 58081 49045 58115 49079
rect 1685 48705 1719 48739
rect 1869 48569 1903 48603
rect 56977 48093 57011 48127
rect 57253 48025 57287 48059
rect 57989 48025 58023 48059
rect 56609 47957 56643 47991
rect 58081 47957 58115 47991
rect 1685 47617 1719 47651
rect 1869 47481 1903 47515
rect 1593 47005 1627 47039
rect 57897 47005 57931 47039
rect 58173 46937 58207 46971
rect 1777 46869 1811 46903
rect 1593 46529 1627 46563
rect 1777 46325 1811 46359
rect 1685 45849 1719 45883
rect 57989 45849 58023 45883
rect 1777 45781 1811 45815
rect 58081 45781 58115 45815
rect 17969 45509 18003 45543
rect 36553 45509 36587 45543
rect 17601 45441 17635 45475
rect 17694 45441 17728 45475
rect 17877 45441 17911 45475
rect 18107 45441 18141 45475
rect 36277 45441 36311 45475
rect 36461 45441 36495 45475
rect 36697 45441 36731 45475
rect 36829 45305 36863 45339
rect 18245 45237 18279 45271
rect 38209 45033 38243 45067
rect 1593 44829 1627 44863
rect 37657 44829 37691 44863
rect 37933 44829 37967 44863
rect 38030 44829 38064 44863
rect 56977 44829 57011 44863
rect 1869 44761 1903 44795
rect 37841 44761 37875 44795
rect 57253 44761 57287 44795
rect 57989 44761 58023 44795
rect 58265 44693 58299 44727
rect 1685 44353 1719 44387
rect 1777 44149 1811 44183
rect 35449 43877 35483 43911
rect 35817 43809 35851 43843
rect 34897 43741 34931 43775
rect 35317 43741 35351 43775
rect 57897 43741 57931 43775
rect 1685 43673 1719 43707
rect 35081 43673 35115 43707
rect 35173 43673 35207 43707
rect 58173 43673 58207 43707
rect 1777 43605 1811 43639
rect 34253 43333 34287 43367
rect 1593 43265 1627 43299
rect 33977 43265 34011 43299
rect 34161 43265 34195 43299
rect 34397 43265 34431 43299
rect 1777 43061 1811 43095
rect 34529 43061 34563 43095
rect 37473 42789 37507 42823
rect 33333 42653 33367 42687
rect 33425 42653 33459 42687
rect 33701 42653 33735 42687
rect 33977 42653 34011 42687
rect 34161 42653 34195 42687
rect 36921 42653 36955 42687
rect 37197 42653 37231 42687
rect 37289 42653 37323 42687
rect 37105 42585 37139 42619
rect 57069 42585 57103 42619
rect 57989 42585 58023 42619
rect 58357 42585 58391 42619
rect 32965 42517 32999 42551
rect 57161 42517 57195 42551
rect 1685 42177 1719 42211
rect 1869 42041 1903 42075
rect 25145 41633 25179 41667
rect 25237 41565 25271 41599
rect 25605 41565 25639 41599
rect 25697 41565 25731 41599
rect 56977 41565 57011 41599
rect 1685 41497 1719 41531
rect 24593 41497 24627 41531
rect 57253 41497 57287 41531
rect 57989 41497 58023 41531
rect 1777 41429 1811 41463
rect 58081 41429 58115 41463
rect 1685 41089 1719 41123
rect 1777 40885 1811 40919
rect 56977 40477 57011 40511
rect 57897 40477 57931 40511
rect 1685 40409 1719 40443
rect 57253 40409 57287 40443
rect 58173 40409 58207 40443
rect 1777 40341 1811 40375
rect 2881 39525 2915 39559
rect 1869 39457 1903 39491
rect 2329 39389 2363 39423
rect 2605 39389 2639 39423
rect 2743 39389 2777 39423
rect 20637 39389 20671 39423
rect 20913 39389 20947 39423
rect 21005 39389 21039 39423
rect 1685 39321 1719 39355
rect 2513 39321 2547 39355
rect 20821 39321 20855 39355
rect 57069 39321 57103 39355
rect 57989 39321 58023 39355
rect 21189 39253 21223 39287
rect 57161 39253 57195 39287
rect 58081 39253 58115 39287
rect 34345 38981 34379 39015
rect 1685 38913 1719 38947
rect 34069 38913 34103 38947
rect 34253 38913 34287 38947
rect 34442 38913 34476 38947
rect 1869 38777 1903 38811
rect 34621 38777 34655 38811
rect 22753 38301 22787 38335
rect 22901 38301 22935 38335
rect 23218 38301 23252 38335
rect 57897 38301 57931 38335
rect 1685 38233 1719 38267
rect 23029 38233 23063 38267
rect 23121 38233 23155 38267
rect 58173 38233 58207 38267
rect 1777 38165 1811 38199
rect 23397 38165 23431 38199
rect 20913 37961 20947 37995
rect 19625 37893 19659 37927
rect 1685 37825 1719 37859
rect 4813 37825 4847 37859
rect 4997 37825 5031 37859
rect 19257 37825 19291 37859
rect 19350 37825 19384 37859
rect 19533 37825 19567 37859
rect 19741 37825 19775 37859
rect 20729 37825 20763 37859
rect 21005 37825 21039 37859
rect 58081 37825 58115 37859
rect 20269 37757 20303 37791
rect 1869 37689 1903 37723
rect 5181 37621 5215 37655
rect 19901 37621 19935 37655
rect 20545 37621 20579 37655
rect 58265 37621 58299 37655
rect 20361 37417 20395 37451
rect 20545 37349 20579 37383
rect 20085 37281 20119 37315
rect 2053 37213 2087 37247
rect 2421 37213 2455 37247
rect 18429 37213 18463 37247
rect 20453 37213 20487 37247
rect 20637 37213 20671 37247
rect 20821 37213 20855 37247
rect 57897 37213 57931 37247
rect 2237 37145 2271 37179
rect 2329 37145 2363 37179
rect 18705 37145 18739 37179
rect 58173 37145 58207 37179
rect 2605 37077 2639 37111
rect 53757 36873 53791 36907
rect 2329 36805 2363 36839
rect 6653 36805 6687 36839
rect 19073 36805 19107 36839
rect 2053 36737 2087 36771
rect 2237 36737 2271 36771
rect 2421 36737 2455 36771
rect 3065 36737 3099 36771
rect 6929 36737 6963 36771
rect 17969 36737 18003 36771
rect 18797 36737 18831 36771
rect 18981 36737 19015 36771
rect 19211 36737 19245 36771
rect 19993 36737 20027 36771
rect 20269 36737 20303 36771
rect 23581 36737 23615 36771
rect 54309 36737 54343 36771
rect 54677 36737 54711 36771
rect 6745 36669 6779 36703
rect 18061 36669 18095 36703
rect 20453 36669 20487 36703
rect 24225 36669 24259 36703
rect 54401 36669 54435 36703
rect 54585 36669 54619 36703
rect 2605 36601 2639 36635
rect 18337 36601 18371 36635
rect 19349 36601 19383 36635
rect 20085 36601 20119 36635
rect 3249 36533 3283 36567
rect 6653 36533 6687 36567
rect 7113 36533 7147 36567
rect 18153 36533 18187 36567
rect 3065 36329 3099 36363
rect 54033 36329 54067 36363
rect 1869 36261 1903 36295
rect 18889 36261 18923 36295
rect 21189 36261 21223 36295
rect 2513 36125 2547 36159
rect 2881 36125 2915 36159
rect 5549 36125 5583 36159
rect 5641 36125 5675 36159
rect 5917 36125 5951 36159
rect 6193 36125 6227 36159
rect 6377 36125 6411 36159
rect 18061 36125 18095 36159
rect 18337 36125 18371 36159
rect 18613 36125 18647 36159
rect 18705 36125 18739 36159
rect 19993 36125 20027 36159
rect 20141 36125 20175 36159
rect 20361 36125 20395 36159
rect 20499 36125 20533 36159
rect 21097 36125 21131 36159
rect 21373 36125 21407 36159
rect 22477 36125 22511 36159
rect 22753 36125 22787 36159
rect 22845 36125 22879 36159
rect 23673 36125 23707 36159
rect 40325 36125 40359 36159
rect 40693 36125 40727 36159
rect 53481 36125 53515 36159
rect 53757 36125 53791 36159
rect 53901 36125 53935 36159
rect 1685 36057 1719 36091
rect 2697 36057 2731 36091
rect 2789 36057 2823 36091
rect 18521 36057 18555 36091
rect 20269 36057 20303 36091
rect 22661 36057 22695 36091
rect 23489 36057 23523 36091
rect 24041 36057 24075 36091
rect 40509 36057 40543 36091
rect 40601 36057 40635 36091
rect 53665 36057 53699 36091
rect 57989 36057 58023 36091
rect 58357 36057 58391 36091
rect 5181 35989 5215 36023
rect 20637 35989 20671 36023
rect 21557 35989 21591 36023
rect 23029 35989 23063 36023
rect 40877 35989 40911 36023
rect 24317 35785 24351 35819
rect 1869 35717 1903 35751
rect 19809 35717 19843 35751
rect 23213 35717 23247 35751
rect 23857 35717 23891 35751
rect 1685 35649 1719 35683
rect 19533 35649 19567 35683
rect 19717 35649 19751 35683
rect 19901 35649 19935 35683
rect 20637 35649 20671 35683
rect 22201 35649 22235 35683
rect 24133 35649 24167 35683
rect 36001 35649 36035 35683
rect 21189 35581 21223 35615
rect 23949 35581 23983 35615
rect 36277 35581 36311 35615
rect 20085 35445 20119 35479
rect 23857 35445 23891 35479
rect 20085 35241 20119 35275
rect 21833 35241 21867 35275
rect 1869 35173 1903 35207
rect 20729 35173 20763 35207
rect 35633 35173 35667 35207
rect 40601 35173 40635 35207
rect 20361 35105 20395 35139
rect 22017 35105 22051 35139
rect 19533 35037 19567 35071
rect 19809 35037 19843 35071
rect 19901 35037 19935 35071
rect 20637 35037 20671 35071
rect 20913 35037 20947 35071
rect 21833 35037 21867 35071
rect 22109 35037 22143 35071
rect 36001 35037 36035 35071
rect 36093 35037 36127 35071
rect 36369 35037 36403 35071
rect 36645 35037 36679 35071
rect 36829 35037 36863 35071
rect 40049 35037 40083 35071
rect 40325 35037 40359 35071
rect 40417 35037 40451 35071
rect 57897 35037 57931 35071
rect 1685 34969 1719 35003
rect 19717 34969 19751 35003
rect 40233 34969 40267 35003
rect 58173 34969 58207 35003
rect 21097 34901 21131 34935
rect 22293 34901 22327 34935
rect 23949 34697 23983 34731
rect 58265 34697 58299 34731
rect 22477 34629 22511 34663
rect 26341 34629 26375 34663
rect 22109 34561 22143 34595
rect 22257 34561 22291 34595
rect 22385 34561 22419 34595
rect 22615 34561 22649 34595
rect 23397 34561 23431 34595
rect 23581 34561 23615 34595
rect 23673 34561 23707 34595
rect 23765 34561 23799 34595
rect 25973 34561 26007 34595
rect 26121 34561 26155 34595
rect 26249 34561 26283 34595
rect 26438 34561 26472 34595
rect 58081 34561 58115 34595
rect 23029 34493 23063 34527
rect 22753 34357 22787 34391
rect 26617 34357 26651 34391
rect 21465 34085 21499 34119
rect 22569 34017 22603 34051
rect 20821 33949 20855 33983
rect 20969 33949 21003 33983
rect 21286 33949 21320 33983
rect 22017 33949 22051 33983
rect 22477 33949 22511 33983
rect 1685 33881 1719 33915
rect 21097 33881 21131 33915
rect 21189 33881 21223 33915
rect 1777 33813 1811 33847
rect 1869 33541 1903 33575
rect 1685 33473 1719 33507
rect 22017 33473 22051 33507
rect 22109 33473 22143 33507
rect 22293 33473 22327 33507
rect 22753 33405 22787 33439
rect 26801 32997 26835 33031
rect 22845 32929 22879 32963
rect 58173 32929 58207 32963
rect 22569 32861 22603 32895
rect 26709 32861 26743 32895
rect 26985 32861 27019 32895
rect 57897 32861 57931 32895
rect 1685 32793 1719 32827
rect 57069 32793 57103 32827
rect 1777 32725 1811 32759
rect 27169 32725 27203 32759
rect 57161 32725 57195 32759
rect 1685 32385 1719 32419
rect 1777 32181 1811 32215
rect 25881 31909 25915 31943
rect 25053 31841 25087 31875
rect 58081 31841 58115 31875
rect 25329 31773 25363 31807
rect 25605 31773 25639 31807
rect 25697 31773 25731 31807
rect 57897 31773 57931 31807
rect 25513 31705 25547 31739
rect 25973 31433 26007 31467
rect 25605 31365 25639 31399
rect 25697 31365 25731 31399
rect 1685 31297 1719 31331
rect 19625 31297 19659 31331
rect 19901 31297 19935 31331
rect 25329 31297 25363 31331
rect 25477 31297 25511 31331
rect 25794 31297 25828 31331
rect 58081 31297 58115 31331
rect 20085 31229 20119 31263
rect 19717 31161 19751 31195
rect 1777 31093 1811 31127
rect 58265 31093 58299 31127
rect 20085 30889 20119 30923
rect 19441 30685 19475 30719
rect 19589 30685 19623 30719
rect 19947 30685 19981 30719
rect 1685 30617 1719 30651
rect 19717 30617 19751 30651
rect 19809 30617 19843 30651
rect 1777 30549 1811 30583
rect 23673 30277 23707 30311
rect 23765 30277 23799 30311
rect 25329 30277 25363 30311
rect 1593 30209 1627 30243
rect 23489 30209 23523 30243
rect 23857 30209 23891 30243
rect 25145 30209 25179 30243
rect 25421 30209 25455 30243
rect 25513 30209 25547 30243
rect 1777 30141 1811 30175
rect 24041 30005 24075 30039
rect 25697 30005 25731 30039
rect 25881 29801 25915 29835
rect 25973 29801 26007 29835
rect 24041 29733 24075 29767
rect 58173 29665 58207 29699
rect 1593 29597 1627 29631
rect 23489 29597 23523 29631
rect 23857 29597 23891 29631
rect 24593 29597 24627 29631
rect 24869 29597 24903 29631
rect 24961 29597 24995 29631
rect 26065 29597 26099 29631
rect 26157 29597 26191 29631
rect 26341 29597 26375 29631
rect 57897 29597 57931 29631
rect 1869 29529 1903 29563
rect 23673 29529 23707 29563
rect 23765 29529 23799 29563
rect 24777 29529 24811 29563
rect 57069 29529 57103 29563
rect 25145 29461 25179 29495
rect 25605 29461 25639 29495
rect 57161 29461 57195 29495
rect 17969 29189 18003 29223
rect 24317 29189 24351 29223
rect 17785 29121 17819 29155
rect 18245 29121 18279 29155
rect 24547 29121 24581 29155
rect 25605 29121 25639 29155
rect 25881 29121 25915 29155
rect 24464 29053 24498 29087
rect 24685 29053 24719 29087
rect 25697 29053 25731 29087
rect 26341 29053 26375 29087
rect 24777 28985 24811 29019
rect 1593 28509 1627 28543
rect 57897 28509 57931 28543
rect 1869 28441 1903 28475
rect 58173 28441 58207 28475
rect 2881 28169 2915 28203
rect 1593 28033 1627 28067
rect 2513 28033 2547 28067
rect 2667 28033 2701 28067
rect 58081 28033 58115 28067
rect 1777 27965 1811 27999
rect 58265 27829 58299 27863
rect 1593 27421 1627 27455
rect 1869 27353 1903 27387
rect 2881 27081 2915 27115
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 2667 26945 2701 26979
rect 1777 26877 1811 26911
rect 58173 26401 58207 26435
rect 57897 26333 57931 26367
rect 57069 26265 57103 26299
rect 57161 26197 57195 26231
rect 18153 25925 18187 25959
rect 1593 25857 1627 25891
rect 17969 25857 18003 25891
rect 1777 25789 1811 25823
rect 18245 25789 18279 25823
rect 2881 25313 2915 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 2667 25245 2701 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 58173 25177 58207 25211
rect 1593 24769 1627 24803
rect 58081 24769 58115 24803
rect 1777 24701 1811 24735
rect 58265 24565 58299 24599
rect 4169 24361 4203 24395
rect 1593 24157 1627 24191
rect 3985 24157 4019 24191
rect 4139 24157 4173 24191
rect 1869 24089 1903 24123
rect 17233 23817 17267 23851
rect 16865 23681 16899 23715
rect 17019 23681 17053 23715
rect 26801 23273 26835 23307
rect 23397 23205 23431 23239
rect 18521 23137 18555 23171
rect 26433 23137 26467 23171
rect 58173 23137 58207 23171
rect 1593 23069 1627 23103
rect 18153 23069 18187 23103
rect 18613 23069 18647 23103
rect 24593 23069 24627 23103
rect 26617 23069 26651 23103
rect 57897 23069 57931 23103
rect 1869 23001 1903 23035
rect 23029 23001 23063 23035
rect 24860 23001 24894 23035
rect 23489 22933 23523 22967
rect 25973 22933 26007 22967
rect 17693 22661 17727 22695
rect 25605 22661 25639 22695
rect 1593 22593 1627 22627
rect 17509 22593 17543 22627
rect 22845 22593 22879 22627
rect 27353 22593 27387 22627
rect 58081 22593 58115 22627
rect 1777 22525 1811 22559
rect 17785 22525 17819 22559
rect 27169 22525 27203 22559
rect 25881 22457 25915 22491
rect 24041 22389 24075 22423
rect 26065 22389 26099 22423
rect 27537 22389 27571 22423
rect 58265 22389 58299 22423
rect 23949 22185 23983 22219
rect 17693 22117 17727 22151
rect 22753 22117 22787 22151
rect 17785 22049 17819 22083
rect 22477 22049 22511 22083
rect 23765 22049 23799 22083
rect 1593 21981 1627 22015
rect 17509 21981 17543 22015
rect 22385 21981 22419 22015
rect 23673 21981 23707 22015
rect 24593 21981 24627 22015
rect 27353 21981 27387 22015
rect 27721 21981 27755 22015
rect 28457 21981 28491 22015
rect 28549 21981 28583 22015
rect 57897 21981 57931 22015
rect 1869 21913 1903 21947
rect 27537 21913 27571 21947
rect 27629 21913 27663 21947
rect 58173 21913 58207 21947
rect 25789 21845 25823 21879
rect 27905 21845 27939 21879
rect 28733 21845 28767 21879
rect 22753 21641 22787 21675
rect 23305 21641 23339 21675
rect 25697 21641 25731 21675
rect 28549 21641 28583 21675
rect 20913 21573 20947 21607
rect 21129 21573 21163 21607
rect 27436 21573 27470 21607
rect 1685 21505 1719 21539
rect 22385 21505 22419 21539
rect 23581 21505 23615 21539
rect 24317 21505 24351 21539
rect 29193 21505 29227 21539
rect 58081 21505 58115 21539
rect 22293 21437 22327 21471
rect 23489 21437 23523 21471
rect 23673 21437 23707 21471
rect 23765 21437 23799 21471
rect 27169 21437 27203 21471
rect 29009 21437 29043 21471
rect 1777 21301 1811 21335
rect 21097 21301 21131 21335
rect 21281 21301 21315 21335
rect 29377 21301 29411 21335
rect 58265 21301 58299 21335
rect 21097 21097 21131 21131
rect 29745 21097 29779 21131
rect 21281 21029 21315 21063
rect 27537 20961 27571 20995
rect 30297 20961 30331 20995
rect 20085 20893 20119 20927
rect 20269 20893 20303 20927
rect 21741 20893 21775 20927
rect 24777 20893 24811 20927
rect 20913 20825 20947 20859
rect 27077 20825 27111 20859
rect 27782 20825 27816 20859
rect 20453 20757 20487 20791
rect 21113 20757 21147 20791
rect 22937 20757 22971 20791
rect 28917 20757 28951 20791
rect 30113 20757 30147 20791
rect 30205 20757 30239 20791
rect 30849 20757 30883 20791
rect 19533 20553 19567 20587
rect 22845 20553 22879 20587
rect 26433 20553 26467 20587
rect 27445 20553 27479 20587
rect 22753 20485 22787 20519
rect 1593 20417 1627 20451
rect 18705 20417 18739 20451
rect 18889 20417 18923 20451
rect 19349 20417 19383 20451
rect 19533 20417 19567 20451
rect 20260 20417 20294 20451
rect 22661 20417 22695 20451
rect 23581 20417 23615 20451
rect 26341 20417 26375 20451
rect 26525 20417 26559 20451
rect 27353 20417 27387 20451
rect 27537 20417 27571 20451
rect 28457 20417 28491 20451
rect 28724 20417 28758 20451
rect 30389 20417 30423 20451
rect 30645 20417 30679 20451
rect 32321 20417 32355 20451
rect 32505 20417 32539 20451
rect 38761 20417 38795 20451
rect 1777 20349 1811 20383
rect 19993 20349 20027 20383
rect 23029 20349 23063 20383
rect 38577 20349 38611 20383
rect 22477 20281 22511 20315
rect 27169 20281 27203 20315
rect 18705 20213 18739 20247
rect 21373 20213 21407 20247
rect 24777 20213 24811 20247
rect 27721 20213 27755 20247
rect 29837 20213 29871 20247
rect 31769 20213 31803 20247
rect 32689 20213 32723 20247
rect 38945 20213 38979 20247
rect 25145 20009 25179 20043
rect 38577 20009 38611 20043
rect 18613 19941 18647 19975
rect 21189 19941 21223 19975
rect 29837 19941 29871 19975
rect 24041 19873 24075 19907
rect 27353 19873 27387 19907
rect 32413 19873 32447 19907
rect 39129 19873 39163 19907
rect 40509 19873 40543 19907
rect 48145 19873 48179 19907
rect 58173 19873 58207 19907
rect 1593 19805 1627 19839
rect 17969 19805 18003 19839
rect 18153 19805 18187 19839
rect 18613 19805 18647 19839
rect 18889 19805 18923 19839
rect 19809 19805 19843 19839
rect 21741 19805 21775 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 26249 19805 26283 19839
rect 30113 19805 30147 19839
rect 31309 19805 31343 19839
rect 36461 19805 36495 19839
rect 36645 19805 36679 19839
rect 38301 19805 38335 19839
rect 39037 19805 39071 19839
rect 40713 19805 40747 19839
rect 48329 19805 48363 19839
rect 57897 19805 57931 19839
rect 1869 19737 1903 19771
rect 20076 19737 20110 19771
rect 24593 19737 24627 19771
rect 30389 19737 30423 19771
rect 18061 19669 18095 19703
rect 18797 19669 18831 19703
rect 24869 19669 24903 19703
rect 30297 19669 30331 19703
rect 36829 19669 36863 19703
rect 38945 19669 38979 19703
rect 40877 19669 40911 19703
rect 48513 19669 48547 19703
rect 20361 19465 20395 19499
rect 23765 19465 23799 19499
rect 25513 19465 25547 19499
rect 27261 19465 27295 19499
rect 30021 19465 30055 19499
rect 33517 19465 33551 19499
rect 35081 19465 35115 19499
rect 35449 19465 35483 19499
rect 38669 19465 38703 19499
rect 40509 19465 40543 19499
rect 58265 19465 58299 19499
rect 27629 19397 27663 19431
rect 48145 19397 48179 19431
rect 1593 19329 1627 19363
rect 1869 19329 1903 19363
rect 17509 19329 17543 19363
rect 17693 19329 17727 19363
rect 18337 19329 18371 19363
rect 19165 19329 19199 19363
rect 22385 19329 22419 19363
rect 22652 19329 22686 19363
rect 24317 19329 24351 19363
rect 28825 19329 28859 19363
rect 32321 19329 32355 19363
rect 36461 19329 36495 19363
rect 37473 19329 37507 19363
rect 40877 19329 40911 19363
rect 42717 19329 42751 19363
rect 47869 19329 47903 19363
rect 48053 19329 48087 19363
rect 48283 19329 48317 19363
rect 48881 19329 48915 19363
rect 49065 19329 49099 19363
rect 58081 19329 58115 19363
rect 18429 19261 18463 19295
rect 18705 19261 18739 19295
rect 27721 19261 27755 19295
rect 27905 19261 27939 19295
rect 35541 19261 35575 19295
rect 35725 19261 35759 19295
rect 36277 19261 36311 19295
rect 40969 19261 41003 19295
rect 41153 19261 41187 19295
rect 2421 19125 2455 19159
rect 17509 19125 17543 19159
rect 36645 19125 36679 19159
rect 40233 19125 40267 19159
rect 42993 19125 43027 19159
rect 48421 19125 48455 19159
rect 49249 19125 49283 19159
rect 22937 18921 22971 18955
rect 32597 18921 32631 18955
rect 48421 18921 48455 18955
rect 21281 18853 21315 18887
rect 30297 18853 30331 18887
rect 39681 18853 39715 18887
rect 40141 18853 40175 18887
rect 41889 18853 41923 18887
rect 42441 18853 42475 18887
rect 17601 18785 17635 18819
rect 17877 18785 17911 18819
rect 18521 18785 18555 18819
rect 18705 18785 18739 18819
rect 18797 18785 18831 18819
rect 24593 18785 24627 18819
rect 36921 18785 36955 18819
rect 39129 18785 39163 18819
rect 42993 18785 43027 18819
rect 1593 18717 1627 18751
rect 16681 18717 16715 18751
rect 16865 18717 16899 18751
rect 17509 18717 17543 18751
rect 18613 18717 18647 18751
rect 19901 18717 19935 18751
rect 21741 18717 21775 18751
rect 24860 18717 24894 18751
rect 26893 18717 26927 18751
rect 30573 18717 30607 18751
rect 31401 18717 31435 18751
rect 34897 18717 34931 18751
rect 35081 18717 35115 18751
rect 35817 18717 35851 18751
rect 38945 18717 38979 18751
rect 40509 18717 40543 18751
rect 40776 18717 40810 18751
rect 42809 18717 42843 18751
rect 43637 18717 43671 18751
rect 44005 18717 44039 18751
rect 45385 18717 45419 18751
rect 45569 18717 45603 18751
rect 47869 18717 47903 18751
rect 48237 18717 48271 18751
rect 48881 18717 48915 18751
rect 49019 18717 49053 18751
rect 49249 18717 49283 18751
rect 57897 18717 57931 18751
rect 1869 18649 1903 18683
rect 20168 18649 20202 18683
rect 30849 18649 30883 18683
rect 42901 18649 42935 18683
rect 43821 18649 43855 18683
rect 43913 18649 43947 18683
rect 48053 18649 48087 18683
rect 48145 18649 48179 18683
rect 49157 18649 49191 18683
rect 58173 18649 58207 18683
rect 2421 18581 2455 18615
rect 16773 18581 16807 18615
rect 18337 18581 18371 18615
rect 25973 18581 26007 18615
rect 28089 18581 28123 18615
rect 30757 18581 30791 18615
rect 35265 18581 35299 18615
rect 38577 18581 38611 18615
rect 39037 18581 39071 18615
rect 44189 18581 44223 18615
rect 45753 18581 45787 18615
rect 49433 18581 49467 18615
rect 18613 18377 18647 18411
rect 24501 18377 24535 18411
rect 27169 18377 27203 18411
rect 29469 18377 29503 18411
rect 31401 18377 31435 18411
rect 36461 18377 36495 18411
rect 37473 18377 37507 18411
rect 40141 18377 40175 18411
rect 40693 18377 40727 18411
rect 44281 18377 44315 18411
rect 46857 18377 46891 18411
rect 49525 18377 49559 18411
rect 58265 18377 58299 18411
rect 22661 18309 22695 18343
rect 35348 18309 35382 18343
rect 41061 18309 41095 18343
rect 45744 18309 45778 18343
rect 48412 18309 48446 18343
rect 15393 18241 15427 18275
rect 15577 18241 15611 18275
rect 17500 18241 17534 18275
rect 19165 18241 19199 18275
rect 23305 18241 23339 18275
rect 26249 18241 26283 18275
rect 27346 18247 27380 18281
rect 27629 18241 27663 18275
rect 27813 18241 27847 18275
rect 28273 18241 28307 18275
rect 32321 18241 32355 18275
rect 37841 18241 37875 18275
rect 39028 18241 39062 18275
rect 41705 18241 41739 18275
rect 43157 18241 43191 18275
rect 50261 18241 50295 18275
rect 58081 18241 58115 18275
rect 17233 18173 17267 18207
rect 20269 18173 20303 18207
rect 22569 18173 22603 18207
rect 22753 18173 22787 18207
rect 26341 18173 26375 18207
rect 31493 18173 31527 18207
rect 31585 18173 31619 18207
rect 35081 18173 35115 18207
rect 37933 18173 37967 18207
rect 38117 18173 38151 18207
rect 38761 18173 38795 18207
rect 40509 18173 40543 18207
rect 41153 18173 41187 18207
rect 41245 18173 41279 18207
rect 42901 18173 42935 18207
rect 45477 18173 45511 18207
rect 48145 18173 48179 18207
rect 50077 18173 50111 18207
rect 22201 18105 22235 18139
rect 26617 18105 26651 18139
rect 15761 18037 15795 18071
rect 31033 18037 31067 18071
rect 33517 18037 33551 18071
rect 50445 18037 50479 18071
rect 26801 17833 26835 17867
rect 28457 17833 28491 17867
rect 33057 17833 33091 17867
rect 42441 17833 42475 17867
rect 44281 17833 44315 17867
rect 45753 17833 45787 17867
rect 51733 17833 51767 17867
rect 16037 17765 16071 17799
rect 20821 17765 20855 17799
rect 24593 17765 24627 17799
rect 15117 17697 15151 17731
rect 24961 17697 24995 17731
rect 29101 17697 29135 17731
rect 31769 17697 31803 17731
rect 33701 17697 33735 17731
rect 48145 17697 48179 17731
rect 1593 17629 1627 17663
rect 14289 17629 14323 17663
rect 14473 17629 14507 17663
rect 15025 17629 15059 17663
rect 15209 17629 15243 17663
rect 16589 17629 16623 17663
rect 19441 17629 19475 17663
rect 21741 17629 21775 17663
rect 24777 17629 24811 17663
rect 24869 17629 24903 17663
rect 25053 17629 25087 17663
rect 25605 17629 25639 17663
rect 28825 17629 28859 17663
rect 30297 17629 30331 17663
rect 33517 17629 33551 17663
rect 34897 17629 34931 17663
rect 35909 17629 35943 17663
rect 37841 17629 37875 17663
rect 40049 17629 40083 17663
rect 42165 17629 42199 17663
rect 42257 17629 42291 17663
rect 42901 17629 42935 17663
rect 45201 17629 45235 17663
rect 45569 17629 45603 17663
rect 47133 17629 47167 17663
rect 47409 17629 47443 17663
rect 47501 17629 47535 17663
rect 50353 17629 50387 17663
rect 1869 17561 1903 17595
rect 15669 17561 15703 17595
rect 18889 17561 18923 17595
rect 19686 17561 19720 17595
rect 24041 17561 24075 17595
rect 35173 17561 35207 17595
rect 36176 17561 36210 17595
rect 38108 17561 38142 17595
rect 40316 17561 40350 17595
rect 43168 17561 43202 17595
rect 45385 17561 45419 17595
rect 45477 17561 45511 17595
rect 47317 17561 47351 17595
rect 48412 17561 48446 17595
rect 50598 17561 50632 17595
rect 14381 17493 14415 17527
rect 16129 17493 16163 17527
rect 28917 17493 28951 17527
rect 33425 17493 33459 17527
rect 37289 17493 37323 17527
rect 39221 17493 39255 17527
rect 41429 17493 41463 17527
rect 47685 17493 47719 17527
rect 49525 17493 49559 17527
rect 20361 17289 20395 17323
rect 22385 17289 22419 17323
rect 24133 17289 24167 17323
rect 25881 17289 25915 17323
rect 26249 17289 26283 17323
rect 27537 17289 27571 17323
rect 33793 17289 33827 17323
rect 37841 17289 37875 17323
rect 39773 17289 39807 17323
rect 40693 17289 40727 17323
rect 45569 17289 45603 17323
rect 49893 17289 49927 17323
rect 17592 17221 17626 17255
rect 35725 17221 35759 17255
rect 35909 17221 35943 17255
rect 41889 17221 41923 17255
rect 42993 17221 43027 17255
rect 48780 17221 48814 17255
rect 1593 17153 1627 17187
rect 14013 17153 14047 17187
rect 19165 17153 19199 17187
rect 22201 17153 22235 17187
rect 22937 17153 22971 17187
rect 26341 17153 26375 17187
rect 27353 17153 27387 17187
rect 27997 17153 28031 17187
rect 31401 17153 31435 17187
rect 31493 17153 31527 17187
rect 32597 17153 32631 17187
rect 36737 17153 36771 17187
rect 37473 17153 37507 17187
rect 37657 17153 37691 17187
rect 38393 17153 38427 17187
rect 38660 17153 38694 17187
rect 40785 17153 40819 17187
rect 41705 17153 41739 17187
rect 42717 17153 42751 17187
rect 42901 17153 42935 17187
rect 43085 17153 43119 17187
rect 44456 17153 44490 17187
rect 1777 17085 1811 17119
rect 17325 17085 17359 17119
rect 22017 17085 22051 17119
rect 26525 17085 26559 17119
rect 27169 17085 27203 17119
rect 31585 17085 31619 17119
rect 36001 17085 36035 17119
rect 36553 17085 36587 17119
rect 40969 17085 41003 17119
rect 41521 17085 41555 17119
rect 44189 17085 44223 17119
rect 48513 17085 48547 17119
rect 18705 17017 18739 17051
rect 2421 16949 2455 16983
rect 15393 16949 15427 16983
rect 29193 16949 29227 16983
rect 31033 16949 31067 16983
rect 35449 16949 35483 16983
rect 36921 16949 36955 16983
rect 40325 16949 40359 16983
rect 43269 16949 43303 16983
rect 57161 16745 57195 16779
rect 15577 16677 15611 16711
rect 25973 16677 26007 16711
rect 38117 16677 38151 16711
rect 41797 16677 41831 16711
rect 45569 16677 45603 16711
rect 13461 16609 13495 16643
rect 14841 16609 14875 16643
rect 15117 16609 15151 16643
rect 24593 16609 24627 16643
rect 29745 16609 29779 16643
rect 35541 16609 35575 16643
rect 36185 16609 36219 16643
rect 38577 16609 38611 16643
rect 38669 16609 38703 16643
rect 40877 16609 40911 16643
rect 41429 16609 41463 16643
rect 45201 16609 45235 16643
rect 47501 16609 47535 16643
rect 47869 16609 47903 16643
rect 48329 16609 48363 16643
rect 1593 16541 1627 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 14749 16541 14783 16575
rect 15945 16541 15979 16575
rect 16129 16541 16163 16575
rect 16589 16541 16623 16575
rect 18889 16541 18923 16575
rect 19901 16541 19935 16575
rect 21741 16541 21775 16575
rect 24849 16541 24883 16575
rect 26893 16541 26927 16575
rect 30012 16541 30046 16575
rect 31861 16541 31895 16575
rect 35357 16541 35391 16575
rect 41613 16541 41647 16575
rect 42901 16541 42935 16575
rect 43085 16541 43119 16575
rect 43729 16541 43763 16575
rect 43913 16541 43947 16575
rect 44097 16541 44131 16575
rect 45385 16541 45419 16575
rect 47685 16541 47719 16575
rect 48585 16541 48619 16575
rect 57897 16541 57931 16575
rect 58173 16541 58207 16575
rect 1869 16473 1903 16507
rect 15853 16473 15887 16507
rect 20168 16473 20202 16507
rect 36452 16473 36486 16507
rect 43269 16473 43303 16507
rect 44005 16473 44039 16507
rect 57069 16473 57103 16507
rect 13185 16405 13219 16439
rect 15761 16405 15795 16439
rect 21281 16405 21315 16439
rect 23121 16405 23155 16439
rect 28089 16405 28123 16439
rect 31125 16405 31159 16439
rect 33057 16405 33091 16439
rect 34897 16405 34931 16439
rect 35265 16405 35299 16439
rect 37565 16405 37599 16439
rect 38485 16405 38519 16439
rect 40233 16405 40267 16439
rect 40601 16405 40635 16439
rect 40693 16405 40727 16439
rect 44281 16405 44315 16439
rect 49709 16405 49743 16439
rect 13001 16201 13035 16235
rect 25053 16201 25087 16235
rect 29009 16201 29043 16235
rect 33701 16201 33735 16235
rect 35633 16201 35667 16235
rect 36461 16201 36495 16235
rect 41705 16201 41739 16235
rect 48697 16201 48731 16235
rect 49525 16201 49559 16235
rect 22284 16133 22318 16167
rect 27885 16133 27919 16167
rect 43085 16133 43119 16167
rect 43177 16133 43211 16167
rect 44180 16133 44214 16167
rect 48329 16133 48363 16167
rect 48421 16133 48455 16167
rect 1593 16065 1627 16099
rect 12173 16065 12207 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 13461 16065 13495 16099
rect 14013 16065 14047 16099
rect 17500 16065 17534 16099
rect 19165 16065 19199 16099
rect 22017 16065 22051 16099
rect 23857 16065 23891 16099
rect 27629 16065 27663 16099
rect 29469 16065 29503 16099
rect 32321 16065 32355 16099
rect 32577 16065 32611 16099
rect 34520 16065 34554 16099
rect 37473 16065 37507 16099
rect 37729 16065 37763 16099
rect 39589 16065 39623 16099
rect 39773 16065 39807 16099
rect 40233 16065 40267 16099
rect 40417 16065 40451 16099
rect 42901 16065 42935 16099
rect 43269 16065 43303 16099
rect 46397 16065 46431 16099
rect 48145 16065 48179 16099
rect 48513 16065 48547 16099
rect 49157 16065 49191 16099
rect 49341 16065 49375 16099
rect 1777 15997 1811 16031
rect 11989 15997 12023 16031
rect 12265 15997 12299 16031
rect 12357 15997 12391 16031
rect 12449 15997 12483 16031
rect 13369 15997 13403 16031
rect 17233 15997 17267 16031
rect 34253 15997 34287 16031
rect 36553 15997 36587 16031
rect 36645 15997 36679 16031
rect 39405 15997 39439 16031
rect 41797 15997 41831 16031
rect 41889 15997 41923 16031
rect 43913 15997 43947 16031
rect 46213 15997 46247 16031
rect 18613 15929 18647 15963
rect 36093 15929 36127 15963
rect 45293 15929 45327 15963
rect 2421 15861 2455 15895
rect 12909 15861 12943 15895
rect 15209 15861 15243 15895
rect 20361 15861 20395 15895
rect 23397 15861 23431 15895
rect 30665 15861 30699 15895
rect 38853 15861 38887 15895
rect 40601 15861 40635 15895
rect 41337 15861 41371 15895
rect 43453 15861 43487 15895
rect 46581 15861 46615 15895
rect 17785 15657 17819 15691
rect 42901 15657 42935 15691
rect 45753 15657 45787 15691
rect 48145 15657 48179 15691
rect 22569 15589 22603 15623
rect 30297 15589 30331 15623
rect 32873 15589 32907 15623
rect 37473 15589 37507 15623
rect 38669 15589 38703 15623
rect 13737 15521 13771 15555
rect 14749 15521 14783 15555
rect 25789 15521 25823 15555
rect 28089 15521 28123 15555
rect 30849 15521 30883 15555
rect 34161 15521 34195 15555
rect 35541 15521 35575 15555
rect 38117 15521 38151 15555
rect 50353 15521 50387 15555
rect 11437 15453 11471 15487
rect 14473 15453 14507 15487
rect 16589 15453 16623 15487
rect 19533 15453 19567 15487
rect 19800 15453 19834 15487
rect 21373 15453 21407 15487
rect 26341 15453 26375 15487
rect 30665 15453 30699 15487
rect 31493 15453 31527 15487
rect 34069 15453 34103 15487
rect 34897 15453 34931 15487
rect 35081 15453 35115 15487
rect 37933 15453 37967 15487
rect 38854 15431 38888 15465
rect 38946 15453 38980 15487
rect 39175 15453 39209 15487
rect 39313 15453 39347 15487
rect 41613 15453 41647 15487
rect 44189 15453 44223 15487
rect 45201 15453 45235 15487
rect 45569 15453 45603 15487
rect 49065 15453 49099 15487
rect 49433 15453 49467 15487
rect 50537 15453 50571 15487
rect 57897 15453 57931 15487
rect 16129 15385 16163 15419
rect 31760 15385 31794 15419
rect 35786 15385 35820 15419
rect 39062 15385 39096 15419
rect 40049 15385 40083 15419
rect 40233 15385 40267 15419
rect 44465 15385 44499 15419
rect 45385 15385 45419 15419
rect 45477 15385 45511 15419
rect 46857 15385 46891 15419
rect 49249 15385 49283 15419
rect 49341 15385 49375 15419
rect 58173 15385 58207 15419
rect 20913 15317 20947 15351
rect 25145 15317 25179 15351
rect 25513 15317 25547 15351
rect 25605 15317 25639 15351
rect 30757 15317 30791 15351
rect 33609 15317 33643 15351
rect 33977 15317 34011 15351
rect 34989 15317 35023 15351
rect 36921 15317 36955 15351
rect 37841 15317 37875 15351
rect 40417 15317 40451 15351
rect 49617 15317 49651 15351
rect 50721 15317 50755 15351
rect 16221 15113 16255 15147
rect 25145 15113 25179 15147
rect 29285 15113 29319 15147
rect 30849 15113 30883 15147
rect 31309 15113 31343 15147
rect 32321 15113 32355 15147
rect 41981 15113 42015 15147
rect 43085 15113 43119 15147
rect 45845 15113 45879 15147
rect 32689 15045 32723 15079
rect 32781 15045 32815 15079
rect 33968 15045 34002 15079
rect 40868 15045 40902 15079
rect 46581 15045 46615 15079
rect 48688 15045 48722 15079
rect 1593 14977 1627 15011
rect 10977 14977 11011 15011
rect 11161 14977 11195 15011
rect 14013 14977 14047 15011
rect 19165 14977 19199 15011
rect 22109 14977 22143 15011
rect 22376 14977 22410 15011
rect 23949 14977 23983 15011
rect 27261 14977 27295 15011
rect 28089 14977 28123 15011
rect 31217 14977 31251 15011
rect 35725 14977 35759 15011
rect 35909 14977 35943 15011
rect 36001 14977 36035 15011
rect 36737 14977 36771 15011
rect 37657 14977 37691 15011
rect 39221 14977 39255 15011
rect 40601 14977 40635 15011
rect 42901 14977 42935 15011
rect 43637 14977 43671 15011
rect 44005 14977 44039 15011
rect 44465 14977 44499 15011
rect 44732 14977 44766 15011
rect 46305 14977 46339 15011
rect 1777 14909 1811 14943
rect 2421 14909 2455 14943
rect 11897 14909 11931 14943
rect 12173 14909 12207 14943
rect 17049 14909 17083 14943
rect 17325 14909 17359 14943
rect 31401 14909 31435 14943
rect 32873 14909 32907 14943
rect 33701 14909 33735 14943
rect 35817 14909 35851 14943
rect 36553 14909 36587 14943
rect 36921 14909 36955 14943
rect 37473 14909 37507 14943
rect 39313 14909 39347 14943
rect 39497 14909 39531 14943
rect 42717 14909 42751 14943
rect 48421 14909 48455 14943
rect 23489 14841 23523 14875
rect 37841 14841 37875 14875
rect 49801 14841 49835 14875
rect 10977 14773 11011 14807
rect 13277 14773 13311 14807
rect 18613 14773 18647 14807
rect 21373 14773 21407 14807
rect 27537 14773 27571 14807
rect 35081 14773 35115 14807
rect 35541 14773 35575 14807
rect 38853 14773 38887 14807
rect 10977 14569 11011 14603
rect 24593 14569 24627 14603
rect 32965 14569 32999 14603
rect 34989 14569 35023 14603
rect 42717 14569 42751 14603
rect 46765 14569 46799 14603
rect 48605 14569 48639 14603
rect 20821 14501 20855 14535
rect 28089 14501 28123 14535
rect 31125 14501 31159 14535
rect 33793 14501 33827 14535
rect 36093 14501 36127 14535
rect 37473 14501 37507 14535
rect 40049 14501 40083 14535
rect 10609 14433 10643 14467
rect 12541 14433 12575 14467
rect 14473 14433 14507 14467
rect 14749 14433 14783 14467
rect 19441 14433 19475 14467
rect 28549 14433 28583 14467
rect 28733 14433 28767 14467
rect 33977 14433 34011 14467
rect 34161 14433 34195 14467
rect 35541 14433 35575 14467
rect 35633 14433 35667 14467
rect 35909 14433 35943 14467
rect 38025 14433 38059 14467
rect 40693 14433 40727 14467
rect 1593 14365 1627 14399
rect 10793 14365 10827 14399
rect 11437 14365 11471 14399
rect 16589 14365 16623 14399
rect 21741 14365 21775 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 25329 14365 25363 14399
rect 28457 14365 28491 14399
rect 29745 14365 29779 14399
rect 31585 14365 31619 14399
rect 34069 14365 34103 14399
rect 34253 14365 34287 14399
rect 35170 14365 35204 14399
rect 36280 14365 36314 14399
rect 37197 14365 37231 14399
rect 37309 14365 37343 14399
rect 38292 14365 38326 14399
rect 40233 14365 40267 14399
rect 40325 14365 40359 14399
rect 40417 14365 40451 14399
rect 41245 14365 41279 14399
rect 41337 14365 41371 14399
rect 42073 14365 42107 14399
rect 42221 14365 42255 14399
rect 42538 14365 42572 14399
rect 43269 14365 43303 14399
rect 44005 14365 44039 14399
rect 44189 14365 44223 14399
rect 44281 14365 44315 14399
rect 44373 14365 44407 14399
rect 45385 14365 45419 14399
rect 47225 14365 47259 14399
rect 57989 14365 58023 14399
rect 1869 14297 1903 14331
rect 18889 14297 18923 14331
rect 19686 14297 19720 14331
rect 30012 14297 30046 14331
rect 31830 14297 31864 14331
rect 36645 14297 36679 14331
rect 40555 14297 40589 14331
rect 42349 14297 42383 14331
rect 42441 14297 42475 14331
rect 45652 14297 45686 14331
rect 47492 14297 47526 14331
rect 15853 14229 15887 14263
rect 22937 14229 22971 14263
rect 26525 14229 26559 14263
rect 35173 14229 35207 14263
rect 36369 14229 36403 14263
rect 36461 14229 36495 14263
rect 39405 14229 39439 14263
rect 41521 14229 41555 14263
rect 43453 14229 43487 14263
rect 44557 14229 44591 14263
rect 58081 14229 58115 14263
rect 2421 14025 2455 14059
rect 11161 14025 11195 14059
rect 16221 14025 16255 14059
rect 28365 14025 28399 14059
rect 31309 14025 31343 14059
rect 36369 14025 36403 14059
rect 37657 14025 37691 14059
rect 41889 14025 41923 14059
rect 43453 14025 43487 14059
rect 44741 14025 44775 14059
rect 47225 14025 47259 14059
rect 48145 14025 48179 14059
rect 10701 13957 10735 13991
rect 22744 13957 22778 13991
rect 30196 13957 30230 13991
rect 39120 13957 39154 13991
rect 41613 13957 41647 13991
rect 46857 13957 46891 13991
rect 1593 13889 1627 13923
rect 10057 13889 10091 13923
rect 12265 13889 12299 13923
rect 12449 13889 12483 13923
rect 13185 13889 13219 13923
rect 14013 13889 14047 13923
rect 16865 13889 16899 13923
rect 19165 13889 19199 13923
rect 24317 13889 24351 13923
rect 27169 13889 27203 13923
rect 29929 13889 29963 13923
rect 32873 13889 32907 13923
rect 33149 13889 33183 13923
rect 35245 13889 35279 13923
rect 37565 13889 37599 13923
rect 38853 13889 38887 13923
rect 41337 13889 41371 13923
rect 41521 13889 41555 13923
rect 41705 13889 41739 13923
rect 43361 13889 43395 13923
rect 43545 13889 43579 13923
rect 44543 13889 44577 13923
rect 46673 13889 46707 13923
rect 46949 13889 46983 13923
rect 47041 13889 47075 13923
rect 47961 13889 47995 13923
rect 1777 13821 1811 13855
rect 9873 13821 9907 13855
rect 11989 13821 12023 13855
rect 12173 13821 12207 13855
rect 12357 13821 12391 13855
rect 13277 13821 13311 13855
rect 17141 13821 17175 13855
rect 21465 13821 21499 13855
rect 22477 13821 22511 13855
rect 34253 13821 34287 13855
rect 34989 13821 35023 13855
rect 44373 13821 44407 13855
rect 47777 13821 47811 13855
rect 10977 13753 11011 13787
rect 13553 13753 13587 13787
rect 40233 13753 40267 13787
rect 10241 13685 10275 13719
rect 18429 13685 18463 13719
rect 23857 13685 23891 13719
rect 25513 13685 25547 13719
rect 11253 13481 11287 13515
rect 37473 13481 37507 13515
rect 38117 13481 38151 13515
rect 10609 13413 10643 13447
rect 16037 13413 16071 13447
rect 22937 13413 22971 13447
rect 29745 13413 29779 13447
rect 36553 13413 36587 13447
rect 12265 13345 12299 13379
rect 13553 13345 13587 13379
rect 13645 13345 13679 13379
rect 19441 13345 19475 13379
rect 27629 13345 27663 13379
rect 30297 13345 30331 13379
rect 35173 13345 35207 13379
rect 58173 13345 58207 13379
rect 1593 13277 1627 13311
rect 10609 13277 10643 13311
rect 10793 13277 10827 13311
rect 11437 13277 11471 13311
rect 11713 13277 11747 13311
rect 12357 13277 12391 13311
rect 13369 13277 13403 13311
rect 13461 13277 13495 13311
rect 14381 13277 14415 13311
rect 14657 13277 14691 13311
rect 14749 13277 14783 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 15761 13277 15795 13311
rect 15905 13277 15939 13311
rect 16589 13277 16623 13311
rect 18889 13277 18923 13311
rect 21741 13277 21775 13311
rect 24593 13277 24627 13311
rect 26525 13277 26559 13311
rect 30113 13277 30147 13311
rect 31217 13277 31251 13311
rect 33609 13277 33643 13311
rect 37105 13277 37139 13311
rect 37289 13277 37323 13311
rect 37933 13277 37967 13311
rect 38761 13277 38795 13311
rect 39129 13277 39163 13311
rect 40049 13277 40083 13311
rect 40325 13277 40359 13311
rect 40417 13277 40451 13311
rect 41061 13277 41095 13311
rect 41245 13277 41279 13311
rect 41337 13277 41371 13311
rect 41521 13277 41555 13311
rect 41613 13277 41647 13311
rect 42073 13277 42107 13311
rect 42165 13277 42199 13311
rect 57897 13277 57931 13311
rect 1869 13209 1903 13243
rect 19686 13209 19720 13243
rect 24838 13209 24872 13243
rect 32965 13209 32999 13243
rect 33425 13209 33459 13243
rect 35418 13209 35452 13243
rect 40233 13209 40267 13243
rect 57069 13209 57103 13243
rect 2329 13141 2363 13175
rect 11621 13141 11655 13175
rect 12725 13141 12759 13175
rect 13185 13141 13219 13175
rect 14565 13141 14599 13175
rect 14933 13141 14967 13175
rect 20821 13141 20855 13175
rect 25973 13141 26007 13175
rect 30205 13141 30239 13175
rect 33701 13141 33735 13175
rect 40601 13141 40635 13175
rect 57161 13141 57195 13175
rect 11161 12937 11195 12971
rect 12541 12937 12575 12971
rect 17877 12937 17911 12971
rect 25237 12937 25271 12971
rect 27721 12937 27755 12971
rect 10149 12869 10183 12903
rect 17785 12869 17819 12903
rect 22284 12869 22318 12903
rect 27445 12869 27479 12903
rect 32505 12869 32539 12903
rect 32597 12869 32631 12903
rect 36461 12869 36495 12903
rect 40969 12869 41003 12903
rect 42993 12869 43027 12903
rect 10057 12801 10091 12835
rect 10241 12801 10275 12835
rect 13185 12801 13219 12835
rect 14013 12801 14047 12835
rect 16957 12801 16991 12835
rect 17141 12801 17175 12835
rect 17953 12801 17987 12835
rect 19165 12801 19199 12835
rect 24041 12801 24075 12835
rect 27169 12801 27203 12835
rect 27353 12801 27387 12835
rect 27583 12801 27617 12835
rect 28181 12801 28215 12835
rect 31309 12801 31343 12835
rect 32321 12801 32355 12835
rect 32689 12801 32723 12835
rect 33885 12801 33919 12835
rect 36093 12801 36127 12835
rect 39681 12801 39715 12835
rect 39865 12801 39899 12835
rect 40693 12801 40727 12835
rect 40877 12801 40911 12835
rect 41061 12801 41095 12835
rect 41889 12801 41923 12835
rect 10701 12733 10735 12767
rect 12081 12733 12115 12767
rect 13277 12733 13311 12767
rect 15117 12733 15151 12767
rect 17049 12733 17083 12767
rect 17601 12733 17635 12767
rect 18337 12733 18371 12767
rect 22017 12733 22051 12767
rect 31401 12733 31435 12767
rect 31493 12733 31527 12767
rect 34161 12733 34195 12767
rect 37473 12733 37507 12767
rect 37749 12733 37783 12767
rect 38945 12733 38979 12767
rect 41705 12733 41739 12767
rect 43085 12733 43119 12767
rect 43177 12733 43211 12767
rect 10977 12665 11011 12699
rect 12357 12665 12391 12699
rect 29377 12665 29411 12699
rect 30941 12665 30975 12699
rect 32873 12665 32907 12699
rect 41245 12665 41279 12699
rect 13461 12597 13495 12631
rect 20361 12597 20395 12631
rect 23397 12597 23431 12631
rect 35449 12597 35483 12631
rect 39957 12597 39991 12631
rect 42073 12597 42107 12631
rect 42625 12597 42659 12631
rect 12633 12393 12667 12427
rect 14381 12393 14415 12427
rect 16037 12393 16071 12427
rect 18797 12393 18831 12427
rect 33149 12393 33183 12427
rect 39129 12393 39163 12427
rect 43085 12393 43119 12427
rect 22937 12325 22971 12359
rect 37565 12325 37599 12359
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 11805 12257 11839 12291
rect 14565 12257 14599 12291
rect 14749 12257 14783 12291
rect 14841 12257 14875 12291
rect 15393 12257 15427 12291
rect 15853 12257 15887 12291
rect 25697 12257 25731 12291
rect 30297 12257 30331 12291
rect 33701 12257 33735 12291
rect 35633 12257 35667 12291
rect 36185 12257 36219 12291
rect 36553 12257 36587 12291
rect 38025 12257 38059 12291
rect 38209 12257 38243 12291
rect 41521 12257 41555 12291
rect 1593 12189 1627 12223
rect 1869 12189 1903 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 13277 12189 13311 12223
rect 14657 12189 14691 12223
rect 16589 12189 16623 12223
rect 19441 12189 19475 12223
rect 21741 12189 21775 12223
rect 24593 12189 24627 12223
rect 27721 12189 27755 12223
rect 30941 12189 30975 12223
rect 31217 12189 31251 12223
rect 33517 12189 33551 12223
rect 35234 12189 35268 12223
rect 35725 12189 35759 12223
rect 36369 12189 36403 12223
rect 37933 12189 37967 12223
rect 38853 12189 38887 12223
rect 38945 12189 38979 12223
rect 40233 12189 40267 12223
rect 41797 12189 41831 12223
rect 57897 12189 57931 12223
rect 12449 12121 12483 12155
rect 12649 12121 12683 12155
rect 13553 12121 13587 12155
rect 15669 12121 15703 12155
rect 19708 12121 19742 12155
rect 27988 12121 28022 12155
rect 30113 12121 30147 12155
rect 33609 12121 33643 12155
rect 40049 12121 40083 12155
rect 58173 12121 58207 12155
rect 12817 12053 12851 12087
rect 15761 12053 15795 12087
rect 20821 12053 20855 12087
rect 29101 12053 29135 12087
rect 29745 12053 29779 12087
rect 30205 12053 30239 12087
rect 32505 12053 32539 12087
rect 35081 12053 35115 12087
rect 35265 12053 35299 12087
rect 40325 12053 40359 12087
rect 15301 11849 15335 11883
rect 17049 11849 17083 11883
rect 20361 11849 20395 11883
rect 23397 11849 23431 11883
rect 25513 11849 25547 11883
rect 27813 11849 27847 11883
rect 33609 11849 33643 11883
rect 34069 11849 34103 11883
rect 39957 11849 39991 11883
rect 41521 11849 41555 11883
rect 44005 11849 44039 11883
rect 15761 11781 15795 11815
rect 28641 11781 28675 11815
rect 32413 11781 32447 11815
rect 35725 11781 35759 11815
rect 36553 11781 36587 11815
rect 36645 11781 36679 11815
rect 41245 11781 41279 11815
rect 42892 11781 42926 11815
rect 1593 11713 1627 11747
rect 11989 11713 12023 11747
rect 12909 11713 12943 11747
rect 13829 11713 13863 11747
rect 14933 11713 14967 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 16313 11713 16347 11747
rect 16990 11713 17024 11747
rect 17969 11713 18003 11747
rect 18245 11713 18279 11747
rect 19165 11713 19199 11747
rect 22017 11713 22051 11747
rect 22273 11713 22307 11747
rect 24317 11713 24351 11747
rect 31217 11713 31251 11747
rect 33425 11713 33459 11747
rect 34437 11713 34471 11747
rect 35357 11713 35391 11747
rect 36369 11713 36403 11747
rect 36737 11713 36771 11747
rect 37729 11713 37763 11747
rect 39313 11713 39347 11747
rect 39497 11713 39531 11747
rect 40141 11713 40175 11747
rect 40233 11713 40267 11747
rect 40417 11713 40451 11747
rect 40509 11713 40543 11747
rect 40969 11713 41003 11747
rect 41153 11713 41187 11747
rect 41337 11713 41371 11747
rect 42625 11713 42659 11747
rect 58081 11713 58115 11747
rect 1777 11645 1811 11679
rect 11713 11645 11747 11679
rect 11897 11645 11931 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 13001 11645 13035 11679
rect 15025 11645 15059 11679
rect 17509 11645 17543 11679
rect 18429 11645 18463 11679
rect 27905 11645 27939 11679
rect 28089 11645 28123 11679
rect 31309 11645 31343 11679
rect 31401 11645 31435 11679
rect 33241 11645 33275 11679
rect 34529 11645 34563 11679
rect 34713 11645 34747 11679
rect 37473 11645 37507 11679
rect 39405 11645 39439 11679
rect 14197 11577 14231 11611
rect 14289 11577 14323 11611
rect 16865 11577 16899 11611
rect 18061 11577 18095 11611
rect 30113 11577 30147 11611
rect 12909 11509 12943 11543
rect 13277 11509 13311 11543
rect 16221 11509 16255 11543
rect 17417 11509 17451 11543
rect 27445 11509 27479 11543
rect 30849 11509 30883 11543
rect 32689 11509 32723 11543
rect 36921 11509 36955 11543
rect 38853 11509 38887 11543
rect 58265 11509 58299 11543
rect 13645 11305 13679 11339
rect 14749 11305 14783 11339
rect 18889 11305 18923 11339
rect 25973 11305 26007 11339
rect 37381 11305 37415 11339
rect 39037 11305 39071 11339
rect 12633 11237 12667 11271
rect 13461 11237 13495 11271
rect 27629 11237 27663 11271
rect 33609 11237 33643 11271
rect 34253 11237 34287 11271
rect 36461 11237 36495 11271
rect 40969 11237 41003 11271
rect 14933 11169 14967 11203
rect 15025 11169 15059 11203
rect 15209 11169 15243 11203
rect 18521 11169 18555 11203
rect 34897 11169 34931 11203
rect 37013 11169 37047 11203
rect 38209 11169 38243 11203
rect 38669 11169 38703 11203
rect 1593 11101 1627 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 15117 11101 15151 11135
rect 15761 11101 15795 11135
rect 18705 11101 18739 11135
rect 20085 11101 20119 11135
rect 20545 11101 20579 11135
rect 20821 11101 20855 11135
rect 21189 11101 21223 11135
rect 21281 11101 21315 11135
rect 21741 11101 21775 11135
rect 24593 11101 24627 11135
rect 26433 11101 26467 11135
rect 30297 11101 30331 11135
rect 32229 11101 32263 11135
rect 32485 11101 32519 11135
rect 34069 11101 34103 11135
rect 35173 11101 35207 11135
rect 37197 11101 37231 11135
rect 37841 11101 37875 11135
rect 38025 11101 38059 11135
rect 38853 11101 38887 11135
rect 40417 11101 40451 11135
rect 40785 11101 40819 11135
rect 41705 11101 41739 11135
rect 43913 11101 43947 11135
rect 44097 11101 44131 11135
rect 44281 11101 44315 11135
rect 52653 11101 52687 11135
rect 52837 11101 52871 11135
rect 53021 11101 53055 11135
rect 57897 11101 57931 11135
rect 1869 11033 1903 11067
rect 13185 11033 13219 11067
rect 24860 11033 24894 11067
rect 30564 11033 30598 11067
rect 40601 11033 40635 11067
rect 40693 11033 40727 11067
rect 43453 11033 43487 11067
rect 52925 11033 52959 11067
rect 58173 11033 58207 11067
rect 16957 10965 16991 10999
rect 22937 10965 22971 10999
rect 31677 10965 31711 10999
rect 53205 10965 53239 10999
rect 14289 10761 14323 10795
rect 15117 10761 15151 10795
rect 24961 10761 24995 10795
rect 29101 10761 29135 10795
rect 30849 10761 30883 10795
rect 31217 10761 31251 10795
rect 31309 10761 31343 10795
rect 32137 10761 32171 10795
rect 37841 10761 37875 10795
rect 50721 10761 50755 10795
rect 13369 10693 13403 10727
rect 13921 10693 13955 10727
rect 14121 10693 14155 10727
rect 33149 10693 33183 10727
rect 33885 10693 33919 10727
rect 41521 10693 41555 10727
rect 43085 10693 43119 10727
rect 44189 10693 44223 10727
rect 49433 10693 49467 10727
rect 1593 10625 1627 10659
rect 13277 10625 13311 10659
rect 13461 10625 13495 10659
rect 14749 10625 14783 10659
rect 14933 10625 14967 10659
rect 15071 10625 15105 10659
rect 15301 10625 15335 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 16865 10625 16899 10659
rect 16957 10625 16991 10659
rect 18075 10625 18109 10659
rect 18521 10625 18555 10659
rect 19165 10625 19199 10659
rect 22201 10625 22235 10659
rect 23765 10625 23799 10659
rect 27261 10625 27295 10659
rect 27905 10625 27939 10659
rect 32505 10625 32539 10659
rect 32597 10625 32631 10659
rect 33701 10625 33735 10659
rect 33977 10625 34011 10659
rect 34345 10625 34379 10659
rect 34437 10625 34471 10659
rect 34713 10625 34747 10659
rect 36001 10625 36035 10659
rect 36277 10625 36311 10659
rect 38669 10625 38703 10659
rect 38853 10625 38887 10659
rect 39497 10625 39531 10659
rect 39681 10625 39715 10659
rect 40601 10625 40635 10659
rect 40693 10625 40727 10659
rect 40877 10625 40911 10659
rect 40969 10625 41003 10659
rect 42993 10625 43027 10659
rect 57253 10625 57287 10659
rect 57437 10625 57471 10659
rect 1777 10557 1811 10591
rect 18245 10557 18279 10591
rect 18613 10557 18647 10591
rect 22569 10557 22603 10591
rect 31493 10557 31527 10591
rect 32689 10557 32723 10591
rect 34621 10557 34655 10591
rect 34989 10557 35023 10591
rect 35357 10557 35391 10591
rect 36093 10557 36127 10591
rect 37933 10557 37967 10591
rect 38117 10557 38151 10591
rect 43269 10557 43303 10591
rect 35725 10489 35759 10523
rect 38945 10489 38979 10523
rect 14105 10421 14139 10455
rect 16313 10421 16347 10455
rect 17601 10421 17635 10455
rect 20361 10421 20395 10455
rect 27353 10421 27387 10455
rect 33517 10421 33551 10455
rect 36277 10421 36311 10455
rect 36461 10421 36495 10455
rect 37473 10421 37507 10455
rect 39497 10421 39531 10455
rect 40417 10421 40451 10455
rect 41797 10421 41831 10455
rect 42625 10421 42659 10455
rect 45477 10421 45511 10455
rect 57345 10421 57379 10455
rect 11805 10217 11839 10251
rect 14473 10217 14507 10251
rect 24685 10217 24719 10251
rect 29009 10217 29043 10251
rect 34069 10217 34103 10251
rect 35449 10217 35483 10251
rect 58265 10217 58299 10251
rect 11621 10149 11655 10183
rect 36553 10149 36587 10183
rect 11345 10081 11379 10115
rect 15117 10081 15151 10115
rect 15485 10081 15519 10115
rect 17049 10081 17083 10115
rect 17693 10081 17727 10115
rect 18245 10081 18279 10115
rect 18613 10081 18647 10115
rect 23213 10081 23247 10115
rect 23765 10081 23799 10115
rect 25145 10081 25179 10115
rect 25789 10081 25823 10115
rect 30205 10081 30239 10115
rect 30297 10081 30331 10115
rect 41429 10081 41463 10115
rect 43085 10081 43119 10115
rect 44189 10081 44223 10115
rect 56885 10081 56919 10115
rect 14473 10013 14507 10047
rect 14657 10013 14691 10047
rect 15301 10013 15335 10047
rect 16129 10013 16163 10047
rect 16241 10013 16275 10047
rect 16957 10013 16991 10047
rect 17233 10013 17267 10047
rect 18153 10013 18187 10047
rect 18429 10013 18463 10047
rect 19717 10013 19751 10047
rect 19868 10013 19902 10047
rect 19993 10013 20027 10047
rect 20085 10013 20119 10047
rect 20821 10013 20855 10047
rect 21189 10013 21223 10047
rect 21373 10013 21407 10047
rect 22109 10013 22143 10047
rect 23305 10013 23339 10047
rect 23673 10013 23707 10047
rect 27629 10013 27663 10047
rect 30113 10013 30147 10047
rect 31309 10013 31343 10047
rect 34069 10013 34103 10047
rect 34345 10013 34379 10047
rect 34897 10013 34931 10047
rect 35081 10013 35115 10047
rect 35173 10013 35207 10047
rect 35265 10013 35299 10047
rect 36001 10013 36035 10047
rect 36185 10013 36219 10047
rect 36277 10013 36311 10047
rect 36369 10013 36403 10047
rect 37105 10013 37139 10047
rect 37372 10013 37406 10047
rect 40325 10013 40359 10047
rect 40473 10013 40507 10047
rect 40693 10013 40727 10047
rect 40790 10013 40824 10047
rect 41705 10013 41739 10047
rect 43913 10013 43947 10047
rect 15945 9945 15979 9979
rect 16331 9945 16365 9979
rect 16497 9945 16531 9979
rect 22661 9945 22695 9979
rect 25237 9945 25271 9979
rect 26056 9945 26090 9979
rect 27896 9945 27930 9979
rect 38945 9945 38979 9979
rect 39129 9945 39163 9979
rect 39313 9945 39347 9979
rect 40601 9945 40635 9979
rect 57130 9945 57164 9979
rect 19533 9877 19567 9911
rect 20637 9877 20671 9911
rect 25145 9877 25179 9911
rect 27169 9877 27203 9911
rect 29745 9877 29779 9911
rect 32505 9877 32539 9911
rect 34253 9877 34287 9911
rect 38485 9877 38519 9911
rect 40969 9877 41003 9911
rect 24409 9673 24443 9707
rect 29009 9673 29043 9707
rect 30573 9673 30607 9707
rect 31585 9673 31619 9707
rect 32321 9673 32355 9707
rect 32689 9673 32723 9707
rect 40325 9673 40359 9707
rect 44005 9673 44039 9707
rect 56977 9673 57011 9707
rect 58265 9673 58299 9707
rect 19165 9605 19199 9639
rect 21005 9605 21039 9639
rect 25145 9605 25179 9639
rect 29377 9605 29411 9639
rect 29469 9605 29503 9639
rect 30757 9605 30791 9639
rect 31401 9605 31435 9639
rect 33977 9605 34011 9639
rect 35909 9605 35943 9639
rect 40049 9605 40083 9639
rect 42892 9605 42926 9639
rect 44925 9605 44959 9639
rect 1593 9537 1627 9571
rect 11713 9537 11747 9571
rect 14565 9537 14599 9571
rect 15209 9537 15243 9571
rect 16865 9537 16899 9571
rect 17785 9537 17819 9571
rect 17877 9537 17911 9571
rect 18061 9537 18095 9571
rect 18153 9537 18187 9571
rect 18705 9537 18739 9571
rect 19901 9537 19935 9571
rect 20269 9537 20303 9571
rect 20637 9537 20671 9571
rect 21465 9537 21499 9571
rect 22201 9537 22235 9571
rect 23857 9537 23891 9571
rect 24501 9537 24535 9571
rect 24593 9537 24627 9571
rect 25605 9537 25639 9571
rect 25789 9537 25823 9571
rect 25973 9537 26007 9571
rect 27169 9537 27203 9571
rect 30205 9537 30239 9571
rect 30389 9537 30423 9571
rect 30527 9537 30561 9571
rect 31217 9537 31251 9571
rect 31539 9537 31573 9571
rect 31767 9537 31801 9571
rect 32505 9537 32539 9571
rect 32781 9537 32815 9571
rect 33701 9537 33735 9571
rect 33885 9537 33919 9571
rect 34069 9537 34103 9571
rect 34805 9537 34839 9571
rect 35725 9537 35759 9571
rect 35993 9537 36027 9571
rect 36093 9537 36127 9571
rect 36737 9537 36771 9571
rect 36921 9537 36955 9571
rect 37841 9537 37875 9571
rect 38393 9537 38427 9571
rect 38945 9537 38979 9571
rect 39129 9537 39163 9571
rect 39221 9537 39255 9571
rect 39681 9537 39715 9571
rect 39774 9537 39808 9571
rect 39957 9537 39991 9571
rect 40187 9537 40221 9571
rect 41429 9537 41463 9571
rect 41797 9537 41831 9571
rect 42625 9537 42659 9571
rect 56793 9537 56827 9571
rect 57069 9537 57103 9571
rect 58081 9537 58115 9571
rect 1777 9469 1811 9503
rect 12173 9469 12207 9503
rect 14657 9469 14691 9503
rect 15853 9469 15887 9503
rect 16313 9469 16347 9503
rect 16957 9469 16991 9503
rect 23213 9469 23247 9503
rect 24041 9469 24075 9503
rect 26433 9469 26467 9503
rect 26525 9469 26559 9503
rect 28365 9469 28399 9503
rect 29561 9469 29595 9503
rect 41521 9469 41555 9503
rect 41889 9469 41923 9503
rect 45017 9469 45051 9503
rect 45109 9469 45143 9503
rect 11989 9401 12023 9435
rect 16129 9401 16163 9435
rect 36737 9401 36771 9435
rect 56793 9401 56827 9435
rect 15301 9333 15335 9367
rect 17601 9333 17635 9367
rect 34253 9333 34287 9367
rect 34989 9333 35023 9367
rect 36277 9333 36311 9367
rect 38945 9333 38979 9367
rect 40877 9333 40911 9367
rect 44557 9333 44591 9367
rect 17417 9129 17451 9163
rect 20085 9129 20119 9163
rect 24593 9129 24627 9163
rect 26617 9129 26651 9163
rect 28457 9129 28491 9163
rect 29009 9129 29043 9163
rect 38669 9129 38703 9163
rect 16405 9061 16439 9095
rect 32137 9061 32171 9095
rect 44005 9061 44039 9095
rect 23857 8993 23891 9027
rect 25237 8993 25271 9027
rect 32965 8993 32999 9027
rect 34161 8993 34195 9027
rect 35909 8993 35943 9027
rect 41061 8993 41095 9027
rect 1593 8925 1627 8959
rect 15669 8925 15703 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 17049 8925 17083 8959
rect 17509 8925 17543 8959
rect 18521 8925 18555 8959
rect 18609 8925 18643 8959
rect 19441 8925 19475 8959
rect 19589 8925 19623 8959
rect 19809 8925 19843 8959
rect 19947 8925 19981 8959
rect 20545 8925 20579 8959
rect 22937 8925 22971 8959
rect 23305 8925 23339 8959
rect 24593 8925 24627 8959
rect 24777 8925 24811 8959
rect 27077 8925 27111 8959
rect 29009 8925 29043 8959
rect 29193 8925 29227 8959
rect 29745 8925 29779 8959
rect 29837 8925 29871 8959
rect 30757 8925 30791 8959
rect 31033 8925 31067 8959
rect 33149 8925 33183 8959
rect 33885 8925 33919 8959
rect 34897 8925 34931 8959
rect 35173 8925 35207 8959
rect 36185 8925 36219 8959
rect 38025 8925 38059 8959
rect 38118 8925 38152 8959
rect 38393 8925 38427 8959
rect 38490 8925 38524 8959
rect 39497 8925 39531 8959
rect 40049 8925 40083 8959
rect 40245 8925 40279 8959
rect 40785 8925 40819 8959
rect 42625 8925 42659 8959
rect 42892 8925 42926 8959
rect 57069 8925 57103 8959
rect 57253 8925 57287 8959
rect 57897 8925 57931 8959
rect 1869 8857 1903 8891
rect 18061 8857 18095 8891
rect 18153 8857 18187 8891
rect 18705 8857 18739 8891
rect 19717 8857 19751 8891
rect 22845 8857 22879 8891
rect 23397 8857 23431 8891
rect 25504 8857 25538 8891
rect 27344 8857 27378 8891
rect 30297 8857 30331 8891
rect 33425 8857 33459 8891
rect 37565 8857 37599 8891
rect 38301 8857 38335 8891
rect 39129 8857 39163 8891
rect 39313 8857 39347 8891
rect 40141 8857 40175 8891
rect 58173 8857 58207 8891
rect 15761 8789 15795 8823
rect 20361 8789 20395 8823
rect 21833 8789 21867 8823
rect 33333 8789 33367 8823
rect 57161 8789 57195 8823
rect 16221 8585 16255 8619
rect 18705 8585 18739 8619
rect 21465 8585 21499 8619
rect 27537 8585 27571 8619
rect 28365 8585 28399 8619
rect 28733 8585 28767 8619
rect 33241 8585 33275 8619
rect 35725 8585 35759 8619
rect 39405 8585 39439 8619
rect 41245 8585 41279 8619
rect 17325 8517 17359 8551
rect 18521 8517 18555 8551
rect 25145 8517 25179 8551
rect 27629 8517 27663 8551
rect 32597 8517 32631 8551
rect 33517 8517 33551 8551
rect 38270 8517 38304 8551
rect 40417 8517 40451 8551
rect 1593 8449 1627 8483
rect 10425 8449 10459 8483
rect 16037 8449 16071 8483
rect 17049 8449 17083 8483
rect 18153 8449 18187 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 19993 8449 20027 8483
rect 20269 8449 20303 8483
rect 20453 8449 20487 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 22109 8449 22143 8483
rect 23765 8449 23799 8483
rect 25605 8449 25639 8483
rect 25973 8449 26007 8483
rect 26065 8449 26099 8483
rect 28825 8449 28859 8483
rect 29837 8449 29871 8483
rect 30104 8449 30138 8483
rect 32229 8449 32263 8483
rect 33701 8449 33735 8483
rect 33793 8449 33827 8483
rect 34437 8449 34471 8483
rect 34529 8449 34563 8483
rect 34653 8449 34687 8483
rect 35633 8449 35667 8483
rect 36277 8449 36311 8483
rect 36425 8449 36459 8483
rect 36553 8449 36587 8483
rect 36645 8449 36679 8483
rect 36742 8449 36776 8483
rect 38025 8449 38059 8483
rect 40049 8449 40083 8483
rect 40142 8449 40176 8483
rect 40325 8449 40359 8483
rect 40514 8449 40548 8483
rect 41429 8449 41463 8483
rect 41521 8449 41555 8483
rect 41705 8449 41739 8483
rect 41797 8449 41831 8483
rect 42717 8449 42751 8483
rect 43637 8449 43671 8483
rect 44557 8449 44591 8483
rect 57161 8449 57195 8483
rect 1777 8381 1811 8415
rect 10149 8381 10183 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 10609 8381 10643 8415
rect 22845 8381 22879 8415
rect 24501 8381 24535 8415
rect 27813 8381 27847 8415
rect 28917 8381 28951 8415
rect 34897 8381 34931 8415
rect 42993 8381 43027 8415
rect 43821 8381 43855 8415
rect 44741 8381 44775 8415
rect 27169 8313 27203 8347
rect 33977 8313 34011 8347
rect 40693 8313 40727 8347
rect 57345 8313 57379 8347
rect 18521 8245 18555 8279
rect 19257 8245 19291 8279
rect 31217 8245 31251 8279
rect 33517 8245 33551 8279
rect 34345 8245 34379 8279
rect 36921 8245 36955 8279
rect 10241 8041 10275 8075
rect 16589 8041 16623 8075
rect 17141 8041 17175 8075
rect 27721 8041 27755 8075
rect 29837 8041 29871 8075
rect 39129 8041 39163 8075
rect 40785 8041 40819 8075
rect 58265 8041 58299 8075
rect 10149 7973 10183 8007
rect 36185 7973 36219 8007
rect 56149 7973 56183 8007
rect 17417 7905 17451 7939
rect 17509 7905 17543 7939
rect 17601 7905 17635 7939
rect 19717 7905 19751 7939
rect 21005 7905 21039 7939
rect 21097 7905 21131 7939
rect 22017 7905 22051 7939
rect 22845 7905 22879 7939
rect 25145 7905 25179 7939
rect 25881 7905 25915 7939
rect 28273 7905 28307 7939
rect 32965 7905 32999 7939
rect 34069 7905 34103 7939
rect 36645 7905 36679 7939
rect 36829 7905 36863 7939
rect 56885 7905 56919 7939
rect 1593 7837 1627 7871
rect 16497 7837 16531 7871
rect 17325 7837 17359 7871
rect 18153 7837 18187 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18567 7837 18601 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 21465 7837 21499 7871
rect 22477 7837 22511 7871
rect 24685 7837 24719 7871
rect 28181 7837 28215 7871
rect 29009 7837 29043 7871
rect 30021 7837 30055 7871
rect 30113 7837 30147 7871
rect 30297 7837 30331 7871
rect 30389 7837 30423 7871
rect 33609 7837 33643 7871
rect 33701 7837 33735 7871
rect 33885 7837 33919 7871
rect 35081 7837 35115 7871
rect 35229 7837 35263 7871
rect 35449 7837 35483 7871
rect 35546 7837 35580 7871
rect 37473 7837 37507 7871
rect 38577 7837 38611 7871
rect 38761 7837 38795 7871
rect 38945 7837 38979 7871
rect 40037 7837 40071 7871
rect 40233 7837 40267 7871
rect 40693 7837 40727 7871
rect 41935 7837 41969 7871
rect 42070 7837 42104 7871
rect 42170 7837 42204 7871
rect 42349 7837 42383 7871
rect 42809 7837 42843 7871
rect 56425 7837 56459 7871
rect 57141 7837 57175 7871
rect 1869 7769 1903 7803
rect 9781 7769 9815 7803
rect 19625 7769 19659 7803
rect 20269 7769 20303 7803
rect 21557 7769 21591 7803
rect 26126 7769 26160 7803
rect 31217 7769 31251 7803
rect 35357 7769 35391 7803
rect 36553 7769 36587 7803
rect 37841 7769 37875 7803
rect 38853 7769 38887 7803
rect 43054 7769 43088 7803
rect 56149 7769 56183 7803
rect 56333 7769 56367 7803
rect 18705 7701 18739 7735
rect 27261 7701 27295 7735
rect 28089 7701 28123 7735
rect 29101 7701 29135 7735
rect 35725 7701 35759 7735
rect 40141 7701 40175 7735
rect 41705 7701 41739 7735
rect 44189 7701 44223 7735
rect 9597 7497 9631 7531
rect 23305 7497 23339 7531
rect 25881 7497 25915 7531
rect 26249 7497 26283 7531
rect 31125 7497 31159 7531
rect 31309 7497 31343 7531
rect 32689 7497 32723 7531
rect 34069 7497 34103 7531
rect 41705 7497 41739 7531
rect 42717 7497 42751 7531
rect 44465 7497 44499 7531
rect 8677 7429 8711 7463
rect 9689 7429 9723 7463
rect 26341 7429 26375 7463
rect 28641 7429 28675 7463
rect 35449 7429 35483 7463
rect 38945 7429 38979 7463
rect 56333 7429 56367 7463
rect 56517 7429 56551 7463
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 9413 7361 9447 7395
rect 10333 7361 10367 7395
rect 10425 7361 10459 7395
rect 17049 7361 17083 7395
rect 17325 7361 17359 7395
rect 17877 7361 17911 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 19717 7361 19751 7395
rect 20821 7361 20855 7395
rect 20913 7361 20947 7395
rect 22017 7361 22051 7395
rect 24685 7361 24719 7395
rect 27169 7361 27203 7395
rect 31306 7361 31340 7395
rect 31769 7361 31803 7395
rect 35081 7361 35115 7395
rect 35174 7361 35208 7395
rect 35357 7361 35391 7395
rect 35546 7361 35580 7395
rect 36173 7367 36207 7401
rect 36461 7361 36495 7395
rect 37473 7361 37507 7395
rect 37657 7361 37691 7395
rect 37933 7361 37967 7395
rect 38117 7361 38151 7395
rect 38761 7361 38795 7395
rect 41613 7361 41647 7395
rect 41797 7361 41831 7395
rect 42625 7361 42659 7395
rect 42809 7361 42843 7395
rect 43361 7361 43395 7395
rect 44649 7361 44683 7395
rect 44833 7361 44867 7395
rect 44925 7361 44959 7395
rect 56609 7361 56643 7395
rect 57069 7361 57103 7395
rect 58081 7361 58115 7395
rect 58265 7361 58299 7395
rect 7941 7293 7975 7327
rect 10149 7293 10183 7327
rect 10517 7293 10551 7327
rect 10609 7293 10643 7327
rect 17141 7293 17175 7327
rect 18153 7293 18187 7327
rect 18981 7293 19015 7327
rect 19165 7293 19199 7327
rect 20361 7293 20395 7327
rect 20453 7293 20487 7327
rect 21373 7293 21407 7327
rect 25053 7293 25087 7327
rect 25421 7293 25455 7327
rect 26525 7293 26559 7327
rect 27537 7293 27571 7327
rect 32781 7293 32815 7327
rect 32873 7293 32907 7327
rect 33885 7293 33919 7327
rect 34345 7293 34379 7327
rect 34437 7293 34471 7327
rect 36645 7293 36679 7327
rect 37841 7293 37875 7327
rect 38577 7293 38611 7327
rect 41981 7293 42015 7327
rect 43637 7293 43671 7327
rect 57345 7293 57379 7327
rect 27445 7225 27479 7259
rect 35725 7225 35759 7259
rect 36277 7225 36311 7259
rect 37749 7225 37783 7259
rect 41429 7225 41463 7259
rect 58173 7225 58207 7259
rect 9229 7157 9263 7191
rect 17233 7157 17267 7191
rect 24850 7157 24884 7191
rect 24961 7157 24995 7191
rect 27307 7157 27341 7191
rect 27813 7157 27847 7191
rect 29929 7157 29963 7191
rect 31677 7157 31711 7191
rect 32321 7157 32355 7191
rect 56333 7157 56367 7191
rect 10885 6953 10919 6987
rect 17601 6953 17635 6987
rect 18889 6953 18923 6987
rect 24593 6953 24627 6987
rect 38301 6953 38335 6987
rect 42809 6953 42843 6987
rect 58265 6953 58299 6987
rect 36461 6885 36495 6919
rect 9689 6817 9723 6851
rect 9965 6817 9999 6851
rect 18245 6817 18279 6851
rect 18613 6817 18647 6851
rect 21741 6817 21775 6851
rect 25605 6817 25639 6851
rect 30389 6817 30423 6851
rect 30481 6817 30515 6851
rect 32413 6817 32447 6851
rect 35474 6817 35508 6851
rect 37933 6817 37967 6851
rect 40141 6817 40175 6851
rect 42073 6817 42107 6851
rect 44005 6817 44039 6851
rect 56885 6817 56919 6851
rect 1593 6749 1627 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10701 6749 10735 6783
rect 16313 6749 16347 6783
rect 17417 6749 17451 6783
rect 17601 6749 17635 6783
rect 18521 6749 18555 6783
rect 19809 6749 19843 6783
rect 20177 6749 20211 6783
rect 20453 6749 20487 6783
rect 20821 6749 20855 6783
rect 21189 6749 21223 6783
rect 22017 6749 22051 6783
rect 22293 6749 22327 6783
rect 22477 6749 22511 6783
rect 22753 6749 22787 6783
rect 23673 6749 23707 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 24777 6749 24811 6783
rect 24869 6749 24903 6783
rect 25053 6749 25087 6783
rect 25145 6749 25179 6783
rect 27445 6749 27479 6783
rect 31125 6749 31159 6783
rect 31493 6749 31527 6783
rect 32597 6749 32631 6783
rect 32689 6749 32723 6783
rect 32873 6749 32907 6783
rect 32965 6749 32999 6783
rect 33425 6749 33459 6783
rect 33573 6749 33607 6783
rect 33793 6749 33827 6783
rect 33931 6749 33965 6783
rect 34897 6749 34931 6783
rect 35375 6749 35409 6783
rect 36185 6749 36219 6783
rect 37197 6749 37231 6783
rect 37381 6749 37415 6783
rect 37473 6727 37507 6761
rect 38117 6749 38151 6783
rect 40049 6749 40083 6783
rect 40969 6749 41003 6783
rect 41153 6749 41187 6783
rect 41797 6749 41831 6783
rect 42985 6749 43019 6783
rect 43117 6749 43151 6783
rect 43269 6749 43303 6783
rect 43361 6749 43395 6783
rect 43821 6749 43855 6783
rect 57141 6749 57175 6783
rect 1869 6681 1903 6715
rect 18730 6681 18764 6715
rect 25872 6681 25906 6715
rect 27712 6681 27746 6715
rect 31309 6681 31343 6715
rect 31401 6681 31435 6715
rect 33701 6681 33735 6715
rect 41337 6681 41371 6715
rect 17785 6613 17819 6647
rect 23121 6613 23155 6647
rect 26985 6613 27019 6647
rect 28825 6613 28859 6647
rect 29929 6613 29963 6647
rect 30297 6613 30331 6647
rect 31677 6613 31711 6647
rect 34069 6613 34103 6647
rect 35081 6613 35115 6647
rect 37013 6613 37047 6647
rect 10149 6409 10183 6443
rect 17325 6409 17359 6443
rect 21189 6409 21223 6443
rect 27537 6409 27571 6443
rect 27997 6409 28031 6443
rect 28365 6409 28399 6443
rect 39497 6409 39531 6443
rect 9689 6341 9723 6375
rect 28457 6341 28491 6375
rect 29285 6341 29319 6375
rect 34253 6341 34287 6375
rect 35265 6341 35299 6375
rect 35357 6341 35391 6375
rect 37740 6341 37774 6375
rect 44097 6341 44131 6375
rect 55781 6341 55815 6375
rect 55965 6341 55999 6375
rect 1593 6273 1627 6307
rect 10885 6273 10919 6307
rect 11713 6273 11747 6307
rect 16865 6273 16899 6307
rect 18889 6273 18923 6307
rect 19993 6273 20027 6307
rect 20269 6273 20303 6307
rect 20729 6273 20763 6307
rect 21373 6273 21407 6307
rect 22017 6273 22051 6307
rect 22293 6273 22327 6307
rect 22753 6273 22787 6307
rect 23213 6273 23247 6307
rect 24961 6273 24995 6307
rect 25513 6273 25547 6307
rect 27353 6273 27387 6307
rect 29469 6273 29503 6307
rect 29561 6273 29595 6307
rect 29745 6273 29779 6307
rect 29837 6273 29871 6307
rect 30297 6273 30331 6307
rect 31401 6273 31435 6307
rect 32321 6273 32355 6307
rect 32588 6273 32622 6307
rect 34437 6273 34471 6307
rect 34529 6273 34563 6307
rect 34989 6273 35023 6307
rect 35127 6273 35161 6307
rect 35495 6273 35529 6307
rect 36369 6273 36403 6307
rect 36553 6273 36587 6307
rect 37473 6273 37507 6307
rect 39313 6273 39347 6307
rect 42901 6273 42935 6307
rect 43545 6273 43579 6307
rect 43637 6273 43671 6307
rect 56057 6273 56091 6307
rect 56609 6273 56643 6307
rect 58081 6273 58115 6307
rect 1777 6205 1811 6239
rect 19165 6205 19199 6239
rect 25789 6205 25823 6239
rect 27169 6205 27203 6239
rect 28641 6205 28675 6239
rect 30573 6205 30607 6239
rect 36093 6205 36127 6239
rect 56885 6205 56919 6239
rect 9965 6137 9999 6171
rect 11069 6137 11103 6171
rect 17141 6137 17175 6171
rect 22109 6137 22143 6171
rect 30849 6137 30883 6171
rect 33701 6137 33735 6171
rect 34253 6137 34287 6171
rect 36369 6137 36403 6171
rect 58265 6137 58299 6171
rect 11897 6069 11931 6103
rect 16313 6069 16347 6103
rect 18429 6069 18463 6103
rect 30665 6069 30699 6103
rect 31493 6069 31527 6103
rect 35633 6069 35667 6103
rect 38853 6069 38887 6103
rect 55781 6069 55815 6103
rect 13277 5865 13311 5899
rect 24593 5865 24627 5899
rect 30297 5865 30331 5899
rect 37749 5865 37783 5899
rect 41705 5865 41739 5899
rect 44557 5865 44591 5899
rect 45293 5865 45327 5899
rect 24041 5797 24075 5831
rect 26617 5797 26651 5831
rect 32045 5797 32079 5831
rect 33517 5797 33551 5831
rect 10885 5729 10919 5763
rect 19901 5729 19935 5763
rect 19993 5729 20027 5763
rect 20913 5729 20947 5763
rect 22845 5729 22879 5763
rect 25237 5729 25271 5763
rect 27169 5729 27203 5763
rect 30941 5729 30975 5763
rect 32689 5729 32723 5763
rect 36001 5729 36035 5763
rect 36829 5729 36863 5763
rect 38209 5729 38243 5763
rect 38393 5729 38427 5763
rect 43177 5729 43211 5763
rect 56885 5729 56919 5763
rect 1593 5661 1627 5695
rect 14749 5661 14783 5695
rect 16405 5661 16439 5695
rect 17049 5661 17083 5695
rect 17509 5661 17543 5695
rect 18429 5661 18463 5695
rect 20361 5661 20395 5695
rect 21833 5661 21867 5695
rect 23673 5661 23707 5695
rect 24593 5661 24627 5695
rect 24777 5661 24811 5695
rect 29009 5661 29043 5695
rect 29193 5661 29227 5695
rect 33241 5661 33275 5695
rect 35081 5661 35115 5695
rect 36185 5661 36219 5695
rect 37013 5661 37047 5695
rect 42441 5661 42475 5695
rect 42717 5661 42751 5695
rect 45201 5661 45235 5695
rect 57141 5661 57175 5695
rect 1869 5593 1903 5627
rect 10701 5593 10735 5627
rect 11621 5593 11655 5627
rect 12357 5593 12391 5627
rect 12541 5593 12575 5627
rect 13185 5593 13219 5627
rect 15025 5593 15059 5627
rect 17785 5593 17819 5627
rect 18705 5593 18739 5627
rect 20453 5593 20487 5627
rect 23857 5593 23891 5627
rect 25482 5593 25516 5627
rect 27436 5593 27470 5627
rect 30757 5593 30791 5627
rect 34161 5593 34195 5627
rect 35357 5593 35391 5627
rect 39037 5593 39071 5627
rect 41613 5593 41647 5627
rect 42625 5593 42659 5627
rect 43729 5593 43763 5627
rect 44465 5593 44499 5627
rect 11713 5525 11747 5559
rect 28549 5525 28583 5559
rect 29101 5525 29135 5559
rect 30665 5525 30699 5559
rect 32413 5525 32447 5559
rect 32505 5525 32539 5559
rect 33701 5525 33735 5559
rect 36369 5525 36403 5559
rect 37197 5525 37231 5559
rect 38117 5525 38151 5559
rect 39129 5525 39163 5559
rect 43821 5525 43855 5559
rect 58265 5525 58299 5559
rect 9597 5321 9631 5355
rect 23949 5321 23983 5355
rect 27721 5321 27755 5355
rect 28089 5321 28123 5355
rect 29009 5321 29043 5355
rect 40601 5321 40635 5355
rect 43545 5321 43579 5355
rect 45017 5321 45051 5355
rect 57253 5321 57287 5355
rect 11161 5253 11195 5287
rect 15853 5253 15887 5287
rect 18521 5253 18555 5287
rect 25390 5253 25424 5287
rect 34437 5253 34471 5287
rect 36369 5253 36403 5287
rect 37565 5253 37599 5287
rect 39037 5253 39071 5287
rect 39957 5253 39991 5287
rect 41245 5253 41279 5287
rect 41429 5253 41463 5287
rect 1593 5185 1627 5219
rect 8769 5185 8803 5219
rect 9781 5185 9815 5219
rect 9873 5185 9907 5219
rect 10057 5185 10091 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 13369 5185 13403 5219
rect 14013 5185 14047 5219
rect 16957 5185 16991 5219
rect 17049 5185 17083 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 19441 5185 19475 5219
rect 19717 5185 19751 5219
rect 20453 5185 20487 5219
rect 22201 5185 22235 5219
rect 22845 5185 22879 5219
rect 24317 5185 24351 5219
rect 25145 5185 25179 5219
rect 28917 5185 28951 5219
rect 29101 5185 29135 5219
rect 29561 5185 29595 5219
rect 29828 5185 29862 5219
rect 31585 5185 31619 5219
rect 32321 5185 32355 5219
rect 33517 5185 33551 5219
rect 33701 5185 33735 5219
rect 34161 5185 34195 5219
rect 35081 5185 35115 5219
rect 36185 5185 36219 5219
rect 38301 5185 38335 5219
rect 39773 5185 39807 5219
rect 40509 5185 40543 5219
rect 42717 5185 42751 5219
rect 43361 5185 43395 5219
rect 44833 5185 44867 5219
rect 45661 5185 45695 5219
rect 46581 5185 46615 5219
rect 57161 5185 57195 5219
rect 57345 5185 57379 5219
rect 58081 5185 58115 5219
rect 1777 5117 1811 5151
rect 9965 5117 9999 5151
rect 14749 5117 14783 5151
rect 16313 5117 16347 5151
rect 18981 5117 19015 5151
rect 21005 5117 21039 5151
rect 24409 5117 24443 5151
rect 24593 5117 24627 5151
rect 28181 5117 28215 5151
rect 28365 5117 28399 5151
rect 31401 5117 31435 5151
rect 32413 5117 32447 5151
rect 35357 5117 35391 5151
rect 36001 5117 36035 5151
rect 38485 5117 38519 5151
rect 44649 5117 44683 5151
rect 46765 5117 46799 5151
rect 12633 5049 12667 5083
rect 13553 5049 13587 5083
rect 15025 5049 15059 5083
rect 16129 5049 16163 5083
rect 18797 5049 18831 5083
rect 31769 5049 31803 5083
rect 33517 5049 33551 5083
rect 58265 5049 58299 5083
rect 8861 4981 8895 5015
rect 12817 4981 12851 5015
rect 14197 4981 14231 5015
rect 15209 4981 15243 5015
rect 26525 4981 26559 5015
rect 30941 4981 30975 5015
rect 32413 4981 32447 5015
rect 32689 4981 32723 5015
rect 33241 4981 33275 5015
rect 37657 4981 37691 5015
rect 39129 4981 39163 5015
rect 42809 4981 42843 5015
rect 45753 4981 45787 5015
rect 9229 4777 9263 4811
rect 10701 4777 10735 4811
rect 13645 4777 13679 4811
rect 26525 4777 26559 4811
rect 28549 4777 28583 4811
rect 29837 4777 29871 4811
rect 32413 4777 32447 4811
rect 34989 4777 35023 4811
rect 37841 4777 37875 4811
rect 40969 4777 41003 4811
rect 42993 4777 43027 4811
rect 54217 4777 54251 4811
rect 57345 4777 57379 4811
rect 7021 4709 7055 4743
rect 8585 4709 8619 4743
rect 10517 4709 10551 4743
rect 11713 4709 11747 4743
rect 11805 4709 11839 4743
rect 12541 4709 12575 4743
rect 13461 4709 13495 4743
rect 15025 4709 15059 4743
rect 15209 4709 15243 4743
rect 22109 4709 22143 4743
rect 38853 4709 38887 4743
rect 40325 4709 40359 4743
rect 44097 4709 44131 4743
rect 9597 4641 9631 4675
rect 10241 4641 10275 4675
rect 11345 4641 11379 4675
rect 12265 4641 12299 4675
rect 21281 4641 21315 4675
rect 22753 4641 22787 4675
rect 23949 4641 23983 4675
rect 25145 4641 25179 4675
rect 27445 4641 27479 4675
rect 27537 4641 27571 4675
rect 30297 4641 30331 4675
rect 30481 4641 30515 4675
rect 35541 4641 35575 4675
rect 46121 4641 46155 4675
rect 58173 4641 58207 4675
rect 9413 4573 9447 4607
rect 9505 4573 9539 4607
rect 9689 4573 9723 4607
rect 15669 4573 15703 4607
rect 16589 4573 16623 4607
rect 17509 4573 17543 4607
rect 18429 4573 18463 4607
rect 19533 4573 19567 4607
rect 20913 4573 20947 4607
rect 22017 4573 22051 4607
rect 22293 4573 22327 4607
rect 27353 4573 27387 4607
rect 28457 4573 28491 4607
rect 28825 4573 28859 4607
rect 30205 4573 30239 4607
rect 31033 4573 31067 4607
rect 33609 4573 33643 4607
rect 34069 4573 34103 4607
rect 36185 4573 36219 4607
rect 37197 4573 37231 4607
rect 38025 4573 38059 4607
rect 38117 4573 38151 4607
rect 40785 4573 40819 4607
rect 41613 4573 41647 4607
rect 42349 4573 42383 4607
rect 42497 4573 42531 4607
rect 42814 4573 42848 4607
rect 43545 4573 43579 4607
rect 43821 4573 43855 4607
rect 43913 4573 43947 4607
rect 57897 4573 57931 4607
rect 6837 4505 6871 4539
rect 7665 4505 7699 4539
rect 8401 4505 8435 4539
rect 13185 4505 13219 4539
rect 14749 4505 14783 4539
rect 15945 4505 15979 4539
rect 16865 4505 16899 4539
rect 17785 4505 17819 4539
rect 18705 4505 18739 4539
rect 19809 4505 19843 4539
rect 23673 4505 23707 4539
rect 25390 4505 25424 4539
rect 31300 4505 31334 4539
rect 32965 4505 32999 4539
rect 33149 4505 33183 4539
rect 34345 4505 34379 4539
rect 36461 4505 36495 4539
rect 37841 4505 37875 4539
rect 38669 4505 38703 4539
rect 40141 4505 40175 4539
rect 42625 4505 42659 4539
rect 42717 4505 42751 4539
rect 43729 4505 43763 4539
rect 45293 4505 45327 4539
rect 46366 4505 46400 4539
rect 54125 4505 54159 4539
rect 57253 4505 57287 4539
rect 7757 4437 7791 4471
rect 12725 4437 12759 4471
rect 23305 4437 23339 4471
rect 23765 4437 23799 4471
rect 26985 4437 27019 4471
rect 29009 4437 29043 4471
rect 35357 4437 35391 4471
rect 35449 4437 35483 4471
rect 37289 4437 37323 4471
rect 41705 4437 41739 4471
rect 45385 4437 45419 4471
rect 47501 4437 47535 4471
rect 13277 4233 13311 4267
rect 19717 4233 19751 4267
rect 20729 4233 20763 4267
rect 20821 4233 20855 4267
rect 23313 4233 23347 4267
rect 23949 4233 23983 4267
rect 29561 4233 29595 4267
rect 31769 4233 31803 4267
rect 32321 4233 32355 4267
rect 32689 4233 32723 4267
rect 35633 4233 35667 4267
rect 39497 4233 39531 4267
rect 45937 4233 45971 4267
rect 54585 4233 54619 4267
rect 2881 4165 2915 4199
rect 3617 4165 3651 4199
rect 4353 4165 4387 4199
rect 5825 4165 5859 4199
rect 7113 4165 7147 4199
rect 16129 4165 16163 4199
rect 16957 4165 16991 4199
rect 19827 4165 19861 4199
rect 19993 4165 20027 4199
rect 20453 4165 20487 4199
rect 22937 4165 22971 4199
rect 24317 4165 24351 4199
rect 27537 4165 27571 4199
rect 37565 4165 37599 4199
rect 38669 4165 38703 4199
rect 40141 4165 40175 4199
rect 41613 4165 41647 4199
rect 45109 4165 45143 4199
rect 45845 4165 45879 4199
rect 49157 4165 49191 4199
rect 50721 4165 50755 4199
rect 51549 4165 51583 4199
rect 53021 4165 53055 4199
rect 53757 4165 53791 4199
rect 58173 4165 58207 4199
rect 1593 4097 1627 4131
rect 3801 4097 3835 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 10333 4097 10367 4131
rect 12173 4097 12207 4131
rect 13185 4097 13219 4131
rect 14013 4097 14047 4131
rect 14933 4097 14967 4131
rect 15853 4097 15887 4131
rect 18521 4097 18555 4131
rect 19628 4097 19662 4131
rect 20637 4097 20671 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 22753 4097 22787 4131
rect 23029 4097 23063 4131
rect 23173 4097 23207 4131
rect 25145 4097 25179 4131
rect 25412 4097 25446 4131
rect 28549 4097 28583 4131
rect 30645 4097 30679 4131
rect 32781 4097 32815 4131
rect 33609 4097 33643 4131
rect 36461 4097 36495 4131
rect 39313 4097 39347 4131
rect 40877 4097 40911 4131
rect 42625 4097 42659 4131
rect 43269 4097 43303 4131
rect 43637 4097 43671 4131
rect 44373 4097 44407 4131
rect 46581 4097 46615 4131
rect 46765 4097 46799 4131
rect 48237 4097 48271 4131
rect 48421 4097 48455 4131
rect 49341 4097 49375 4131
rect 50905 4097 50939 4131
rect 51733 4097 51767 4131
rect 53205 4097 53239 4131
rect 53941 4097 53975 4131
rect 54401 4097 54435 4131
rect 55137 4097 55171 4131
rect 57253 4097 57287 4131
rect 58357 4097 58391 4131
rect 1777 4029 1811 4063
rect 7757 4029 7791 4063
rect 8677 4029 8711 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 12633 4029 12667 4063
rect 14289 4029 14323 4063
rect 15209 4029 15243 4063
rect 17601 4029 17635 4063
rect 18705 4029 18739 4063
rect 19441 4029 19475 4063
rect 24409 4029 24443 4063
rect 24593 4029 24627 4063
rect 27629 4029 27663 4063
rect 27721 4029 27755 4063
rect 28365 4029 28399 4063
rect 29653 4029 29687 4063
rect 29745 4029 29779 4063
rect 30389 4029 30423 4063
rect 32873 4029 32907 4063
rect 33885 4029 33919 4063
rect 35725 4029 35759 4063
rect 35817 4029 35851 4063
rect 36645 4029 36679 4063
rect 40325 4029 40359 4063
rect 41061 4029 41095 4063
rect 43361 4029 43395 4063
rect 43545 4029 43579 4063
rect 45293 4029 45327 4063
rect 57069 4029 57103 4063
rect 3065 3961 3099 3995
rect 6009 3961 6043 3995
rect 8033 3961 8067 3995
rect 8217 3961 8251 3995
rect 10701 3961 10735 3995
rect 12541 3961 12575 3995
rect 17877 3961 17911 3995
rect 55321 3961 55355 3995
rect 4445 3893 4479 3927
rect 7205 3893 7239 3927
rect 9873 3893 9907 3927
rect 10793 3893 10827 3927
rect 18061 3893 18095 3927
rect 22201 3893 22235 3927
rect 26525 3893 26559 3927
rect 27169 3893 27203 3927
rect 28733 3893 28767 3927
rect 29193 3893 29227 3927
rect 35265 3893 35299 3927
rect 37657 3893 37691 3927
rect 38761 3893 38795 3927
rect 41705 3893 41739 3927
rect 44465 3893 44499 3927
rect 48605 3893 48639 3927
rect 57437 3893 57471 3927
rect 16037 3689 16071 3723
rect 22937 3689 22971 3723
rect 24041 3689 24075 3723
rect 24593 3689 24627 3723
rect 36277 3689 36311 3723
rect 38945 3689 38979 3723
rect 41981 3689 42015 3723
rect 45385 3689 45419 3723
rect 46121 3689 46155 3723
rect 47869 3689 47903 3723
rect 48605 3689 48639 3723
rect 49341 3689 49375 3723
rect 50537 3689 50571 3723
rect 52009 3689 52043 3723
rect 54217 3689 54251 3723
rect 5457 3621 5491 3655
rect 8401 3621 8435 3655
rect 9689 3621 9723 3655
rect 11529 3621 11563 3655
rect 11713 3621 11747 3655
rect 19441 3621 19475 3655
rect 33425 3621 33459 3655
rect 37381 3621 37415 3655
rect 44005 3621 44039 3655
rect 47041 3621 47075 3655
rect 52837 3621 52871 3655
rect 58265 3621 58299 3655
rect 4721 3553 4755 3587
rect 6929 3553 6963 3587
rect 10609 3553 10643 3587
rect 12633 3553 12667 3587
rect 17785 3553 17819 3587
rect 22845 3553 22879 3587
rect 23673 3553 23707 3587
rect 25145 3553 25179 3587
rect 25789 3553 25823 3587
rect 27997 3553 28031 3587
rect 29745 3553 29779 3587
rect 34897 3553 34931 3587
rect 40325 3553 40359 3587
rect 40785 3553 40819 3587
rect 51365 3553 51399 3587
rect 56885 3553 56919 3587
rect 1593 3485 1627 3519
rect 3249 3485 3283 3519
rect 3433 3485 3467 3519
rect 5273 3485 5307 3519
rect 7481 3485 7515 3519
rect 10333 3485 10367 3519
rect 11253 3485 11287 3519
rect 12357 3485 12391 3519
rect 13277 3485 13311 3519
rect 14749 3485 14783 3519
rect 15025 3485 15059 3519
rect 16589 3485 16623 3519
rect 17509 3485 17543 3519
rect 18429 3485 18463 3519
rect 18705 3485 18739 3519
rect 19625 3485 19659 3519
rect 20637 3485 20671 3519
rect 20821 3485 20855 3519
rect 21833 3485 21867 3519
rect 22661 3485 22695 3519
rect 22937 3485 22971 3519
rect 23857 3485 23891 3519
rect 26056 3485 26090 3519
rect 27721 3485 27755 3519
rect 29049 3485 29083 3519
rect 32045 3485 32079 3519
rect 33885 3485 33919 3519
rect 35164 3485 35198 3519
rect 36737 3485 36771 3519
rect 36885 3485 36919 3519
rect 37243 3485 37277 3519
rect 37841 3485 37875 3519
rect 40693 3485 40727 3519
rect 41061 3485 41095 3519
rect 41153 3485 41187 3519
rect 42165 3485 42199 3519
rect 42349 3485 42383 3519
rect 42717 3485 42751 3519
rect 42809 3485 42843 3519
rect 43361 3485 43395 3519
rect 43509 3485 43543 3519
rect 43826 3485 43860 3519
rect 46029 3485 46063 3519
rect 48513 3485 48547 3519
rect 51181 3485 51215 3519
rect 51917 3485 51951 3519
rect 53389 3485 53423 3519
rect 55965 3485 55999 3519
rect 1869 3417 1903 3451
rect 4537 3417 4571 3451
rect 6009 3417 6043 3451
rect 6745 3417 6779 3451
rect 8125 3417 8159 3451
rect 9413 3417 9447 3451
rect 13553 3417 13587 3451
rect 15761 3417 15795 3451
rect 16865 3417 16899 3451
rect 19993 3417 20027 3451
rect 21189 3417 21223 3451
rect 21649 3417 21683 3451
rect 22035 3417 22069 3451
rect 22201 3417 22235 3451
rect 25053 3417 25087 3451
rect 28825 3417 28859 3451
rect 29193 3417 29227 3451
rect 30012 3417 30046 3451
rect 32312 3417 32346 3451
rect 34161 3417 34195 3451
rect 37013 3417 37047 3451
rect 37105 3417 37139 3451
rect 38117 3417 38151 3451
rect 38853 3417 38887 3451
rect 43637 3417 43671 3451
rect 43729 3417 43763 3451
rect 45293 3417 45327 3451
rect 46857 3417 46891 3451
rect 47777 3417 47811 3451
rect 49249 3417 49283 3451
rect 50445 3417 50479 3451
rect 52653 3417 52687 3451
rect 54125 3417 54159 3451
rect 56241 3417 56275 3451
rect 57130 3417 57164 3451
rect 6101 3349 6135 3383
rect 7573 3349 7607 3383
rect 8585 3349 8619 3383
rect 9873 3349 9907 3383
rect 19717 3349 19751 3383
rect 19809 3349 19843 3383
rect 20361 3349 20395 3383
rect 20913 3349 20947 3383
rect 21005 3349 21039 3383
rect 21925 3349 21959 3383
rect 23121 3349 23155 3383
rect 24961 3349 24995 3383
rect 27169 3349 27203 3383
rect 28733 3349 28767 3383
rect 28917 3349 28951 3383
rect 31125 3349 31159 3383
rect 53481 3349 53515 3383
rect 2973 3145 3007 3179
rect 4445 3145 4479 3179
rect 8401 3145 8435 3179
rect 20913 3145 20947 3179
rect 23029 3145 23063 3179
rect 23121 3145 23155 3179
rect 24409 3145 24443 3179
rect 25145 3145 25179 3179
rect 25513 3145 25547 3179
rect 28733 3145 28767 3179
rect 29929 3145 29963 3179
rect 30297 3145 30331 3179
rect 36277 3145 36311 3179
rect 39497 3145 39531 3179
rect 40601 3145 40635 3179
rect 44465 3145 44499 3179
rect 45201 3145 45235 3179
rect 46397 3145 46431 3179
rect 47961 3145 47995 3179
rect 49801 3145 49835 3179
rect 51273 3145 51307 3179
rect 53849 3145 53883 3179
rect 54769 3145 54803 3179
rect 58265 3145 58299 3179
rect 5089 3077 5123 3111
rect 7297 3077 7331 3111
rect 7481 3077 7515 3111
rect 7941 3077 7975 3111
rect 9137 3077 9171 3111
rect 10057 3077 10091 3111
rect 15025 3077 15059 3111
rect 19073 3077 19107 3111
rect 21189 3077 21223 3111
rect 22109 3077 22143 3111
rect 26433 3077 26467 3111
rect 27721 3077 27755 3111
rect 28549 3077 28583 3111
rect 28917 3077 28951 3111
rect 33517 3077 33551 3111
rect 35164 3077 35198 3111
rect 38669 3077 38703 3111
rect 41245 3077 41279 3111
rect 41429 3077 41463 3111
rect 42625 3077 42659 3111
rect 49709 3077 49743 3111
rect 51917 3077 51951 3111
rect 53021 3077 53055 3111
rect 55781 3077 55815 3111
rect 58173 3077 58207 3111
rect 1593 3009 1627 3043
rect 2881 3009 2915 3043
rect 3617 3009 3651 3043
rect 4353 3009 4387 3043
rect 5827 3009 5861 3043
rect 8861 3009 8895 3043
rect 9781 3009 9815 3043
rect 10701 3009 10735 3043
rect 12173 3009 12207 3043
rect 12449 3009 12483 3043
rect 13093 3009 13127 3043
rect 14013 3009 14047 3043
rect 14749 3009 14783 3043
rect 15853 3009 15887 3043
rect 17141 3009 17175 3043
rect 18797 3009 18831 3043
rect 19717 3009 19751 3043
rect 20637 3009 20671 3043
rect 20821 3009 20855 3043
rect 21045 3009 21079 3043
rect 22937 3009 22971 3043
rect 23305 3009 23339 3043
rect 24317 3009 24351 3043
rect 27445 3009 27479 3043
rect 28687 3009 28721 3043
rect 31309 3009 31343 3043
rect 32321 3009 32355 3043
rect 33241 3009 33275 3043
rect 34253 3009 34287 3043
rect 34437 3009 34471 3043
rect 34897 3009 34931 3043
rect 37473 3009 37507 3043
rect 38393 3009 38427 3043
rect 39405 3009 39439 3043
rect 40325 3009 40359 3043
rect 43269 3009 43303 3043
rect 43637 3009 43671 3043
rect 43821 3009 43855 3043
rect 44281 3009 44315 3043
rect 45109 3009 45143 3043
rect 46305 3009 46339 3043
rect 47869 3009 47903 3043
rect 48789 3009 48823 3043
rect 50445 3009 50479 3043
rect 51089 3009 51123 3043
rect 53757 3009 53791 3043
rect 54677 3009 54711 3043
rect 55505 3009 55539 3043
rect 56425 3009 56459 3043
rect 1777 2941 1811 2975
rect 10977 2941 11011 2975
rect 13369 2941 13403 2975
rect 14289 2941 14323 2975
rect 16129 2941 16163 2975
rect 17417 2941 17451 2975
rect 18337 2941 18371 2975
rect 19993 2941 20027 2975
rect 24593 2941 24627 2975
rect 25605 2941 25639 2975
rect 25789 2941 25823 2975
rect 30389 2941 30423 2975
rect 30573 2941 30607 2975
rect 31493 2941 31527 2975
rect 32505 2941 32539 2975
rect 37657 2941 37691 2975
rect 43361 2941 43395 2975
rect 53205 2941 53239 2975
rect 56609 2941 56643 2975
rect 8217 2873 8251 2907
rect 15577 2873 15611 2907
rect 22293 2873 22327 2907
rect 22753 2873 22787 2907
rect 23949 2873 23983 2907
rect 28365 2873 28399 2907
rect 52101 2873 52135 2907
rect 3709 2805 3743 2839
rect 5181 2805 5215 2839
rect 5917 2805 5951 2839
rect 49065 2805 49099 2839
rect 50537 2805 50571 2839
rect 8585 2601 8619 2635
rect 14657 2601 14691 2635
rect 25145 2601 25179 2635
rect 34161 2601 34195 2635
rect 40233 2601 40267 2635
rect 41337 2601 41371 2635
rect 42809 2601 42843 2635
rect 45845 2601 45879 2635
rect 46949 2601 46983 2635
rect 47961 2601 47995 2635
rect 49065 2601 49099 2635
rect 50537 2601 50571 2635
rect 54033 2601 54067 2635
rect 58265 2601 58299 2635
rect 4537 2533 4571 2567
rect 7665 2533 7699 2567
rect 8493 2533 8527 2567
rect 11897 2533 11931 2567
rect 22017 2533 22051 2567
rect 23029 2533 23063 2567
rect 6009 2465 6043 2499
rect 10057 2465 10091 2499
rect 14105 2465 14139 2499
rect 25697 2465 25731 2499
rect 29009 2465 29043 2499
rect 36093 2465 36127 2499
rect 52101 2465 52135 2499
rect 55689 2465 55723 2499
rect 1593 2397 1627 2431
rect 3249 2397 3283 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 10701 2397 10735 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 19993 2397 20027 2431
rect 20913 2397 20947 2431
rect 21097 2397 21131 2431
rect 22313 2397 22347 2431
rect 22569 2397 22603 2431
rect 23213 2397 23247 2431
rect 23351 2397 23385 2431
rect 27445 2397 27479 2431
rect 28733 2397 28767 2431
rect 30113 2397 30147 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 34161 2397 34195 2431
rect 34345 2397 34379 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 37473 2397 37507 2431
rect 38393 2397 38427 2431
rect 42625 2397 42659 2431
rect 44189 2397 44223 2431
rect 47869 2397 47903 2431
rect 50353 2397 50387 2431
rect 51917 2397 51951 2431
rect 55505 2397 55539 2431
rect 56425 2397 56459 2431
rect 58173 2397 58207 2431
rect 1869 2329 1903 2363
rect 4353 2329 4387 2363
rect 5089 2329 5123 2363
rect 5825 2329 5859 2363
rect 6745 2329 6779 2363
rect 6929 2329 6963 2363
rect 7481 2329 7515 2363
rect 8125 2329 8159 2363
rect 10977 2329 11011 2363
rect 12633 2329 12667 2363
rect 13553 2329 13587 2363
rect 15209 2329 15243 2363
rect 16129 2329 16163 2363
rect 17785 2329 17819 2363
rect 18705 2329 18739 2363
rect 20269 2329 20303 2363
rect 21465 2329 21499 2363
rect 22201 2329 22235 2363
rect 23581 2329 23615 2363
rect 26433 2329 26467 2363
rect 27721 2329 27755 2363
rect 30389 2329 30423 2363
rect 31309 2329 31343 2363
rect 32597 2329 32631 2363
rect 33517 2329 33551 2363
rect 35173 2329 35207 2363
rect 37749 2329 37783 2363
rect 38669 2329 38703 2363
rect 40141 2329 40175 2363
rect 41061 2329 41095 2363
rect 43453 2329 43487 2363
rect 44373 2329 44407 2363
rect 45753 2329 45787 2363
rect 46673 2329 46707 2363
rect 48789 2329 48823 2363
rect 51181 2329 51215 2363
rect 53021 2329 53055 2363
rect 53941 2329 53975 2363
rect 56701 2329 56735 2363
rect 3341 2261 3375 2295
rect 5181 2261 5215 2295
rect 16865 2261 16899 2295
rect 21189 2261 21223 2295
rect 21281 2261 21315 2295
rect 22385 2261 22419 2295
rect 23397 2261 23431 2295
rect 25513 2261 25547 2295
rect 25605 2261 25639 2295
rect 26525 2261 26559 2295
rect 36737 2261 36771 2295
rect 43545 2261 43579 2295
rect 51273 2261 51307 2295
rect 53113 2261 53147 2295
<< metal1 >>
rect 41230 61684 41236 61736
rect 41288 61724 41294 61736
rect 51442 61724 51448 61736
rect 41288 61696 51448 61724
rect 41288 61684 41294 61696
rect 51442 61684 51448 61696
rect 51500 61684 51506 61736
rect 24946 61616 24952 61668
rect 25004 61656 25010 61668
rect 40310 61656 40316 61668
rect 25004 61628 40316 61656
rect 25004 61616 25010 61628
rect 40310 61616 40316 61628
rect 40368 61616 40374 61668
rect 40402 61616 40408 61668
rect 40460 61656 40466 61668
rect 42702 61656 42708 61668
rect 40460 61628 42708 61656
rect 40460 61616 40466 61628
rect 42702 61616 42708 61628
rect 42760 61616 42766 61668
rect 28350 61548 28356 61600
rect 28408 61588 28414 61600
rect 40678 61588 40684 61600
rect 28408 61560 40684 61588
rect 28408 61548 28414 61560
rect 40678 61548 40684 61560
rect 40736 61548 40742 61600
rect 1104 61498 58880 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 58880 61498
rect 1104 61424 58880 61446
rect 7650 61384 7656 61396
rect 2240 61356 7656 61384
rect 2240 61257 2268 61356
rect 7650 61344 7656 61356
rect 7708 61344 7714 61396
rect 11057 61387 11115 61393
rect 11057 61353 11069 61387
rect 11103 61384 11115 61387
rect 15286 61384 15292 61396
rect 11103 61356 15292 61384
rect 11103 61353 11115 61356
rect 11057 61347 11115 61353
rect 15286 61344 15292 61356
rect 15344 61344 15350 61396
rect 18049 61387 18107 61393
rect 18049 61353 18061 61387
rect 18095 61384 18107 61387
rect 22830 61384 22836 61396
rect 18095 61356 22836 61384
rect 18095 61353 18107 61356
rect 18049 61347 18107 61353
rect 22830 61344 22836 61356
rect 22888 61344 22894 61396
rect 33413 61387 33471 61393
rect 33413 61353 33425 61387
rect 33459 61384 33471 61387
rect 40402 61384 40408 61396
rect 33459 61356 40408 61384
rect 33459 61353 33471 61356
rect 33413 61347 33471 61353
rect 40402 61344 40408 61356
rect 40460 61344 40466 61396
rect 40678 61344 40684 61396
rect 40736 61384 40742 61396
rect 47949 61387 48007 61393
rect 47949 61384 47961 61387
rect 40736 61356 47961 61384
rect 40736 61344 40742 61356
rect 47949 61353 47961 61356
rect 47995 61353 48007 61387
rect 51442 61384 51448 61396
rect 51403 61356 51448 61384
rect 47949 61347 48007 61353
rect 51442 61344 51448 61356
rect 51500 61344 51506 61396
rect 6270 61276 6276 61328
rect 6328 61316 6334 61328
rect 40221 61319 40279 61325
rect 40221 61316 40233 61319
rect 6328 61288 40233 61316
rect 6328 61276 6334 61288
rect 40221 61285 40233 61288
rect 40267 61285 40279 61319
rect 40221 61279 40279 61285
rect 40310 61276 40316 61328
rect 40368 61316 40374 61328
rect 44545 61319 44603 61325
rect 44545 61316 44557 61319
rect 40368 61288 44557 61316
rect 40368 61276 40374 61288
rect 44545 61285 44557 61288
rect 44591 61285 44603 61319
rect 44545 61279 44603 61285
rect 46750 61276 46756 61328
rect 46808 61316 46814 61328
rect 48777 61319 48835 61325
rect 48777 61316 48789 61319
rect 46808 61288 48789 61316
rect 46808 61276 46814 61288
rect 48777 61285 48789 61288
rect 48823 61285 48835 61319
rect 48777 61279 48835 61285
rect 48958 61276 48964 61328
rect 49016 61316 49022 61328
rect 49016 61288 55214 61316
rect 49016 61276 49022 61288
rect 2225 61251 2283 61257
rect 2225 61217 2237 61251
rect 2271 61217 2283 61251
rect 2225 61211 2283 61217
rect 3053 61251 3111 61257
rect 3053 61217 3065 61251
rect 3099 61248 3111 61251
rect 17402 61248 17408 61260
rect 3099 61220 17408 61248
rect 3099 61217 3111 61220
rect 3053 61211 3111 61217
rect 17402 61208 17408 61220
rect 17460 61208 17466 61260
rect 20622 61208 20628 61260
rect 20680 61248 20686 61260
rect 21453 61251 21511 61257
rect 21453 61248 21465 61251
rect 20680 61220 21465 61248
rect 20680 61208 20686 61220
rect 21453 61217 21465 61220
rect 21499 61217 21511 61251
rect 21453 61211 21511 61217
rect 25501 61251 25559 61257
rect 25501 61217 25513 61251
rect 25547 61248 25559 61251
rect 28258 61248 28264 61260
rect 25547 61220 28264 61248
rect 25547 61217 25559 61220
rect 25501 61211 25559 61217
rect 28258 61208 28264 61220
rect 28316 61208 28322 61260
rect 32677 61251 32735 61257
rect 32677 61217 32689 61251
rect 32723 61248 32735 61251
rect 39574 61248 39580 61260
rect 32723 61220 39580 61248
rect 32723 61217 32735 61220
rect 32677 61211 32735 61217
rect 39574 61208 39580 61220
rect 39632 61208 39638 61260
rect 41138 61208 41144 61260
rect 41196 61248 41202 61260
rect 52273 61251 52331 61257
rect 52273 61248 52285 61251
rect 41196 61220 52285 61248
rect 41196 61208 41202 61220
rect 52273 61217 52285 61220
rect 52319 61217 52331 61251
rect 55186 61248 55214 61288
rect 56781 61251 56839 61257
rect 56781 61248 56793 61251
rect 55186 61220 56793 61248
rect 52273 61211 52331 61217
rect 56781 61217 56793 61220
rect 56827 61217 56839 61251
rect 56781 61211 56839 61217
rect 1670 61180 1676 61192
rect 1631 61152 1676 61180
rect 1670 61140 1676 61152
rect 1728 61140 1734 61192
rect 2774 61140 2780 61192
rect 2832 61180 2838 61192
rect 4706 61180 4712 61192
rect 2832 61152 2877 61180
rect 4667 61152 4712 61180
rect 2832 61140 2838 61152
rect 4706 61140 4712 61152
rect 4764 61140 4770 61192
rect 5629 61183 5687 61189
rect 5629 61149 5641 61183
rect 5675 61180 5687 61183
rect 5994 61180 6000 61192
rect 5675 61152 6000 61180
rect 5675 61149 5687 61152
rect 5629 61143 5687 61149
rect 5994 61140 6000 61152
rect 6052 61140 6058 61192
rect 6638 61180 6644 61192
rect 6599 61152 6644 61180
rect 6638 61140 6644 61152
rect 6696 61140 6702 61192
rect 7558 61180 7564 61192
rect 7519 61152 7564 61180
rect 7558 61140 7564 61152
rect 7616 61140 7622 61192
rect 9214 61180 9220 61192
rect 9175 61152 9220 61180
rect 9214 61140 9220 61152
rect 9272 61140 9278 61192
rect 10226 61180 10232 61192
rect 10187 61152 10232 61180
rect 10226 61140 10232 61152
rect 10284 61140 10290 61192
rect 10965 61183 11023 61189
rect 10965 61149 10977 61183
rect 11011 61180 11023 61183
rect 11146 61180 11152 61192
rect 11011 61152 11152 61180
rect 11011 61149 11023 61152
rect 10965 61143 11023 61149
rect 11146 61140 11152 61152
rect 11204 61140 11210 61192
rect 12066 61180 12072 61192
rect 12027 61152 12072 61180
rect 12066 61140 12072 61152
rect 12124 61140 12130 61192
rect 12802 61180 12808 61192
rect 12763 61152 12808 61180
rect 12802 61140 12808 61152
rect 12860 61140 12866 61192
rect 14918 61180 14924 61192
rect 14879 61152 14924 61180
rect 14918 61140 14924 61152
rect 14976 61140 14982 61192
rect 16114 61180 16120 61192
rect 16075 61152 16120 61180
rect 16114 61140 16120 61152
rect 16172 61140 16178 61192
rect 17126 61180 17132 61192
rect 17087 61152 17132 61180
rect 17126 61140 17132 61152
rect 17184 61140 17190 61192
rect 17954 61180 17960 61192
rect 17915 61152 17960 61180
rect 17954 61140 17960 61152
rect 18012 61140 18018 61192
rect 18690 61180 18696 61192
rect 18651 61152 18696 61180
rect 18690 61140 18696 61152
rect 18748 61140 18754 61192
rect 19794 61180 19800 61192
rect 19755 61152 19800 61180
rect 19794 61140 19800 61152
rect 19852 61140 19858 61192
rect 20533 61183 20591 61189
rect 20533 61149 20545 61183
rect 20579 61180 20591 61183
rect 20714 61180 20720 61192
rect 20579 61152 20720 61180
rect 20579 61149 20591 61152
rect 20533 61143 20591 61149
rect 20714 61140 20720 61152
rect 20772 61140 20778 61192
rect 21266 61180 21272 61192
rect 21227 61152 21272 61180
rect 21266 61140 21272 61152
rect 21324 61140 21330 61192
rect 22370 61180 22376 61192
rect 22331 61152 22376 61180
rect 22370 61140 22376 61152
rect 22428 61140 22434 61192
rect 23658 61140 23664 61192
rect 23716 61180 23722 61192
rect 23845 61183 23903 61189
rect 23845 61180 23857 61183
rect 23716 61152 23857 61180
rect 23716 61140 23722 61152
rect 23845 61149 23857 61152
rect 23891 61149 23903 61183
rect 23845 61143 23903 61149
rect 25130 61140 25136 61192
rect 25188 61180 25194 61192
rect 25225 61183 25283 61189
rect 25225 61180 25237 61183
rect 25188 61152 25237 61180
rect 25188 61140 25194 61152
rect 25225 61149 25237 61152
rect 25271 61149 25283 61183
rect 25225 61143 25283 61149
rect 25866 61140 25872 61192
rect 25924 61180 25930 61192
rect 26237 61183 26295 61189
rect 26237 61180 26249 61183
rect 25924 61152 26249 61180
rect 25924 61140 25930 61152
rect 26237 61149 26249 61152
rect 26283 61149 26295 61183
rect 26237 61143 26295 61149
rect 26602 61140 26608 61192
rect 26660 61180 26666 61192
rect 27249 61183 27307 61189
rect 27249 61180 27261 61183
rect 26660 61152 27261 61180
rect 26660 61140 26666 61152
rect 27249 61149 27261 61152
rect 27295 61149 27307 61183
rect 27249 61143 27307 61149
rect 28074 61140 28080 61192
rect 28132 61180 28138 61192
rect 28169 61183 28227 61189
rect 28169 61180 28181 61183
rect 28132 61152 28181 61180
rect 28132 61140 28138 61152
rect 28169 61149 28181 61152
rect 28215 61149 28227 61183
rect 29822 61180 29828 61192
rect 29783 61152 29828 61180
rect 28169 61143 28227 61149
rect 29822 61140 29828 61152
rect 29880 61140 29886 61192
rect 31202 61180 31208 61192
rect 31163 61152 31208 61180
rect 31202 61140 31208 61152
rect 31260 61140 31266 61192
rect 31754 61140 31760 61192
rect 31812 61180 31818 61192
rect 32401 61183 32459 61189
rect 32401 61180 32413 61183
rect 31812 61152 32413 61180
rect 31812 61140 31818 61152
rect 32401 61149 32413 61152
rect 32447 61149 32459 61183
rect 32401 61143 32459 61149
rect 32490 61140 32496 61192
rect 32548 61180 32554 61192
rect 33321 61183 33379 61189
rect 33321 61180 33333 61183
rect 32548 61152 33333 61180
rect 32548 61140 32554 61152
rect 33321 61149 33333 61152
rect 33367 61149 33379 61183
rect 33321 61143 33379 61149
rect 33502 61140 33508 61192
rect 33560 61180 33566 61192
rect 34057 61183 34115 61189
rect 34057 61180 34069 61183
rect 33560 61152 34069 61180
rect 33560 61140 33566 61152
rect 34057 61149 34069 61152
rect 34103 61149 34115 61183
rect 34057 61143 34115 61149
rect 34238 61140 34244 61192
rect 34296 61180 34302 61192
rect 34977 61183 35035 61189
rect 34977 61180 34989 61183
rect 34296 61152 34989 61180
rect 34296 61140 34302 61152
rect 34977 61149 34989 61152
rect 35023 61149 35035 61183
rect 34977 61143 35035 61149
rect 35066 61140 35072 61192
rect 35124 61180 35130 61192
rect 35124 61152 35848 61180
rect 35124 61140 35130 61152
rect 4893 61115 4951 61121
rect 4893 61081 4905 61115
rect 4939 61112 4951 61115
rect 5534 61112 5540 61124
rect 4939 61084 5540 61112
rect 4939 61081 4951 61084
rect 4893 61075 4951 61081
rect 5534 61072 5540 61084
rect 5592 61072 5598 61124
rect 6917 61115 6975 61121
rect 6917 61081 6929 61115
rect 6963 61081 6975 61115
rect 7834 61112 7840 61124
rect 7795 61084 7840 61112
rect 6917 61075 6975 61081
rect 5718 61044 5724 61056
rect 5679 61016 5724 61044
rect 5718 61004 5724 61016
rect 5776 61004 5782 61056
rect 6932 61044 6960 61075
rect 7834 61072 7840 61084
rect 7892 61072 7898 61124
rect 10502 61112 10508 61124
rect 9048 61084 10508 61112
rect 9048 61044 9076 61084
rect 10502 61072 10508 61084
rect 10560 61072 10566 61124
rect 15194 61112 15200 61124
rect 15155 61084 15200 61112
rect 15194 61072 15200 61084
rect 15252 61072 15258 61124
rect 16301 61115 16359 61121
rect 16301 61081 16313 61115
rect 16347 61112 16359 61115
rect 17494 61112 17500 61124
rect 16347 61084 17500 61112
rect 16347 61081 16359 61084
rect 16301 61075 16359 61081
rect 17494 61072 17500 61084
rect 17552 61072 17558 61124
rect 19978 61112 19984 61124
rect 19939 61084 19984 61112
rect 19978 61072 19984 61084
rect 20036 61072 20042 61124
rect 22278 61112 22284 61124
rect 21284 61084 22284 61112
rect 9306 61044 9312 61056
rect 6932 61016 9076 61044
rect 9267 61016 9312 61044
rect 9306 61004 9312 61016
rect 9364 61004 9370 61056
rect 10318 61044 10324 61056
rect 10279 61016 10324 61044
rect 10318 61004 10324 61016
rect 10376 61004 10382 61056
rect 12158 61044 12164 61056
rect 12119 61016 12164 61044
rect 12158 61004 12164 61016
rect 12216 61004 12222 61056
rect 12894 61044 12900 61056
rect 12855 61016 12900 61044
rect 12894 61004 12900 61016
rect 12952 61004 12958 61056
rect 17310 61044 17316 61056
rect 17271 61016 17316 61044
rect 17310 61004 17316 61016
rect 17368 61004 17374 61056
rect 18598 61004 18604 61056
rect 18656 61044 18662 61056
rect 18785 61047 18843 61053
rect 18785 61044 18797 61047
rect 18656 61016 18797 61044
rect 18656 61004 18662 61016
rect 18785 61013 18797 61016
rect 18831 61013 18843 61047
rect 18785 61007 18843 61013
rect 20625 61047 20683 61053
rect 20625 61013 20637 61047
rect 20671 61044 20683 61047
rect 21284 61044 21312 61084
rect 22278 61072 22284 61084
rect 22336 61072 22342 61124
rect 26421 61115 26479 61121
rect 26421 61081 26433 61115
rect 26467 61112 26479 61115
rect 26878 61112 26884 61124
rect 26467 61084 26884 61112
rect 26467 61081 26479 61084
rect 26421 61075 26479 61081
rect 26878 61072 26884 61084
rect 26936 61072 26942 61124
rect 28442 61112 28448 61124
rect 28403 61084 28448 61112
rect 28442 61072 28448 61084
rect 28500 61072 28506 61124
rect 31570 61112 31576 61124
rect 31531 61084 31576 61112
rect 31570 61072 31576 61084
rect 31628 61072 31634 61124
rect 34698 61072 34704 61124
rect 34756 61112 34762 61124
rect 35713 61115 35771 61121
rect 35713 61112 35725 61115
rect 34756 61084 35725 61112
rect 34756 61072 34762 61084
rect 35713 61081 35725 61084
rect 35759 61081 35771 61115
rect 35820 61112 35848 61152
rect 35894 61140 35900 61192
rect 35952 61180 35958 61192
rect 36449 61183 36507 61189
rect 36449 61180 36461 61183
rect 35952 61152 36461 61180
rect 35952 61140 35958 61152
rect 36449 61149 36461 61152
rect 36495 61149 36507 61183
rect 36449 61143 36507 61149
rect 36906 61140 36912 61192
rect 36964 61180 36970 61192
rect 37553 61183 37611 61189
rect 37553 61180 37565 61183
rect 36964 61152 37565 61180
rect 36964 61140 36970 61152
rect 37553 61149 37565 61152
rect 37599 61149 37611 61183
rect 37553 61143 37611 61149
rect 37642 61140 37648 61192
rect 37700 61180 37706 61192
rect 38289 61183 38347 61189
rect 38289 61180 38301 61183
rect 37700 61152 38301 61180
rect 37700 61140 37706 61152
rect 38289 61149 38301 61152
rect 38335 61149 38347 61183
rect 38289 61143 38347 61149
rect 38654 61140 38660 61192
rect 38712 61180 38718 61192
rect 38933 61183 38991 61189
rect 38933 61180 38945 61183
rect 38712 61152 38945 61180
rect 38712 61140 38718 61152
rect 38933 61149 38945 61152
rect 38979 61149 38991 61183
rect 38933 61143 38991 61149
rect 39482 61140 39488 61192
rect 39540 61180 39546 61192
rect 40037 61183 40095 61189
rect 40037 61180 40049 61183
rect 39540 61152 40049 61180
rect 39540 61140 39546 61152
rect 40037 61149 40049 61152
rect 40083 61149 40095 61183
rect 40037 61143 40095 61149
rect 40126 61140 40132 61192
rect 40184 61180 40190 61192
rect 40865 61183 40923 61189
rect 40865 61180 40877 61183
rect 40184 61152 40877 61180
rect 40184 61140 40190 61152
rect 40865 61149 40877 61152
rect 40911 61149 40923 61183
rect 40865 61143 40923 61149
rect 40954 61140 40960 61192
rect 41012 61180 41018 61192
rect 41601 61183 41659 61189
rect 41601 61180 41613 61183
rect 41012 61152 41613 61180
rect 41012 61140 41018 61152
rect 41601 61149 41613 61152
rect 41647 61149 41659 61183
rect 41601 61143 41659 61149
rect 42058 61140 42064 61192
rect 42116 61180 42122 61192
rect 42613 61183 42671 61189
rect 42613 61180 42625 61183
rect 42116 61152 42625 61180
rect 42116 61140 42122 61152
rect 42613 61149 42625 61152
rect 42659 61149 42671 61183
rect 42613 61143 42671 61149
rect 42794 61140 42800 61192
rect 42852 61180 42858 61192
rect 43533 61183 43591 61189
rect 43533 61180 43545 61183
rect 42852 61152 43545 61180
rect 42852 61140 42858 61152
rect 43533 61149 43545 61152
rect 43579 61149 43591 61183
rect 43533 61143 43591 61149
rect 43622 61140 43628 61192
rect 43680 61180 43686 61192
rect 44361 61183 44419 61189
rect 44361 61180 44373 61183
rect 43680 61152 44373 61180
rect 43680 61140 43686 61152
rect 44361 61149 44373 61152
rect 44407 61149 44419 61183
rect 44361 61143 44419 61149
rect 44542 61140 44548 61192
rect 44600 61180 44606 61192
rect 45281 61183 45339 61189
rect 45281 61180 45293 61183
rect 44600 61152 45293 61180
rect 44600 61140 44606 61152
rect 45281 61149 45293 61152
rect 45327 61149 45339 61183
rect 45281 61143 45339 61149
rect 45554 61140 45560 61192
rect 45612 61180 45618 61192
rect 46017 61183 46075 61189
rect 46017 61180 46029 61183
rect 45612 61152 46029 61180
rect 45612 61140 45618 61152
rect 46017 61149 46029 61152
rect 46063 61149 46075 61183
rect 46017 61143 46075 61149
rect 46106 61140 46112 61192
rect 46164 61180 46170 61192
rect 46753 61183 46811 61189
rect 46753 61180 46765 61183
rect 46164 61152 46765 61180
rect 46164 61140 46170 61152
rect 46753 61149 46765 61152
rect 46799 61149 46811 61183
rect 46753 61143 46811 61149
rect 47210 61140 47216 61192
rect 47268 61180 47274 61192
rect 47857 61183 47915 61189
rect 47857 61180 47869 61183
rect 47268 61152 47869 61180
rect 47268 61140 47274 61152
rect 47857 61149 47869 61152
rect 47903 61149 47915 61183
rect 47857 61143 47915 61149
rect 48314 61140 48320 61192
rect 48372 61180 48378 61192
rect 48593 61183 48651 61189
rect 48593 61180 48605 61183
rect 48372 61152 48605 61180
rect 48372 61140 48378 61152
rect 48593 61149 48605 61152
rect 48639 61149 48651 61183
rect 48593 61143 48651 61149
rect 48682 61140 48688 61192
rect 48740 61180 48746 61192
rect 49329 61183 49387 61189
rect 49329 61180 49341 61183
rect 48740 61152 49341 61180
rect 48740 61140 48746 61152
rect 49329 61149 49341 61152
rect 49375 61149 49387 61183
rect 49329 61143 49387 61149
rect 49694 61140 49700 61192
rect 49752 61180 49758 61192
rect 50433 61183 50491 61189
rect 50433 61180 50445 61183
rect 49752 61152 50445 61180
rect 49752 61140 49758 61152
rect 50433 61149 50445 61152
rect 50479 61149 50491 61183
rect 50433 61143 50491 61149
rect 51074 61140 51080 61192
rect 51132 61180 51138 61192
rect 51353 61183 51411 61189
rect 51353 61180 51365 61183
rect 51132 61152 51365 61180
rect 51132 61140 51138 61152
rect 51353 61149 51365 61152
rect 51399 61149 51411 61183
rect 51353 61143 51411 61149
rect 51626 61140 51632 61192
rect 51684 61180 51690 61192
rect 52089 61183 52147 61189
rect 52089 61180 52101 61183
rect 51684 61152 52101 61180
rect 51684 61140 51690 61152
rect 52089 61149 52101 61152
rect 52135 61149 52147 61183
rect 53190 61180 53196 61192
rect 53151 61152 53196 61180
rect 52089 61143 52147 61149
rect 53190 61140 53196 61152
rect 53248 61140 53254 61192
rect 54110 61180 54116 61192
rect 54071 61152 54116 61180
rect 54110 61140 54116 61152
rect 54168 61140 54174 61192
rect 55490 61180 55496 61192
rect 55451 61152 55496 61180
rect 55490 61140 55496 61152
rect 55548 61140 55554 61192
rect 56042 61140 56048 61192
rect 56100 61180 56106 61192
rect 56505 61183 56563 61189
rect 56505 61180 56517 61183
rect 56100 61152 56517 61180
rect 56100 61140 56106 61152
rect 56505 61149 56517 61152
rect 56551 61149 56563 61183
rect 56505 61143 56563 61149
rect 57514 61140 57520 61192
rect 57572 61180 57578 61192
rect 58161 61183 58219 61189
rect 58161 61180 58173 61183
rect 57572 61152 58173 61180
rect 57572 61140 57578 61152
rect 58161 61149 58173 61152
rect 58207 61149 58219 61183
rect 58161 61143 58219 61149
rect 38473 61115 38531 61121
rect 38473 61112 38485 61115
rect 35820 61084 38485 61112
rect 35713 61075 35771 61081
rect 38473 61081 38485 61084
rect 38519 61081 38531 61115
rect 38473 61075 38531 61081
rect 39758 61072 39764 61124
rect 39816 61112 39822 61124
rect 42886 61112 42892 61124
rect 39816 61084 41828 61112
rect 42847 61084 42892 61112
rect 39816 61072 39822 61084
rect 20671 61016 21312 61044
rect 20671 61013 20683 61016
rect 20625 61007 20683 61013
rect 21450 61004 21456 61056
rect 21508 61044 21514 61056
rect 22465 61047 22523 61053
rect 22465 61044 22477 61047
rect 21508 61016 22477 61044
rect 21508 61004 21514 61016
rect 22465 61013 22477 61016
rect 22511 61013 22523 61047
rect 22465 61007 22523 61013
rect 23750 61004 23756 61056
rect 23808 61044 23814 61056
rect 23937 61047 23995 61053
rect 23937 61044 23949 61047
rect 23808 61016 23949 61044
rect 23808 61004 23814 61016
rect 23937 61013 23949 61016
rect 23983 61013 23995 61047
rect 27338 61044 27344 61056
rect 27299 61016 27344 61044
rect 23937 61007 23995 61013
rect 27338 61004 27344 61016
rect 27396 61004 27402 61056
rect 29914 61044 29920 61056
rect 29875 61016 29920 61044
rect 29914 61004 29920 61016
rect 29972 61004 29978 61056
rect 33502 61004 33508 61056
rect 33560 61044 33566 61056
rect 34149 61047 34207 61053
rect 34149 61044 34161 61047
rect 33560 61016 34161 61044
rect 33560 61004 33566 61016
rect 34149 61013 34161 61016
rect 34195 61013 34207 61047
rect 34149 61007 34207 61013
rect 34238 61004 34244 61056
rect 34296 61044 34302 61056
rect 35069 61047 35127 61053
rect 35069 61044 35081 61047
rect 34296 61016 35081 61044
rect 34296 61004 34302 61016
rect 35069 61013 35081 61016
rect 35115 61013 35127 61047
rect 35069 61007 35127 61013
rect 35342 61004 35348 61056
rect 35400 61044 35406 61056
rect 35805 61047 35863 61053
rect 35805 61044 35817 61047
rect 35400 61016 35817 61044
rect 35400 61004 35406 61016
rect 35805 61013 35817 61016
rect 35851 61013 35863 61047
rect 35805 61007 35863 61013
rect 36078 61004 36084 61056
rect 36136 61044 36142 61056
rect 36541 61047 36599 61053
rect 36541 61044 36553 61047
rect 36136 61016 36553 61044
rect 36136 61004 36142 61016
rect 36541 61013 36553 61016
rect 36587 61013 36599 61047
rect 36541 61007 36599 61013
rect 37274 61004 37280 61056
rect 37332 61044 37338 61056
rect 37645 61047 37703 61053
rect 37645 61044 37657 61047
rect 37332 61016 37657 61044
rect 37332 61004 37338 61016
rect 37645 61013 37657 61016
rect 37691 61013 37703 61047
rect 39114 61044 39120 61056
rect 39075 61016 39120 61044
rect 37645 61007 37703 61013
rect 39114 61004 39120 61016
rect 39172 61004 39178 61056
rect 40310 61004 40316 61056
rect 40368 61044 40374 61056
rect 40957 61047 41015 61053
rect 40957 61044 40969 61047
rect 40368 61016 40969 61044
rect 40368 61004 40374 61016
rect 40957 61013 40969 61016
rect 41003 61013 41015 61047
rect 41690 61044 41696 61056
rect 41651 61016 41696 61044
rect 40957 61007 41015 61013
rect 41690 61004 41696 61016
rect 41748 61004 41754 61056
rect 41800 61044 41828 61084
rect 42886 61072 42892 61084
rect 42944 61072 42950 61124
rect 46934 61072 46940 61124
rect 46992 61112 46998 61124
rect 49513 61115 49571 61121
rect 49513 61112 49525 61115
rect 46992 61084 49525 61112
rect 46992 61072 46998 61084
rect 49513 61081 49525 61084
rect 49559 61081 49571 61115
rect 53469 61115 53527 61121
rect 53469 61112 53481 61115
rect 49513 61075 49571 61081
rect 49988 61084 53481 61112
rect 43717 61047 43775 61053
rect 43717 61044 43729 61047
rect 41800 61016 43729 61044
rect 43717 61013 43729 61016
rect 43763 61013 43775 61047
rect 45370 61044 45376 61056
rect 45331 61016 45376 61044
rect 43717 61007 43775 61013
rect 45370 61004 45376 61016
rect 45428 61004 45434 61056
rect 46106 61044 46112 61056
rect 46067 61016 46112 61044
rect 46106 61004 46112 61016
rect 46164 61004 46170 61056
rect 46842 61044 46848 61056
rect 46803 61016 46848 61044
rect 46842 61004 46848 61016
rect 46900 61004 46906 61056
rect 47578 61004 47584 61056
rect 47636 61044 47642 61056
rect 49988 61044 50016 61084
rect 53469 61081 53481 61084
rect 53515 61081 53527 61115
rect 55769 61115 55827 61121
rect 55769 61112 55781 61115
rect 53469 61075 53527 61081
rect 53576 61084 55781 61112
rect 47636 61016 50016 61044
rect 47636 61004 47642 61016
rect 50062 61004 50068 61056
rect 50120 61044 50126 61056
rect 50525 61047 50583 61053
rect 50525 61044 50537 61047
rect 50120 61016 50537 61044
rect 50120 61004 50126 61016
rect 50525 61013 50537 61016
rect 50571 61013 50583 61047
rect 50525 61007 50583 61013
rect 51810 61004 51816 61056
rect 51868 61044 51874 61056
rect 53576 61044 53604 61084
rect 55769 61081 55781 61084
rect 55815 61081 55827 61115
rect 58342 61112 58348 61124
rect 58303 61084 58348 61112
rect 55769 61075 55827 61081
rect 58342 61072 58348 61084
rect 58400 61072 58406 61124
rect 54294 61044 54300 61056
rect 51868 61016 53604 61044
rect 54255 61016 54300 61044
rect 51868 61004 51874 61016
rect 54294 61004 54300 61016
rect 54352 61004 54358 61056
rect 1104 60954 58880 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 58880 60954
rect 1104 60880 58880 60902
rect 10318 60800 10324 60852
rect 10376 60840 10382 60852
rect 22186 60840 22192 60852
rect 10376 60812 22192 60840
rect 10376 60800 10382 60812
rect 22186 60800 22192 60812
rect 22244 60800 22250 60852
rect 27154 60800 27160 60852
rect 27212 60840 27218 60852
rect 46842 60840 46848 60852
rect 27212 60812 46848 60840
rect 27212 60800 27218 60812
rect 46842 60800 46848 60812
rect 46900 60800 46906 60852
rect 3970 60772 3976 60784
rect 3931 60744 3976 60772
rect 3970 60732 3976 60744
rect 4028 60732 4034 60784
rect 5442 60772 5448 60784
rect 5403 60744 5448 60772
rect 5442 60732 5448 60744
rect 5500 60732 5506 60784
rect 8294 60732 8300 60784
rect 8352 60772 8358 60784
rect 8389 60775 8447 60781
rect 8389 60772 8401 60775
rect 8352 60744 8401 60772
rect 8352 60732 8358 60744
rect 8389 60741 8401 60744
rect 8435 60741 8447 60775
rect 9858 60772 9864 60784
rect 9819 60744 9864 60772
rect 8389 60735 8447 60741
rect 9858 60732 9864 60744
rect 9916 60732 9922 60784
rect 13538 60772 13544 60784
rect 13499 60744 13544 60772
rect 13538 60732 13544 60744
rect 13596 60732 13602 60784
rect 14274 60772 14280 60784
rect 14235 60744 14280 60772
rect 14274 60732 14280 60744
rect 14332 60732 14338 60784
rect 15746 60772 15752 60784
rect 15707 60744 15752 60772
rect 15746 60732 15752 60744
rect 15804 60732 15810 60784
rect 19334 60732 19340 60784
rect 19392 60772 19398 60784
rect 19429 60775 19487 60781
rect 19429 60772 19441 60775
rect 19392 60744 19441 60772
rect 19392 60732 19398 60744
rect 19429 60741 19441 60744
rect 19475 60741 19487 60775
rect 23290 60772 23296 60784
rect 23251 60744 23296 60772
rect 19429 60735 19487 60741
rect 23290 60732 23296 60744
rect 23348 60732 23354 60784
rect 24578 60772 24584 60784
rect 24539 60744 24584 60772
rect 24578 60732 24584 60744
rect 24636 60732 24642 60784
rect 27522 60772 27528 60784
rect 27483 60744 27528 60772
rect 27522 60732 27528 60744
rect 27580 60732 27586 60784
rect 28994 60772 29000 60784
rect 28955 60744 29000 60772
rect 28994 60732 29000 60744
rect 29052 60732 29058 60784
rect 30374 60732 30380 60784
rect 30432 60772 30438 60784
rect 30469 60775 30527 60781
rect 30469 60772 30481 60775
rect 30432 60744 30481 60772
rect 30432 60732 30438 60744
rect 30469 60741 30481 60744
rect 30515 60741 30527 60775
rect 36354 60772 36360 60784
rect 36315 60744 36360 60772
rect 30469 60735 30527 60741
rect 36354 60732 36360 60744
rect 36412 60732 36418 60784
rect 41414 60732 41420 60784
rect 41472 60772 41478 60784
rect 41509 60775 41567 60781
rect 41509 60772 41521 60775
rect 41472 60744 41521 60772
rect 41472 60732 41478 60744
rect 41509 60741 41521 60744
rect 41555 60741 41567 60775
rect 46658 60772 46664 60784
rect 46619 60744 46664 60772
rect 41509 60735 41567 60741
rect 46658 60732 46664 60744
rect 46716 60732 46722 60784
rect 50154 60732 50160 60784
rect 50212 60772 50218 60784
rect 50341 60775 50399 60781
rect 50341 60772 50353 60775
rect 50212 60744 50353 60772
rect 50212 60732 50218 60744
rect 50341 60741 50353 60744
rect 50387 60741 50399 60775
rect 50341 60735 50399 60741
rect 52454 60732 52460 60784
rect 52512 60772 52518 60784
rect 53009 60775 53067 60781
rect 53009 60772 53021 60775
rect 52512 60744 53021 60772
rect 52512 60732 52518 60744
rect 53009 60741 53021 60744
rect 53055 60741 53067 60775
rect 53009 60735 53067 60741
rect 1578 60704 1584 60716
rect 1539 60676 1584 60704
rect 1578 60664 1584 60676
rect 1636 60664 1642 60716
rect 3142 60704 3148 60716
rect 3103 60676 3148 60704
rect 3142 60664 3148 60676
rect 3200 60664 3206 60716
rect 14461 60707 14519 60713
rect 14461 60673 14473 60707
rect 14507 60704 14519 60707
rect 21266 60704 21272 60716
rect 14507 60676 21272 60704
rect 14507 60673 14519 60676
rect 14461 60667 14519 60673
rect 21266 60664 21272 60676
rect 21324 60664 21330 60716
rect 22094 60664 22100 60716
rect 22152 60704 22158 60716
rect 22152 60676 22197 60704
rect 22152 60664 22158 60676
rect 24670 60664 24676 60716
rect 24728 60704 24734 60716
rect 35066 60704 35072 60716
rect 24728 60676 35072 60704
rect 24728 60664 24734 60676
rect 35066 60664 35072 60676
rect 35124 60664 35130 60716
rect 41598 60704 41604 60716
rect 36556 60676 41604 60704
rect 1857 60639 1915 60645
rect 1857 60605 1869 60639
rect 1903 60636 1915 60639
rect 4798 60636 4804 60648
rect 1903 60608 4804 60636
rect 1903 60605 1915 60608
rect 1857 60599 1915 60605
rect 4798 60596 4804 60608
rect 4856 60596 4862 60648
rect 8573 60639 8631 60645
rect 8573 60605 8585 60639
rect 8619 60636 8631 60639
rect 13630 60636 13636 60648
rect 8619 60608 13636 60636
rect 8619 60605 8631 60608
rect 8573 60599 8631 60605
rect 13630 60596 13636 60608
rect 13688 60596 13694 60648
rect 13725 60639 13783 60645
rect 13725 60605 13737 60639
rect 13771 60636 13783 60639
rect 22462 60636 22468 60648
rect 13771 60608 22468 60636
rect 13771 60605 13783 60608
rect 13725 60599 13783 60605
rect 22462 60596 22468 60608
rect 22520 60596 22526 60648
rect 22646 60636 22652 60648
rect 22559 60608 22652 60636
rect 22646 60596 22652 60608
rect 22704 60636 22710 60648
rect 36556 60636 36584 60676
rect 41598 60664 41604 60676
rect 41656 60664 41662 60716
rect 54662 60704 54668 60716
rect 54623 60676 54668 60704
rect 54662 60664 54668 60676
rect 54720 60664 54726 60716
rect 55398 60704 55404 60716
rect 55359 60676 55404 60704
rect 55398 60664 55404 60676
rect 55456 60664 55462 60716
rect 56134 60704 56140 60716
rect 56095 60676 56140 60704
rect 56134 60664 56140 60676
rect 56192 60664 56198 60716
rect 56870 60704 56876 60716
rect 56831 60676 56876 60704
rect 56870 60664 56876 60676
rect 56928 60664 56934 60716
rect 58066 60704 58072 60716
rect 58027 60676 58072 60704
rect 58066 60664 58072 60676
rect 58124 60664 58130 60716
rect 22704 60608 36584 60636
rect 22704 60596 22710 60608
rect 36630 60596 36636 60648
rect 36688 60636 36694 60648
rect 46934 60636 46940 60648
rect 36688 60608 46940 60636
rect 36688 60596 36694 60608
rect 46934 60596 46940 60608
rect 46992 60596 46998 60648
rect 4157 60571 4215 60577
rect 4157 60537 4169 60571
rect 4203 60568 4215 60571
rect 4614 60568 4620 60580
rect 4203 60540 4620 60568
rect 4203 60537 4215 60540
rect 4157 60531 4215 60537
rect 4614 60528 4620 60540
rect 4672 60528 4678 60580
rect 5629 60571 5687 60577
rect 5629 60537 5641 60571
rect 5675 60568 5687 60571
rect 19613 60571 19671 60577
rect 5675 60540 17264 60568
rect 5675 60537 5687 60540
rect 5629 60531 5687 60537
rect 3326 60500 3332 60512
rect 3287 60472 3332 60500
rect 3326 60460 3332 60472
rect 3384 60460 3390 60512
rect 9950 60500 9956 60512
rect 9911 60472 9956 60500
rect 9950 60460 9956 60472
rect 10008 60460 10014 60512
rect 15838 60500 15844 60512
rect 15799 60472 15844 60500
rect 15838 60460 15844 60472
rect 15896 60460 15902 60512
rect 17236 60500 17264 60540
rect 19613 60537 19625 60571
rect 19659 60568 19671 60571
rect 20346 60568 20352 60580
rect 19659 60540 20352 60568
rect 19659 60537 19671 60540
rect 19613 60531 19671 60537
rect 20346 60528 20352 60540
rect 20404 60528 20410 60580
rect 23477 60571 23535 60577
rect 23477 60537 23489 60571
rect 23523 60568 23535 60571
rect 24486 60568 24492 60580
rect 23523 60540 24492 60568
rect 23523 60537 23535 60540
rect 23477 60531 23535 60537
rect 24486 60528 24492 60540
rect 24544 60528 24550 60580
rect 25222 60528 25228 60580
rect 25280 60568 25286 60580
rect 58253 60571 58311 60577
rect 58253 60568 58265 60571
rect 25280 60540 58265 60568
rect 25280 60528 25286 60540
rect 58253 60537 58265 60540
rect 58299 60537 58311 60571
rect 58253 60531 58311 60537
rect 22830 60500 22836 60512
rect 17236 60472 22836 60500
rect 22830 60460 22836 60472
rect 22888 60460 22894 60512
rect 24394 60460 24400 60512
rect 24452 60500 24458 60512
rect 24673 60503 24731 60509
rect 24673 60500 24685 60503
rect 24452 60472 24685 60500
rect 24452 60460 24458 60472
rect 24673 60469 24685 60472
rect 24719 60469 24731 60503
rect 24673 60463 24731 60469
rect 27617 60503 27675 60509
rect 27617 60469 27629 60503
rect 27663 60500 27675 60503
rect 28074 60500 28080 60512
rect 27663 60472 28080 60500
rect 27663 60469 27675 60472
rect 27617 60463 27675 60469
rect 28074 60460 28080 60472
rect 28132 60460 28138 60512
rect 28166 60460 28172 60512
rect 28224 60500 28230 60512
rect 28350 60500 28356 60512
rect 28224 60472 28356 60500
rect 28224 60460 28230 60472
rect 28350 60460 28356 60472
rect 28408 60460 28414 60512
rect 29086 60500 29092 60512
rect 29047 60472 29092 60500
rect 29086 60460 29092 60472
rect 29144 60460 29150 60512
rect 30561 60503 30619 60509
rect 30561 60469 30573 60503
rect 30607 60500 30619 60503
rect 35618 60500 35624 60512
rect 30607 60472 35624 60500
rect 30607 60469 30619 60472
rect 30561 60463 30619 60469
rect 35618 60460 35624 60472
rect 35676 60460 35682 60512
rect 35710 60460 35716 60512
rect 35768 60500 35774 60512
rect 36449 60503 36507 60509
rect 36449 60500 36461 60503
rect 35768 60472 36461 60500
rect 35768 60460 35774 60472
rect 36449 60469 36461 60472
rect 36495 60469 36507 60503
rect 36449 60463 36507 60469
rect 41601 60503 41659 60509
rect 41601 60469 41613 60503
rect 41647 60500 41659 60503
rect 41966 60500 41972 60512
rect 41647 60472 41972 60500
rect 41647 60469 41659 60472
rect 41601 60463 41659 60469
rect 41966 60460 41972 60472
rect 42024 60460 42030 60512
rect 44174 60460 44180 60512
rect 44232 60500 44238 60512
rect 46753 60503 46811 60509
rect 46753 60500 46765 60503
rect 44232 60472 46765 60500
rect 44232 60460 44238 60472
rect 46753 60469 46765 60472
rect 46799 60469 46811 60503
rect 50430 60500 50436 60512
rect 50391 60472 50436 60500
rect 46753 60463 46811 60469
rect 50430 60460 50436 60472
rect 50488 60460 50494 60512
rect 53098 60500 53104 60512
rect 53059 60472 53104 60500
rect 53098 60460 53104 60472
rect 53156 60460 53162 60512
rect 54846 60500 54852 60512
rect 54807 60472 54852 60500
rect 54846 60460 54852 60472
rect 54904 60460 54910 60512
rect 55582 60500 55588 60512
rect 55543 60472 55588 60500
rect 55582 60460 55588 60472
rect 55640 60460 55646 60512
rect 56318 60500 56324 60512
rect 56279 60472 56324 60500
rect 56318 60460 56324 60472
rect 56376 60460 56382 60512
rect 57054 60500 57060 60512
rect 57015 60472 57060 60500
rect 57054 60460 57060 60472
rect 57112 60460 57118 60512
rect 1104 60410 58880 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 58880 60410
rect 1104 60336 58880 60358
rect 9950 60256 9956 60308
rect 10008 60296 10014 60308
rect 19242 60296 19248 60308
rect 10008 60268 19248 60296
rect 10008 60256 10014 60268
rect 19242 60256 19248 60268
rect 19300 60256 19306 60308
rect 20272 60268 22876 60296
rect 6549 60231 6607 60237
rect 6549 60197 6561 60231
rect 6595 60228 6607 60231
rect 6638 60228 6644 60240
rect 6595 60200 6644 60228
rect 6595 60197 6607 60200
rect 6549 60191 6607 60197
rect 6638 60188 6644 60200
rect 6696 60188 6702 60240
rect 13630 60188 13636 60240
rect 13688 60228 13694 60240
rect 13688 60200 18644 60228
rect 13688 60188 13694 60200
rect 15838 60120 15844 60172
rect 15896 60160 15902 60172
rect 18049 60163 18107 60169
rect 18049 60160 18061 60163
rect 15896 60132 18061 60160
rect 15896 60120 15902 60132
rect 18049 60129 18061 60132
rect 18095 60129 18107 60163
rect 18049 60123 18107 60129
rect 2590 60092 2596 60104
rect 2551 60064 2596 60092
rect 2590 60052 2596 60064
rect 2648 60052 2654 60104
rect 5994 60092 6000 60104
rect 5955 60064 6000 60092
rect 5994 60052 6000 60064
rect 6052 60052 6058 60104
rect 6270 60092 6276 60104
rect 6231 60064 6276 60092
rect 6270 60052 6276 60064
rect 6328 60052 6334 60104
rect 6417 60095 6475 60101
rect 6417 60061 6429 60095
rect 6463 60092 6475 60095
rect 7006 60092 7012 60104
rect 6463 60064 7012 60092
rect 6463 60061 6475 60064
rect 6417 60055 6475 60061
rect 7006 60052 7012 60064
rect 7064 60052 7070 60104
rect 18616 60101 18644 60200
rect 18233 60095 18291 60101
rect 18233 60061 18245 60095
rect 18279 60061 18291 60095
rect 18233 60055 18291 60061
rect 18601 60095 18659 60101
rect 18601 60061 18613 60095
rect 18647 60061 18659 60095
rect 18601 60055 18659 60061
rect 18785 60095 18843 60101
rect 18785 60061 18797 60095
rect 18831 60092 18843 60095
rect 19426 60092 19432 60104
rect 18831 60064 19432 60092
rect 18831 60061 18843 60064
rect 18785 60055 18843 60061
rect 1670 60024 1676 60036
rect 1631 59996 1676 60024
rect 1670 59984 1676 59996
rect 1728 59984 1734 60036
rect 2038 60024 2044 60036
rect 1999 59996 2044 60024
rect 2038 59984 2044 59996
rect 2096 59984 2102 60036
rect 3878 59984 3884 60036
rect 3936 60024 3942 60036
rect 6181 60027 6239 60033
rect 6181 60024 6193 60027
rect 3936 59996 6193 60024
rect 3936 59984 3942 59996
rect 6181 59993 6193 59996
rect 6227 60024 6239 60027
rect 6730 60024 6736 60036
rect 6227 59996 6736 60024
rect 6227 59993 6239 59996
rect 6181 59987 6239 59993
rect 6730 59984 6736 59996
rect 6788 59984 6794 60036
rect 18248 60024 18276 60055
rect 19426 60052 19432 60064
rect 19484 60052 19490 60104
rect 19978 60092 19984 60104
rect 19939 60064 19984 60092
rect 19978 60052 19984 60064
rect 20036 60052 20042 60104
rect 20272 60101 20300 60268
rect 20530 60228 20536 60240
rect 20491 60200 20536 60228
rect 20530 60188 20536 60200
rect 20588 60188 20594 60240
rect 22646 60228 22652 60240
rect 21100 60200 22652 60228
rect 20257 60095 20315 60101
rect 20257 60061 20269 60095
rect 20303 60061 20315 60095
rect 20257 60055 20315 60061
rect 20401 60095 20459 60101
rect 20401 60061 20413 60095
rect 20447 60092 20459 60095
rect 21100 60092 21128 60200
rect 22646 60188 22652 60200
rect 22704 60188 22710 60240
rect 22848 60228 22876 60268
rect 22922 60256 22928 60308
rect 22980 60296 22986 60308
rect 25958 60296 25964 60308
rect 22980 60268 25964 60296
rect 22980 60256 22986 60268
rect 25958 60256 25964 60268
rect 26016 60256 26022 60308
rect 26786 60256 26792 60308
rect 26844 60296 26850 60308
rect 29730 60296 29736 60308
rect 26844 60268 29736 60296
rect 26844 60256 26850 60268
rect 29730 60256 29736 60268
rect 29788 60256 29794 60308
rect 30006 60256 30012 60308
rect 30064 60296 30070 60308
rect 58250 60296 58256 60308
rect 30064 60268 58256 60296
rect 30064 60256 30070 60268
rect 58250 60256 58256 60268
rect 58308 60256 58314 60308
rect 25866 60228 25872 60240
rect 22848 60200 25872 60228
rect 25866 60188 25872 60200
rect 25924 60188 25930 60240
rect 26050 60188 26056 60240
rect 26108 60228 26114 60240
rect 27433 60231 27491 60237
rect 27433 60228 27445 60231
rect 26108 60200 27445 60228
rect 26108 60188 26114 60200
rect 27433 60197 27445 60200
rect 27479 60197 27491 60231
rect 28718 60228 28724 60240
rect 27433 60191 27491 60197
rect 27724 60200 28724 60228
rect 21266 60120 21272 60172
rect 21324 60160 21330 60172
rect 26970 60160 26976 60172
rect 21324 60132 26976 60160
rect 21324 60120 21330 60132
rect 26970 60120 26976 60132
rect 27028 60120 27034 60172
rect 20447 60064 21128 60092
rect 20447 60061 20459 60064
rect 20401 60055 20459 60061
rect 21174 60052 21180 60104
rect 21232 60092 21238 60104
rect 22278 60092 22284 60104
rect 21232 60064 21277 60092
rect 22239 60064 22284 60092
rect 21232 60052 21238 60064
rect 22278 60052 22284 60064
rect 22336 60052 22342 60104
rect 22646 60052 22652 60104
rect 22704 60101 22710 60104
rect 22704 60092 22712 60101
rect 22704 60064 22749 60092
rect 22704 60055 22712 60064
rect 22704 60052 22710 60055
rect 23014 60052 23020 60104
rect 23072 60092 23078 60104
rect 23842 60101 23848 60104
rect 23385 60095 23443 60101
rect 23385 60092 23397 60095
rect 23072 60064 23397 60092
rect 23072 60052 23078 60064
rect 23385 60061 23397 60064
rect 23431 60061 23443 60095
rect 23385 60055 23443 60061
rect 23805 60095 23848 60101
rect 23805 60061 23817 60095
rect 23805 60055 23848 60061
rect 23842 60052 23848 60055
rect 23900 60052 23906 60104
rect 23934 60052 23940 60104
rect 23992 60101 23998 60104
rect 23992 60095 24012 60101
rect 24000 60061 24012 60095
rect 23992 60055 24012 60061
rect 24673 60095 24731 60101
rect 24673 60061 24685 60095
rect 24719 60090 24731 60095
rect 24762 60090 24768 60104
rect 24719 60062 24768 60090
rect 24719 60061 24731 60062
rect 24673 60055 24731 60061
rect 23992 60052 23998 60055
rect 24762 60052 24768 60062
rect 24820 60052 24826 60104
rect 25130 60092 25136 60104
rect 25091 60064 25136 60092
rect 25130 60052 25136 60064
rect 25188 60052 25194 60104
rect 25222 60052 25228 60104
rect 25280 60092 25286 60104
rect 25498 60092 25504 60104
rect 25280 60064 25325 60092
rect 25459 60064 25504 60092
rect 25280 60052 25286 60064
rect 25498 60052 25504 60064
rect 25556 60052 25562 60104
rect 25777 60095 25835 60101
rect 25777 60092 25789 60095
rect 25608 60064 25789 60092
rect 20165 60027 20223 60033
rect 20165 60024 20177 60027
rect 18248 59996 20177 60024
rect 20165 59993 20177 59996
rect 20211 60024 20223 60027
rect 21545 60027 21603 60033
rect 21545 60024 21557 60027
rect 20211 59996 21557 60024
rect 20211 59993 20223 59996
rect 20165 59987 20223 59993
rect 21545 59993 21557 59996
rect 21591 60024 21603 60027
rect 22465 60027 22523 60033
rect 22465 60024 22477 60027
rect 21591 59996 22477 60024
rect 21591 59993 21603 59996
rect 21545 59987 21603 59993
rect 22465 59993 22477 59996
rect 22511 59993 22523 60027
rect 22465 59987 22523 59993
rect 2498 59916 2504 59968
rect 2556 59956 2562 59968
rect 2685 59959 2743 59965
rect 2685 59956 2697 59959
rect 2556 59928 2697 59956
rect 2556 59916 2562 59928
rect 2685 59925 2697 59928
rect 2731 59925 2743 59959
rect 17678 59956 17684 59968
rect 17639 59928 17684 59956
rect 2685 59919 2743 59925
rect 17678 59916 17684 59928
rect 17736 59916 17742 59968
rect 22480 59956 22508 59987
rect 22554 59984 22560 60036
rect 22612 60024 22618 60036
rect 22612 59996 22657 60024
rect 22612 59984 22618 59996
rect 22738 59984 22744 60036
rect 22796 60024 22802 60036
rect 22850 60027 22908 60033
rect 22850 60024 22862 60027
rect 22796 59996 22862 60024
rect 22796 59984 22802 59996
rect 22850 59993 22862 59996
rect 22896 59993 22908 60027
rect 23566 60024 23572 60036
rect 23527 59996 23572 60024
rect 22850 59987 22908 59993
rect 23566 59984 23572 59996
rect 23624 59984 23630 60036
rect 23661 60027 23719 60033
rect 23661 59993 23673 60027
rect 23707 60024 23719 60027
rect 24946 60024 24952 60036
rect 23707 59996 24952 60024
rect 23707 59993 23719 59996
rect 23661 59987 23719 59993
rect 24946 59984 24952 59996
rect 25004 59984 25010 60036
rect 25608 60024 25636 60064
rect 25777 60061 25789 60064
rect 25823 60061 25835 60095
rect 25958 60092 25964 60104
rect 25919 60064 25964 60092
rect 25777 60055 25835 60061
rect 25958 60052 25964 60064
rect 26016 60052 26022 60104
rect 26418 60052 26424 60104
rect 26476 60092 26482 60104
rect 26789 60095 26847 60101
rect 26789 60092 26801 60095
rect 26476 60064 26801 60092
rect 26476 60052 26482 60064
rect 26789 60061 26801 60064
rect 26835 60061 26847 60095
rect 26789 60055 26847 60061
rect 26878 60052 26884 60104
rect 26936 60092 26942 60104
rect 27154 60092 27160 60104
rect 26936 60064 26981 60092
rect 27115 60064 27160 60092
rect 26936 60052 26942 60064
rect 27154 60052 27160 60064
rect 27212 60052 27218 60104
rect 27246 60052 27252 60104
rect 27304 60101 27310 60104
rect 27304 60092 27312 60101
rect 27724 60092 27752 60200
rect 28166 60120 28172 60172
rect 28224 60160 28230 60172
rect 28224 60132 28304 60160
rect 28224 60120 28230 60132
rect 27982 60092 27988 60104
rect 27304 60064 27752 60092
rect 27943 60064 27988 60092
rect 27304 60055 27312 60064
rect 27304 60052 27310 60055
rect 27982 60052 27988 60064
rect 28040 60052 28046 60104
rect 28074 60052 28080 60104
rect 28132 60092 28138 60104
rect 28276 60092 28304 60132
rect 28465 60101 28493 60200
rect 28718 60188 28724 60200
rect 28776 60188 28782 60240
rect 28810 60188 28816 60240
rect 28868 60228 28874 60240
rect 56226 60228 56232 60240
rect 28868 60200 33824 60228
rect 28868 60188 28874 60200
rect 28534 60120 28540 60172
rect 28592 60160 28598 60172
rect 29638 60160 29644 60172
rect 28592 60132 29644 60160
rect 28592 60120 28598 60132
rect 29638 60120 29644 60132
rect 29696 60120 29702 60172
rect 30098 60120 30104 60172
rect 30156 60160 30162 60172
rect 33597 60163 33655 60169
rect 33597 60160 33609 60163
rect 30156 60132 33609 60160
rect 30156 60120 30162 60132
rect 33597 60129 33609 60132
rect 33643 60129 33655 60163
rect 33597 60123 33655 60129
rect 33796 60104 33824 60200
rect 41708 60200 56232 60228
rect 37182 60160 37188 60172
rect 34348 60132 37188 60160
rect 28361 60095 28419 60101
rect 28361 60092 28373 60095
rect 28132 60064 28177 60092
rect 28276 60064 28373 60092
rect 28132 60052 28138 60064
rect 28361 60061 28373 60064
rect 28407 60061 28419 60095
rect 28361 60055 28419 60061
rect 28450 60095 28508 60101
rect 28450 60061 28462 60095
rect 28496 60061 28508 60095
rect 28450 60055 28508 60061
rect 28718 60052 28724 60104
rect 28776 60092 28782 60104
rect 28994 60092 29000 60104
rect 28776 60064 29000 60092
rect 28776 60052 28782 60064
rect 28994 60052 29000 60064
rect 29052 60052 29058 60104
rect 29178 60092 29184 60104
rect 29139 60064 29184 60092
rect 29178 60052 29184 60064
rect 29236 60092 29242 60104
rect 29733 60095 29791 60101
rect 29733 60092 29745 60095
rect 29236 60064 29745 60092
rect 29236 60052 29242 60064
rect 29733 60061 29745 60064
rect 29779 60061 29791 60095
rect 29733 60055 29791 60061
rect 29826 60095 29884 60101
rect 29826 60061 29838 60095
rect 29872 60061 29884 60095
rect 29826 60055 29884 60061
rect 27065 60027 27123 60033
rect 27065 60024 27077 60027
rect 25608 59996 27077 60024
rect 25608 59956 25636 59996
rect 27065 59993 27077 59996
rect 27111 60024 27123 60027
rect 28261 60027 28319 60033
rect 28261 60024 28273 60027
rect 27111 59996 28273 60024
rect 27111 59993 27123 59996
rect 27065 59987 27123 59993
rect 28261 59993 28273 59996
rect 28307 60024 28319 60027
rect 28810 60024 28816 60036
rect 28307 59996 28816 60024
rect 28307 59993 28319 59996
rect 28261 59987 28319 59993
rect 28810 59984 28816 59996
rect 28868 59984 28874 60036
rect 29086 59984 29092 60036
rect 29144 60024 29150 60036
rect 29841 60024 29869 60055
rect 30190 60052 30196 60104
rect 30248 60101 30254 60104
rect 30248 60092 30256 60101
rect 33778 60092 33784 60104
rect 30248 60064 30293 60092
rect 33691 60064 33784 60092
rect 30248 60055 30256 60064
rect 30248 60052 30254 60055
rect 33778 60052 33784 60064
rect 33836 60052 33842 60104
rect 34146 60092 34152 60104
rect 34107 60064 34152 60092
rect 34146 60052 34152 60064
rect 34204 60052 34210 60104
rect 34348 60101 34376 60132
rect 37182 60120 37188 60132
rect 37240 60120 37246 60172
rect 41708 60169 41736 60200
rect 56226 60188 56232 60200
rect 56284 60188 56290 60240
rect 41693 60163 41751 60169
rect 41693 60129 41705 60163
rect 41739 60129 41751 60163
rect 41693 60123 41751 60129
rect 41874 60120 41880 60172
rect 41932 60160 41938 60172
rect 43533 60163 43591 60169
rect 43533 60160 43545 60163
rect 41932 60132 43545 60160
rect 41932 60120 41938 60132
rect 43533 60129 43545 60132
rect 43579 60129 43591 60163
rect 43533 60123 43591 60129
rect 53742 60120 53748 60172
rect 53800 60160 53806 60172
rect 57425 60163 57483 60169
rect 57425 60160 57437 60163
rect 53800 60132 57437 60160
rect 53800 60120 53806 60132
rect 57425 60129 57437 60132
rect 57471 60129 57483 60163
rect 57425 60123 57483 60129
rect 34333 60095 34391 60101
rect 34333 60061 34345 60095
rect 34379 60061 34391 60095
rect 36630 60092 36636 60104
rect 34333 60055 34391 60061
rect 35544 60064 36636 60092
rect 30006 60024 30012 60036
rect 29144 59996 29869 60024
rect 29967 59996 30012 60024
rect 29144 59984 29150 59996
rect 30006 59984 30012 59996
rect 30064 59984 30070 60036
rect 30101 60027 30159 60033
rect 30101 59993 30113 60027
rect 30147 60024 30159 60027
rect 35544 60024 35572 60064
rect 36630 60052 36636 60064
rect 36688 60052 36694 60104
rect 41598 60092 41604 60104
rect 41559 60064 41604 60092
rect 41598 60052 41604 60064
rect 41656 60092 41662 60104
rect 41782 60092 41788 60104
rect 41656 60064 41788 60092
rect 41656 60052 41662 60064
rect 41782 60052 41788 60064
rect 41840 60052 41846 60104
rect 41966 60092 41972 60104
rect 41927 60064 41972 60092
rect 41966 60052 41972 60064
rect 42024 60052 42030 60104
rect 43073 60095 43131 60101
rect 43073 60092 43085 60095
rect 42168 60064 43085 60092
rect 30147 59996 35572 60024
rect 30147 59993 30159 59996
rect 30101 59987 30159 59993
rect 35618 59984 35624 60036
rect 35676 60024 35682 60036
rect 42168 60024 42196 60064
rect 43073 60061 43085 60064
rect 43119 60061 43131 60095
rect 43254 60092 43260 60104
rect 43215 60064 43260 60092
rect 43073 60055 43131 60061
rect 43254 60052 43260 60064
rect 43312 60052 43318 60104
rect 43625 60095 43683 60101
rect 43625 60061 43637 60095
rect 43671 60061 43683 60095
rect 56502 60092 56508 60104
rect 56463 60064 56508 60092
rect 43625 60055 43683 60061
rect 42610 60024 42616 60036
rect 35676 59996 42196 60024
rect 42571 59996 42616 60024
rect 35676 59984 35682 59996
rect 42610 59984 42616 59996
rect 42668 59984 42674 60036
rect 43640 60024 43668 60055
rect 56502 60052 56508 60064
rect 56560 60052 56566 60104
rect 57238 60092 57244 60104
rect 57199 60064 57244 60092
rect 57238 60052 57244 60064
rect 57296 60052 57302 60104
rect 57974 60092 57980 60104
rect 57935 60064 57980 60092
rect 57974 60052 57980 60064
rect 58032 60052 58038 60104
rect 50430 60024 50436 60036
rect 43640 59996 50436 60024
rect 50430 59984 50436 59996
rect 50488 59984 50494 60036
rect 58345 60027 58403 60033
rect 58345 59993 58357 60027
rect 58391 60024 58403 60027
rect 58434 60024 58440 60036
rect 58391 59996 58440 60024
rect 58391 59993 58403 59996
rect 58345 59987 58403 59993
rect 58434 59984 58440 59996
rect 58492 59984 58498 60036
rect 22480 59928 25636 59956
rect 25866 59916 25872 59968
rect 25924 59956 25930 59968
rect 26234 59956 26240 59968
rect 25924 59928 26240 59956
rect 25924 59916 25930 59928
rect 26234 59916 26240 59928
rect 26292 59916 26298 59968
rect 26418 59956 26424 59968
rect 26379 59928 26424 59956
rect 26418 59916 26424 59928
rect 26476 59916 26482 59968
rect 27522 59916 27528 59968
rect 27580 59956 27586 59968
rect 28629 59959 28687 59965
rect 28629 59956 28641 59959
rect 27580 59928 28641 59956
rect 27580 59916 27586 59928
rect 28629 59925 28641 59928
rect 28675 59925 28687 59959
rect 28629 59919 28687 59925
rect 29270 59916 29276 59968
rect 29328 59956 29334 59968
rect 30377 59959 30435 59965
rect 30377 59956 30389 59959
rect 29328 59928 30389 59956
rect 29328 59916 29334 59928
rect 30377 59925 30389 59928
rect 30423 59925 30435 59959
rect 30650 59956 30656 59968
rect 30611 59928 30656 59956
rect 30377 59919 30435 59925
rect 30650 59916 30656 59928
rect 30708 59916 30714 59968
rect 32861 59959 32919 59965
rect 32861 59925 32873 59959
rect 32907 59956 32919 59959
rect 33226 59956 33232 59968
rect 32907 59928 33232 59956
rect 32907 59925 32919 59928
rect 32861 59919 32919 59925
rect 33226 59916 33232 59928
rect 33284 59956 33290 59968
rect 34885 59959 34943 59965
rect 34885 59956 34897 59959
rect 33284 59928 34897 59956
rect 33284 59916 33290 59928
rect 34885 59925 34897 59928
rect 34931 59925 34943 59959
rect 41046 59956 41052 59968
rect 41007 59928 41052 59956
rect 34885 59919 34943 59925
rect 41046 59916 41052 59928
rect 41104 59916 41110 59968
rect 56594 59956 56600 59968
rect 56555 59928 56600 59956
rect 56594 59916 56600 59928
rect 56652 59916 56658 59968
rect 1104 59866 58880 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 58880 59866
rect 1104 59792 58880 59814
rect 23566 59752 23572 59764
rect 6886 59724 23572 59752
rect 1762 59644 1768 59696
rect 1820 59684 1826 59696
rect 2409 59687 2467 59693
rect 2409 59684 2421 59687
rect 1820 59656 2421 59684
rect 1820 59644 1826 59656
rect 2409 59653 2421 59656
rect 2455 59653 2467 59687
rect 6730 59684 6736 59696
rect 6691 59656 6736 59684
rect 2409 59647 2467 59653
rect 6730 59644 6736 59656
rect 6788 59684 6794 59696
rect 6886 59684 6914 59724
rect 23566 59712 23572 59724
rect 23624 59712 23630 59764
rect 24857 59755 24915 59761
rect 24857 59721 24869 59755
rect 24903 59752 24915 59755
rect 25498 59752 25504 59764
rect 24903 59724 25504 59752
rect 24903 59721 24915 59724
rect 24857 59715 24915 59721
rect 25498 59712 25504 59724
rect 25556 59712 25562 59764
rect 26786 59752 26792 59764
rect 25700 59724 26792 59752
rect 6788 59656 6914 59684
rect 6788 59644 6794 59656
rect 15286 59644 15292 59696
rect 15344 59684 15350 59696
rect 19061 59687 19119 59693
rect 19061 59684 19073 59687
rect 15344 59656 19073 59684
rect 15344 59644 15350 59656
rect 19061 59653 19073 59656
rect 19107 59653 19119 59687
rect 19061 59647 19119 59653
rect 19242 59644 19248 59696
rect 19300 59684 19306 59696
rect 22646 59684 22652 59696
rect 19300 59656 22652 59684
rect 19300 59644 19306 59656
rect 22646 59644 22652 59656
rect 22704 59644 22710 59696
rect 24578 59684 24584 59696
rect 24539 59656 24584 59684
rect 24578 59644 24584 59656
rect 24636 59644 24642 59696
rect 1578 59616 1584 59628
rect 1539 59588 1584 59616
rect 1578 59576 1584 59588
rect 1636 59576 1642 59628
rect 5534 59576 5540 59628
rect 5592 59616 5598 59628
rect 6549 59619 6607 59625
rect 6549 59616 6561 59619
rect 5592 59588 6561 59616
rect 5592 59576 5598 59588
rect 6549 59585 6561 59588
rect 6595 59585 6607 59619
rect 6822 59616 6828 59628
rect 6783 59588 6828 59616
rect 6549 59579 6607 59585
rect 6822 59576 6828 59588
rect 6880 59576 6886 59628
rect 6917 59619 6975 59625
rect 6917 59585 6929 59619
rect 6963 59616 6975 59619
rect 7006 59616 7012 59628
rect 6963 59588 7012 59616
rect 6963 59585 6975 59588
rect 6917 59579 6975 59585
rect 7006 59576 7012 59588
rect 7064 59576 7070 59628
rect 18782 59616 18788 59628
rect 18743 59588 18788 59616
rect 18782 59576 18788 59588
rect 18840 59576 18846 59628
rect 18969 59619 19027 59625
rect 18969 59585 18981 59619
rect 19015 59585 19027 59619
rect 18969 59579 19027 59585
rect 18984 59480 19012 59579
rect 19150 59576 19156 59628
rect 19208 59625 19214 59628
rect 19208 59616 19216 59625
rect 19208 59588 19253 59616
rect 19208 59579 19216 59588
rect 19208 59576 19214 59579
rect 22186 59576 22192 59628
rect 22244 59616 22250 59628
rect 24305 59619 24363 59625
rect 24305 59616 24317 59619
rect 22244 59588 24317 59616
rect 22244 59576 22250 59588
rect 24305 59585 24317 59588
rect 24351 59585 24363 59619
rect 24489 59619 24547 59625
rect 24489 59616 24501 59619
rect 24305 59579 24363 59585
rect 24412 59588 24501 59616
rect 19426 59508 19432 59560
rect 19484 59548 19490 59560
rect 24412 59548 24440 59588
rect 24489 59585 24501 59588
rect 24535 59585 24547 59619
rect 24489 59579 24547 59585
rect 24673 59619 24731 59625
rect 24673 59585 24685 59619
rect 24719 59616 24731 59619
rect 24762 59616 24768 59628
rect 24719 59588 24768 59616
rect 24719 59585 24731 59588
rect 24673 59579 24731 59585
rect 24762 59576 24768 59588
rect 24820 59576 24826 59628
rect 25593 59619 25651 59625
rect 25593 59585 25605 59619
rect 25639 59616 25651 59619
rect 25700 59616 25728 59724
rect 26786 59712 26792 59724
rect 26844 59712 26850 59764
rect 29178 59712 29184 59764
rect 29236 59752 29242 59764
rect 30650 59752 30656 59764
rect 29236 59724 30656 59752
rect 29236 59712 29242 59724
rect 30650 59712 30656 59724
rect 30708 59712 30714 59764
rect 33778 59712 33784 59764
rect 33836 59752 33842 59764
rect 43254 59752 43260 59764
rect 33836 59724 43260 59752
rect 33836 59712 33842 59724
rect 43254 59712 43260 59724
rect 43312 59712 43318 59764
rect 56226 59712 56232 59764
rect 56284 59752 56290 59764
rect 57425 59755 57483 59761
rect 57425 59752 57437 59755
rect 56284 59724 57437 59752
rect 56284 59712 56290 59724
rect 57425 59721 57437 59724
rect 57471 59721 57483 59755
rect 58250 59752 58256 59764
rect 58211 59724 58256 59752
rect 57425 59715 57483 59721
rect 58250 59712 58256 59724
rect 58308 59712 58314 59764
rect 25866 59684 25872 59696
rect 25827 59656 25872 59684
rect 25866 59644 25872 59656
rect 25924 59644 25930 59696
rect 26970 59644 26976 59696
rect 27028 59684 27034 59696
rect 30098 59684 30104 59696
rect 27028 59656 30104 59684
rect 27028 59644 27034 59656
rect 30098 59644 30104 59656
rect 30156 59644 30162 59696
rect 56410 59644 56416 59696
rect 56468 59684 56474 59696
rect 57333 59687 57391 59693
rect 57333 59684 57345 59687
rect 56468 59656 57345 59684
rect 56468 59644 56474 59656
rect 57333 59653 57345 59656
rect 57379 59653 57391 59687
rect 57333 59647 57391 59653
rect 25639 59588 25728 59616
rect 25639 59585 25651 59588
rect 25593 59579 25651 59585
rect 25774 59576 25780 59628
rect 25832 59616 25838 59628
rect 25966 59619 26024 59625
rect 25832 59588 25877 59616
rect 25832 59576 25838 59588
rect 25966 59585 25978 59619
rect 26012 59585 26024 59619
rect 25966 59579 26024 59585
rect 25976 59548 26004 59579
rect 26234 59576 26240 59628
rect 26292 59616 26298 59628
rect 30006 59616 30012 59628
rect 26292 59588 30012 59616
rect 26292 59576 26298 59588
rect 30006 59576 30012 59588
rect 30064 59576 30070 59628
rect 35526 59576 35532 59628
rect 35584 59616 35590 59628
rect 35584 59588 43208 59616
rect 35584 59576 35590 59588
rect 26142 59548 26148 59560
rect 19484 59520 24440 59548
rect 19484 59508 19490 59520
rect 21082 59480 21088 59492
rect 18984 59452 21088 59480
rect 21082 59440 21088 59452
rect 21140 59440 21146 59492
rect 1762 59412 1768 59424
rect 1723 59384 1768 59412
rect 1762 59372 1768 59384
rect 1820 59372 1826 59424
rect 2314 59372 2320 59424
rect 2372 59412 2378 59424
rect 2501 59415 2559 59421
rect 2501 59412 2513 59415
rect 2372 59384 2513 59412
rect 2372 59372 2378 59384
rect 2501 59381 2513 59384
rect 2547 59381 2559 59415
rect 2501 59375 2559 59381
rect 6822 59372 6828 59424
rect 6880 59412 6886 59424
rect 7101 59415 7159 59421
rect 7101 59412 7113 59415
rect 6880 59384 7113 59412
rect 6880 59372 6886 59384
rect 7101 59381 7113 59384
rect 7147 59381 7159 59415
rect 18506 59412 18512 59424
rect 18467 59384 18512 59412
rect 7101 59375 7159 59381
rect 18506 59372 18512 59384
rect 18564 59412 18570 59424
rect 19150 59412 19156 59424
rect 18564 59384 19156 59412
rect 18564 59372 18570 59384
rect 19150 59372 19156 59384
rect 19208 59372 19214 59424
rect 19242 59372 19248 59424
rect 19300 59412 19306 59424
rect 19337 59415 19395 59421
rect 19337 59412 19349 59415
rect 19300 59384 19349 59412
rect 19300 59372 19306 59384
rect 19337 59381 19349 59384
rect 19383 59381 19395 59415
rect 24412 59412 24440 59520
rect 25700 59520 26148 59548
rect 25130 59440 25136 59492
rect 25188 59480 25194 59492
rect 25590 59480 25596 59492
rect 25188 59452 25596 59480
rect 25188 59440 25194 59452
rect 25590 59440 25596 59452
rect 25648 59440 25654 59492
rect 25700 59412 25728 59520
rect 26142 59508 26148 59520
rect 26200 59508 26206 59560
rect 42702 59548 42708 59560
rect 42663 59520 42708 59548
rect 42702 59508 42708 59520
rect 42760 59508 42766 59560
rect 42794 59508 42800 59560
rect 42852 59548 42858 59560
rect 43073 59551 43131 59557
rect 43073 59548 43085 59551
rect 42852 59520 43085 59548
rect 42852 59508 42858 59520
rect 43073 59517 43085 59520
rect 43119 59517 43131 59551
rect 43180 59548 43208 59588
rect 43254 59576 43260 59628
rect 43312 59616 43318 59628
rect 43625 59619 43683 59625
rect 43312 59588 43357 59616
rect 43312 59576 43318 59588
rect 43625 59585 43637 59619
rect 43671 59616 43683 59619
rect 53098 59616 53104 59628
rect 43671 59588 53104 59616
rect 43671 59585 43683 59588
rect 43625 59579 43683 59585
rect 53098 59576 53104 59588
rect 53156 59576 53162 59628
rect 58158 59616 58164 59628
rect 58119 59588 58164 59616
rect 58158 59576 58164 59588
rect 58216 59576 58222 59628
rect 43533 59551 43591 59557
rect 43533 59548 43545 59551
rect 43180 59520 43545 59548
rect 43073 59511 43131 59517
rect 43533 59517 43545 59520
rect 43579 59517 43591 59551
rect 43533 59511 43591 59517
rect 25774 59440 25780 59492
rect 25832 59480 25838 59492
rect 56318 59480 56324 59492
rect 25832 59452 56324 59480
rect 25832 59440 25838 59452
rect 56318 59440 56324 59452
rect 56376 59440 56382 59492
rect 24412 59384 25728 59412
rect 19337 59375 19395 59381
rect 25958 59372 25964 59424
rect 26016 59412 26022 59424
rect 26145 59415 26203 59421
rect 26145 59412 26157 59415
rect 26016 59384 26157 59412
rect 26016 59372 26022 59384
rect 26145 59381 26157 59384
rect 26191 59381 26203 59415
rect 26145 59375 26203 59381
rect 27982 59372 27988 59424
rect 28040 59412 28046 59424
rect 28997 59415 29055 59421
rect 28997 59412 29009 59415
rect 28040 59384 29009 59412
rect 28040 59372 28046 59384
rect 28997 59381 29009 59384
rect 29043 59412 29055 59415
rect 29822 59412 29828 59424
rect 29043 59384 29828 59412
rect 29043 59381 29055 59384
rect 28997 59375 29055 59381
rect 29822 59372 29828 59384
rect 29880 59372 29886 59424
rect 30006 59372 30012 59424
rect 30064 59412 30070 59424
rect 55582 59412 55588 59424
rect 30064 59384 55588 59412
rect 30064 59372 30070 59384
rect 55582 59372 55588 59384
rect 55640 59372 55646 59424
rect 57146 59372 57152 59424
rect 57204 59412 57210 59424
rect 58986 59412 58992 59424
rect 57204 59384 58992 59412
rect 57204 59372 57210 59384
rect 58986 59372 58992 59384
rect 59044 59372 59050 59424
rect 1104 59322 58880 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 58880 59322
rect 1104 59248 58880 59270
rect 1762 59168 1768 59220
rect 1820 59208 1826 59220
rect 1820 59180 40632 59208
rect 1820 59168 1826 59180
rect 1857 59143 1915 59149
rect 1857 59109 1869 59143
rect 1903 59140 1915 59143
rect 5994 59140 6000 59152
rect 1903 59112 6000 59140
rect 1903 59109 1915 59112
rect 1857 59103 1915 59109
rect 5994 59100 6000 59112
rect 6052 59100 6058 59152
rect 26878 59032 26884 59084
rect 26936 59072 26942 59084
rect 40604 59081 40632 59180
rect 58342 59140 58348 59152
rect 45526 59112 58348 59140
rect 40589 59075 40647 59081
rect 26936 59044 37872 59072
rect 26936 59032 26942 59044
rect 842 58964 848 59016
rect 900 59004 906 59016
rect 1673 59007 1731 59013
rect 1673 59004 1685 59007
rect 900 58976 1685 59004
rect 900 58964 906 58976
rect 1673 58973 1685 58976
rect 1719 58973 1731 59007
rect 37182 59004 37188 59016
rect 37143 58976 37188 59004
rect 1673 58967 1731 58973
rect 37182 58964 37188 58976
rect 37240 58964 37246 59016
rect 37274 58964 37280 59016
rect 37332 59004 37338 59016
rect 37550 59004 37556 59016
rect 37332 58976 37377 59004
rect 37511 58976 37556 59004
rect 37332 58964 37338 58976
rect 37550 58964 37556 58976
rect 37608 58964 37614 59016
rect 37844 59013 37872 59044
rect 40589 59041 40601 59075
rect 40635 59041 40647 59075
rect 40589 59035 40647 59041
rect 41049 59075 41107 59081
rect 41049 59041 41061 59075
rect 41095 59072 41107 59075
rect 41095 59044 41414 59072
rect 41095 59041 41107 59044
rect 41049 59035 41107 59041
rect 41386 59016 41414 59044
rect 37829 59007 37887 59013
rect 37829 58973 37841 59007
rect 37875 58973 37887 59007
rect 37829 58967 37887 58973
rect 38105 59007 38163 59013
rect 38105 58973 38117 59007
rect 38151 58973 38163 59007
rect 40770 59004 40776 59016
rect 40731 58976 40776 59004
rect 38105 58967 38163 58973
rect 34514 58896 34520 58948
rect 34572 58936 34578 58948
rect 36725 58939 36783 58945
rect 36725 58936 36737 58939
rect 34572 58908 36737 58936
rect 34572 58896 34578 58908
rect 36725 58905 36737 58908
rect 36771 58905 36783 58939
rect 38120 58936 38148 58967
rect 40770 58964 40776 58976
rect 40828 58964 40834 59016
rect 41141 59007 41199 59013
rect 41141 58973 41153 59007
rect 41187 59004 41199 59007
rect 41230 59004 41236 59016
rect 41187 58976 41236 59004
rect 41187 58973 41199 58976
rect 41141 58967 41199 58973
rect 41230 58964 41236 58976
rect 41288 58964 41294 59016
rect 41386 59004 41420 59016
rect 41327 58976 41420 59004
rect 41414 58964 41420 58976
rect 41472 59004 41478 59016
rect 41874 59004 41880 59016
rect 41472 58976 41880 59004
rect 41472 58964 41478 58976
rect 41874 58964 41880 58976
rect 41932 58964 41938 59016
rect 45526 58936 45554 59112
rect 58342 59100 58348 59112
rect 58400 59100 58406 59152
rect 57146 59004 57152 59016
rect 57107 58976 57152 59004
rect 57146 58964 57152 58976
rect 57204 58964 57210 59016
rect 57882 59004 57888 59016
rect 57843 58976 57888 59004
rect 57882 58964 57888 58976
rect 57940 58964 57946 59016
rect 38120 58908 45554 58936
rect 58161 58939 58219 58945
rect 36725 58899 36783 58905
rect 58161 58905 58173 58939
rect 58207 58936 58219 58939
rect 58526 58936 58532 58948
rect 58207 58908 58532 58936
rect 58207 58905 58219 58908
rect 58161 58899 58219 58905
rect 58526 58896 58532 58908
rect 58584 58896 58590 58948
rect 40405 58871 40463 58877
rect 40405 58837 40417 58871
rect 40451 58868 40463 58871
rect 40862 58868 40868 58880
rect 40451 58840 40868 58868
rect 40451 58837 40463 58840
rect 40405 58831 40463 58837
rect 40862 58828 40868 58840
rect 40920 58828 40926 58880
rect 57330 58868 57336 58880
rect 57291 58840 57336 58868
rect 57330 58828 57336 58840
rect 57388 58828 57394 58880
rect 1104 58778 58880 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 58880 58778
rect 1104 58704 58880 58726
rect 18782 58624 18788 58676
rect 18840 58664 18846 58676
rect 57330 58664 57336 58676
rect 18840 58636 57336 58664
rect 18840 58624 18846 58636
rect 57330 58624 57336 58636
rect 57388 58624 57394 58676
rect 58158 58596 58164 58608
rect 58119 58568 58164 58596
rect 58158 58556 58164 58568
rect 58216 58556 58222 58608
rect 1578 58528 1584 58540
rect 1539 58500 1584 58528
rect 1578 58488 1584 58500
rect 1636 58488 1642 58540
rect 40589 58531 40647 58537
rect 40589 58528 40601 58531
rect 22066 58500 40601 58528
rect 1762 58460 1768 58472
rect 1723 58432 1768 58460
rect 1762 58420 1768 58432
rect 1820 58420 1826 58472
rect 2038 58420 2044 58472
rect 2096 58460 2102 58472
rect 22066 58460 22094 58500
rect 40589 58497 40601 58500
rect 40635 58497 40647 58531
rect 40589 58491 40647 58497
rect 40770 58488 40776 58540
rect 40828 58528 40834 58540
rect 41138 58528 41144 58540
rect 40828 58500 40921 58528
rect 41099 58500 41144 58528
rect 40828 58488 40834 58500
rect 41138 58488 41144 58500
rect 41196 58488 41202 58540
rect 41325 58531 41383 58537
rect 41325 58497 41337 58531
rect 41371 58528 41383 58531
rect 41414 58528 41420 58540
rect 41371 58500 41420 58528
rect 41371 58497 41383 58500
rect 41325 58491 41383 58497
rect 41414 58488 41420 58500
rect 41472 58488 41478 58540
rect 2096 58432 22094 58460
rect 2096 58420 2102 58432
rect 39298 58420 39304 58472
rect 39356 58460 39362 58472
rect 40788 58460 40816 58488
rect 39356 58432 40816 58460
rect 39356 58420 39362 58432
rect 40402 58324 40408 58336
rect 40363 58296 40408 58324
rect 40402 58284 40408 58296
rect 40460 58284 40466 58336
rect 56502 58284 56508 58336
rect 56560 58324 56566 58336
rect 58253 58327 58311 58333
rect 58253 58324 58265 58327
rect 56560 58296 58265 58324
rect 56560 58284 56566 58296
rect 58253 58293 58265 58296
rect 58299 58293 58311 58327
rect 58253 58287 58311 58293
rect 1104 58234 58880 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 58880 58234
rect 1104 58160 58880 58182
rect 52914 57944 52920 57996
rect 52972 57984 52978 57996
rect 58253 57987 58311 57993
rect 58253 57984 58265 57987
rect 52972 57956 58265 57984
rect 52972 57944 52978 57956
rect 58253 57953 58265 57956
rect 58299 57953 58311 57987
rect 58253 57947 58311 57953
rect 1578 57916 1584 57928
rect 1539 57888 1584 57916
rect 1578 57876 1584 57888
rect 1636 57876 1642 57928
rect 1857 57851 1915 57857
rect 1857 57817 1869 57851
rect 1903 57848 1915 57851
rect 17218 57848 17224 57860
rect 1903 57820 17224 57848
rect 1903 57817 1915 57820
rect 1857 57811 1915 57817
rect 17218 57808 17224 57820
rect 17276 57808 17282 57860
rect 57974 57848 57980 57860
rect 57935 57820 57980 57848
rect 57974 57808 57980 57820
rect 58032 57808 58038 57860
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1578 57440 1584 57452
rect 1539 57412 1584 57440
rect 1578 57400 1584 57412
rect 1636 57400 1642 57452
rect 1765 57239 1823 57245
rect 1765 57205 1777 57239
rect 1811 57236 1823 57239
rect 29638 57236 29644 57248
rect 1811 57208 29644 57236
rect 1811 57205 1823 57208
rect 1765 57199 1823 57205
rect 29638 57196 29644 57208
rect 29696 57196 29702 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 26970 56992 26976 57044
rect 27028 57032 27034 57044
rect 34514 57032 34520 57044
rect 27028 57004 34520 57032
rect 27028 56992 27034 57004
rect 34514 56992 34520 57004
rect 34572 56992 34578 57044
rect 28350 56924 28356 56976
rect 28408 56964 28414 56976
rect 35253 56967 35311 56973
rect 35253 56964 35265 56967
rect 28408 56936 35265 56964
rect 28408 56924 28414 56936
rect 35253 56933 35265 56936
rect 35299 56933 35311 56967
rect 52454 56964 52460 56976
rect 35253 56927 35311 56933
rect 35912 56936 36216 56964
rect 33965 56899 34023 56905
rect 33965 56865 33977 56899
rect 34011 56896 34023 56899
rect 35912 56896 35940 56936
rect 34011 56868 35940 56896
rect 34011 56865 34023 56868
rect 33965 56859 34023 56865
rect 1578 56828 1584 56840
rect 1539 56800 1584 56828
rect 1578 56788 1584 56800
rect 1636 56788 1642 56840
rect 22462 56788 22468 56840
rect 22520 56828 22526 56840
rect 33505 56831 33563 56837
rect 33505 56828 33517 56831
rect 22520 56800 33517 56828
rect 22520 56788 22526 56800
rect 33505 56797 33517 56800
rect 33551 56797 33563 56831
rect 33505 56791 33563 56797
rect 33689 56831 33747 56837
rect 33689 56797 33701 56831
rect 33735 56828 33747 56831
rect 33778 56828 33784 56840
rect 33735 56800 33784 56828
rect 33735 56797 33747 56800
rect 33689 56791 33747 56797
rect 33778 56788 33784 56800
rect 33836 56788 33842 56840
rect 25682 56720 25688 56772
rect 25740 56760 25746 56772
rect 33980 56760 34008 56859
rect 34057 56831 34115 56837
rect 34057 56797 34069 56831
rect 34103 56797 34115 56831
rect 34057 56791 34115 56797
rect 25740 56732 34008 56760
rect 25740 56720 25746 56732
rect 1765 56695 1823 56701
rect 1765 56661 1777 56695
rect 1811 56692 1823 56695
rect 27614 56692 27620 56704
rect 1811 56664 27620 56692
rect 1811 56661 1823 56664
rect 1765 56655 1823 56661
rect 27614 56652 27620 56664
rect 27672 56652 27678 56704
rect 33318 56692 33324 56704
rect 33279 56664 33324 56692
rect 33318 56652 33324 56664
rect 33376 56652 33382 56704
rect 34072 56692 34100 56791
rect 35618 56788 35624 56840
rect 35676 56828 35682 56840
rect 35894 56828 35900 56840
rect 35676 56800 35721 56828
rect 35855 56800 35900 56828
rect 35676 56788 35682 56800
rect 35894 56788 35900 56800
rect 35952 56788 35958 56840
rect 35986 56788 35992 56840
rect 36044 56828 36050 56840
rect 36188 56828 36216 56936
rect 36464 56936 52460 56964
rect 36265 56831 36323 56837
rect 36265 56828 36277 56831
rect 36044 56800 36089 56828
rect 36188 56800 36277 56828
rect 36044 56788 36050 56800
rect 36265 56797 36277 56800
rect 36311 56797 36323 56831
rect 36265 56791 36323 56797
rect 36464 56692 36492 56936
rect 52454 56924 52460 56936
rect 52512 56924 52518 56976
rect 56502 56896 56508 56908
rect 45526 56868 56508 56896
rect 36541 56831 36599 56837
rect 36541 56797 36553 56831
rect 36587 56828 36599 56831
rect 45526 56828 45554 56868
rect 56502 56856 56508 56868
rect 56560 56856 56566 56908
rect 57882 56828 57888 56840
rect 36587 56800 45554 56828
rect 57843 56800 57888 56828
rect 36587 56797 36599 56800
rect 36541 56791 36599 56797
rect 57882 56788 57888 56800
rect 57940 56788 57946 56840
rect 58066 56720 58072 56772
rect 58124 56760 58130 56772
rect 58161 56763 58219 56769
rect 58161 56760 58173 56763
rect 58124 56732 58173 56760
rect 58124 56720 58130 56732
rect 58161 56729 58173 56732
rect 58207 56729 58219 56763
rect 58161 56723 58219 56729
rect 34072 56664 36492 56692
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 35618 56448 35624 56500
rect 35676 56488 35682 56500
rect 36446 56488 36452 56500
rect 35676 56460 36452 56488
rect 35676 56448 35682 56460
rect 36446 56448 36452 56460
rect 36504 56488 36510 56500
rect 37182 56488 37188 56500
rect 36504 56460 37188 56488
rect 36504 56448 36510 56460
rect 37182 56448 37188 56460
rect 37240 56488 37246 56500
rect 41414 56488 41420 56500
rect 37240 56460 41420 56488
rect 37240 56448 37246 56460
rect 41414 56448 41420 56460
rect 41472 56448 41478 56500
rect 27614 56380 27620 56432
rect 27672 56420 27678 56432
rect 58158 56420 58164 56432
rect 27672 56392 41000 56420
rect 58119 56392 58164 56420
rect 27672 56380 27678 56392
rect 29270 56352 29276 56364
rect 29231 56324 29276 56352
rect 29270 56312 29276 56324
rect 29328 56312 29334 56364
rect 29638 56352 29644 56364
rect 29599 56324 29644 56352
rect 29638 56312 29644 56324
rect 29696 56312 29702 56364
rect 29825 56355 29883 56361
rect 29825 56321 29837 56355
rect 29871 56352 29883 56355
rect 30006 56352 30012 56364
rect 29871 56324 30012 56352
rect 29871 56321 29883 56324
rect 29825 56315 29883 56321
rect 30006 56312 30012 56324
rect 30064 56312 30070 56364
rect 35526 56312 35532 56364
rect 35584 56352 35590 56364
rect 35621 56355 35679 56361
rect 35621 56352 35633 56355
rect 35584 56324 35633 56352
rect 35584 56312 35590 56324
rect 35621 56321 35633 56324
rect 35667 56321 35679 56355
rect 36446 56352 36452 56364
rect 36407 56324 36452 56352
rect 35621 56315 35679 56321
rect 36446 56312 36452 56324
rect 36504 56312 36510 56364
rect 40972 56361 41000 56392
rect 58158 56380 58164 56392
rect 58216 56380 58222 56432
rect 40957 56355 41015 56361
rect 40957 56321 40969 56355
rect 41003 56321 41015 56355
rect 40957 56315 41015 56321
rect 41141 56355 41199 56361
rect 41141 56321 41153 56355
rect 41187 56321 41199 56355
rect 41141 56315 41199 56321
rect 41509 56355 41567 56361
rect 41509 56321 41521 56355
rect 41555 56352 41567 56355
rect 46750 56352 46756 56364
rect 41555 56324 46756 56352
rect 41555 56321 41567 56324
rect 41509 56315 41567 56321
rect 27338 56244 27344 56296
rect 27396 56284 27402 56296
rect 29181 56287 29239 56293
rect 29181 56284 29193 56287
rect 27396 56256 29193 56284
rect 27396 56244 27402 56256
rect 29181 56253 29193 56256
rect 29227 56253 29239 56287
rect 29181 56247 29239 56253
rect 39942 56244 39948 56296
rect 40000 56284 40006 56296
rect 41156 56284 41184 56315
rect 46750 56312 46756 56324
rect 46808 56312 46814 56364
rect 41414 56284 41420 56296
rect 40000 56256 41184 56284
rect 41375 56256 41420 56284
rect 40000 56244 40006 56256
rect 41414 56244 41420 56256
rect 41472 56244 41478 56296
rect 28721 56151 28779 56157
rect 28721 56117 28733 56151
rect 28767 56148 28779 56151
rect 32398 56148 32404 56160
rect 28767 56120 32404 56148
rect 28767 56117 28779 56120
rect 28721 56111 28779 56117
rect 32398 56108 32404 56120
rect 32456 56108 32462 56160
rect 40773 56151 40831 56157
rect 40773 56117 40785 56151
rect 40819 56148 40831 56151
rect 42242 56148 42248 56160
rect 40819 56120 42248 56148
rect 40819 56117 40831 56120
rect 40773 56111 40831 56117
rect 42242 56108 42248 56120
rect 42300 56108 42306 56160
rect 52454 56108 52460 56160
rect 52512 56148 52518 56160
rect 58253 56151 58311 56157
rect 58253 56148 58265 56151
rect 52512 56120 58265 56148
rect 52512 56108 52518 56120
rect 58253 56117 58265 56120
rect 58299 56117 58311 56151
rect 58253 56111 58311 56117
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 58342 55944 58348 55956
rect 58303 55916 58348 55944
rect 58342 55904 58348 55916
rect 58400 55904 58406 55956
rect 27522 55808 27528 55820
rect 27264 55780 27528 55808
rect 23566 55700 23572 55752
rect 23624 55740 23630 55752
rect 27264 55749 27292 55780
rect 27522 55768 27528 55780
rect 27580 55768 27586 55820
rect 27249 55743 27307 55749
rect 23624 55712 26740 55740
rect 23624 55700 23630 55712
rect 1670 55672 1676 55684
rect 1631 55644 1676 55672
rect 1670 55632 1676 55644
rect 1728 55632 1734 55684
rect 26602 55672 26608 55684
rect 26563 55644 26608 55672
rect 26602 55632 26608 55644
rect 26660 55632 26666 55684
rect 26712 55672 26740 55712
rect 27249 55709 27261 55743
rect 27295 55709 27307 55743
rect 27249 55703 27307 55709
rect 27338 55700 27344 55752
rect 27396 55740 27402 55752
rect 27617 55743 27675 55749
rect 27396 55712 27441 55740
rect 27396 55700 27402 55712
rect 27617 55709 27629 55743
rect 27663 55709 27675 55743
rect 27617 55703 27675 55709
rect 27801 55743 27859 55749
rect 27801 55709 27813 55743
rect 27847 55740 27859 55743
rect 30006 55740 30012 55752
rect 27847 55712 30012 55740
rect 27847 55709 27859 55712
rect 27801 55703 27859 55709
rect 27356 55672 27384 55700
rect 26712 55644 27384 55672
rect 1765 55607 1823 55613
rect 1765 55573 1777 55607
rect 1811 55604 1823 55607
rect 27632 55604 27660 55703
rect 30006 55700 30012 55712
rect 30064 55700 30070 55752
rect 1811 55576 27660 55604
rect 1811 55573 1823 55576
rect 1765 55567 1823 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1765 55403 1823 55409
rect 1765 55369 1777 55403
rect 1811 55400 1823 55403
rect 1811 55372 6914 55400
rect 1811 55369 1823 55372
rect 1765 55363 1823 55369
rect 6886 55332 6914 55372
rect 6886 55304 22094 55332
rect 1578 55264 1584 55276
rect 1539 55236 1584 55264
rect 1578 55224 1584 55236
rect 1636 55224 1642 55276
rect 22066 55264 22094 55304
rect 39390 55292 39396 55344
rect 39448 55332 39454 55344
rect 39942 55332 39948 55344
rect 39448 55304 39948 55332
rect 39448 55292 39454 55304
rect 39942 55292 39948 55304
rect 40000 55332 40006 55344
rect 41414 55332 41420 55344
rect 40000 55304 40632 55332
rect 40000 55292 40006 55304
rect 40604 55273 40632 55304
rect 40880 55304 41420 55332
rect 40405 55267 40463 55273
rect 40405 55264 40417 55267
rect 22066 55236 40417 55264
rect 40405 55233 40417 55236
rect 40451 55233 40463 55267
rect 40405 55227 40463 55233
rect 40589 55267 40647 55273
rect 40589 55233 40601 55267
rect 40635 55233 40647 55267
rect 40589 55227 40647 55233
rect 40034 55196 40040 55208
rect 39995 55168 40040 55196
rect 40034 55156 40040 55168
rect 40092 55156 40098 55208
rect 40880 55205 40908 55304
rect 41414 55292 41420 55304
rect 41472 55292 41478 55344
rect 40957 55267 41015 55273
rect 40957 55233 40969 55267
rect 41003 55264 41015 55267
rect 44174 55264 44180 55276
rect 41003 55236 44180 55264
rect 41003 55233 41015 55236
rect 40957 55227 41015 55233
rect 44174 55224 44180 55236
rect 44232 55224 44238 55276
rect 40865 55199 40923 55205
rect 40865 55165 40877 55199
rect 40911 55165 40923 55199
rect 40865 55159 40923 55165
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 18046 54680 18052 54732
rect 18104 54720 18110 54732
rect 23566 54720 23572 54732
rect 18104 54692 23572 54720
rect 18104 54680 18110 54692
rect 23566 54680 23572 54692
rect 23624 54680 23630 54732
rect 26050 54720 26056 54732
rect 23768 54692 26056 54720
rect 23477 54655 23535 54661
rect 23477 54621 23489 54655
rect 23523 54652 23535 54655
rect 23768 54652 23796 54692
rect 26050 54680 26056 54692
rect 26108 54680 26114 54732
rect 23523 54624 23796 54652
rect 23845 54655 23903 54661
rect 23523 54621 23535 54624
rect 23477 54615 23535 54621
rect 23845 54621 23857 54655
rect 23891 54621 23903 54655
rect 23845 54615 23903 54621
rect 1670 54584 1676 54596
rect 1631 54556 1676 54584
rect 1670 54544 1676 54556
rect 1728 54544 1734 54596
rect 22830 54584 22836 54596
rect 22791 54556 22836 54584
rect 22830 54544 22836 54556
rect 22888 54544 22894 54596
rect 1765 54519 1823 54525
rect 1765 54485 1777 54519
rect 1811 54516 1823 54519
rect 23860 54516 23888 54615
rect 23934 54612 23940 54664
rect 23992 54652 23998 54664
rect 24029 54655 24087 54661
rect 24029 54652 24041 54655
rect 23992 54624 24041 54652
rect 23992 54612 23998 54624
rect 24029 54621 24041 54624
rect 24075 54652 24087 54655
rect 30006 54652 30012 54664
rect 24075 54624 30012 54652
rect 24075 54621 24087 54624
rect 24029 54615 24087 54621
rect 30006 54612 30012 54624
rect 30064 54612 30070 54664
rect 58342 54652 58348 54664
rect 58303 54624 58348 54652
rect 58342 54612 58348 54624
rect 58400 54612 58406 54664
rect 1811 54488 23888 54516
rect 1811 54485 1823 54488
rect 1765 54479 1823 54485
rect 27522 54476 27528 54528
rect 27580 54516 27586 54528
rect 45370 54516 45376 54528
rect 27580 54488 45376 54516
rect 27580 54476 27586 54488
rect 45370 54476 45376 54488
rect 45428 54476 45434 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1578 54176 1584 54188
rect 1539 54148 1584 54176
rect 1578 54136 1584 54148
rect 1636 54136 1642 54188
rect 1765 53975 1823 53981
rect 1765 53941 1777 53975
rect 1811 53972 1823 53975
rect 10962 53972 10968 53984
rect 1811 53944 10968 53972
rect 1811 53941 1823 53944
rect 1765 53935 1823 53941
rect 10962 53932 10968 53944
rect 11020 53932 11026 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 40862 53660 40868 53712
rect 40920 53700 40926 53712
rect 41874 53700 41880 53712
rect 40920 53672 41880 53700
rect 40920 53660 40926 53672
rect 41874 53660 41880 53672
rect 41932 53660 41938 53712
rect 10962 53592 10968 53644
rect 11020 53632 11026 53644
rect 40497 53635 40555 53641
rect 40497 53632 40509 53635
rect 11020 53604 40509 53632
rect 11020 53592 11026 53604
rect 40497 53601 40509 53604
rect 40543 53601 40555 53635
rect 46106 53632 46112 53644
rect 40497 53595 40555 53601
rect 41064 53604 46112 53632
rect 30006 53524 30012 53576
rect 30064 53564 30070 53576
rect 36446 53564 36452 53576
rect 30064 53536 36452 53564
rect 30064 53524 30070 53536
rect 36446 53524 36452 53536
rect 36504 53564 36510 53576
rect 41064 53573 41092 53604
rect 46106 53592 46112 53604
rect 46164 53592 46170 53644
rect 40681 53567 40739 53573
rect 40681 53564 40693 53567
rect 36504 53536 40693 53564
rect 36504 53524 36510 53536
rect 40681 53533 40693 53536
rect 40727 53533 40739 53567
rect 40681 53527 40739 53533
rect 41049 53567 41107 53573
rect 41049 53533 41061 53567
rect 41095 53533 41107 53567
rect 41049 53527 41107 53533
rect 41233 53567 41291 53573
rect 41233 53533 41245 53567
rect 41279 53564 41291 53567
rect 41414 53564 41420 53576
rect 41279 53536 41420 53564
rect 41279 53533 41291 53536
rect 41233 53527 41291 53533
rect 41414 53524 41420 53536
rect 41472 53524 41478 53576
rect 40313 53431 40371 53437
rect 40313 53397 40325 53431
rect 40359 53428 40371 53431
rect 40402 53428 40408 53440
rect 40359 53400 40408 53428
rect 40359 53397 40371 53400
rect 40313 53391 40371 53397
rect 40402 53388 40408 53400
rect 40460 53388 40466 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 23934 53224 23940 53236
rect 23308 53196 23940 53224
rect 23308 53165 23336 53196
rect 23934 53184 23940 53196
rect 23992 53184 23998 53236
rect 23293 53159 23351 53165
rect 23293 53125 23305 53159
rect 23339 53125 23351 53159
rect 23293 53119 23351 53125
rect 23385 53159 23443 53165
rect 23385 53125 23397 53159
rect 23431 53156 23443 53159
rect 27522 53156 27528 53168
rect 23431 53128 27528 53156
rect 23431 53125 23443 53128
rect 23385 53119 23443 53125
rect 27522 53116 27528 53128
rect 27580 53116 27586 53168
rect 1670 53088 1676 53100
rect 1631 53060 1676 53088
rect 1670 53048 1676 53060
rect 1728 53048 1734 53100
rect 23109 53091 23167 53097
rect 23109 53088 23121 53091
rect 6886 53060 23121 53088
rect 1765 52887 1823 52893
rect 1765 52853 1777 52887
rect 1811 52884 1823 52887
rect 6886 52884 6914 53060
rect 23109 53057 23121 53060
rect 23155 53057 23167 53091
rect 23109 53051 23167 53057
rect 23529 53091 23587 53097
rect 23529 53057 23541 53091
rect 23575 53088 23587 53091
rect 23842 53088 23848 53100
rect 23575 53060 23848 53088
rect 23575 53057 23587 53060
rect 23529 53051 23587 53057
rect 23842 53048 23848 53060
rect 23900 53088 23906 53100
rect 24302 53088 24308 53100
rect 23900 53060 24164 53088
rect 24263 53060 24308 53088
rect 23900 53048 23906 53060
rect 24136 53020 24164 53060
rect 24302 53048 24308 53060
rect 24360 53048 24366 53100
rect 27430 53048 27436 53100
rect 27488 53088 27494 53100
rect 39666 53088 39672 53100
rect 27488 53060 39672 53088
rect 27488 53048 27494 53060
rect 39666 53048 39672 53060
rect 39724 53048 39730 53100
rect 24581 53023 24639 53029
rect 24581 53020 24593 53023
rect 24136 52992 24593 53020
rect 24581 52989 24593 52992
rect 24627 52989 24639 53023
rect 24581 52983 24639 52989
rect 1811 52856 6914 52884
rect 1811 52853 1823 52856
rect 1765 52847 1823 52853
rect 23566 52844 23572 52896
rect 23624 52884 23630 52896
rect 23661 52887 23719 52893
rect 23661 52884 23673 52887
rect 23624 52856 23673 52884
rect 23624 52844 23630 52856
rect 23661 52853 23673 52856
rect 23707 52853 23719 52887
rect 58342 52884 58348 52896
rect 58303 52856 58348 52884
rect 23661 52847 23719 52853
rect 58342 52844 58348 52856
rect 58400 52844 58406 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1854 52544 1860 52556
rect 1815 52516 1860 52544
rect 1854 52504 1860 52516
rect 1912 52504 1918 52556
rect 34606 52504 34612 52556
rect 34664 52544 34670 52556
rect 35986 52544 35992 52556
rect 34664 52516 35992 52544
rect 34664 52504 34670 52516
rect 35986 52504 35992 52516
rect 36044 52504 36050 52556
rect 1578 52476 1584 52488
rect 1539 52448 1584 52476
rect 1578 52436 1584 52448
rect 1636 52436 1642 52488
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1857 52071 1915 52077
rect 1857 52037 1869 52071
rect 1903 52068 1915 52071
rect 7009 52071 7067 52077
rect 7009 52068 7021 52071
rect 1903 52040 7021 52068
rect 1903 52037 1915 52040
rect 1857 52031 1915 52037
rect 7009 52037 7021 52040
rect 7055 52037 7067 52071
rect 7009 52031 7067 52037
rect 1670 52000 1676 52012
rect 1631 51972 1676 52000
rect 1670 51960 1676 51972
rect 1728 51960 1734 52012
rect 6822 52000 6828 52012
rect 6783 51972 6828 52000
rect 6822 51960 6828 51972
rect 6880 51960 6886 52012
rect 7098 52000 7104 52012
rect 7059 51972 7104 52000
rect 7098 51960 7104 51972
rect 7156 51960 7162 52012
rect 6641 51799 6699 51805
rect 6641 51765 6653 51799
rect 6687 51796 6699 51799
rect 6730 51796 6736 51808
rect 6687 51768 6736 51796
rect 6687 51765 6699 51768
rect 6641 51759 6699 51765
rect 6730 51756 6736 51768
rect 6788 51756 6794 51808
rect 17310 51756 17316 51808
rect 17368 51796 17374 51808
rect 26326 51796 26332 51808
rect 17368 51768 26332 51796
rect 17368 51756 17374 51768
rect 26326 51756 26332 51768
rect 26384 51756 26390 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58342 51388 58348 51400
rect 58303 51360 58348 51388
rect 58342 51348 58348 51360
rect 58400 51348 58406 51400
rect 1670 51320 1676 51332
rect 1631 51292 1676 51320
rect 1670 51280 1676 51292
rect 1728 51280 1734 51332
rect 1857 51323 1915 51329
rect 1857 51289 1869 51323
rect 1903 51320 1915 51323
rect 3970 51320 3976 51332
rect 1903 51292 3976 51320
rect 1903 51289 1915 51292
rect 1857 51283 1915 51289
rect 3970 51280 3976 51292
rect 4028 51280 4034 51332
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 4614 51048 4620 51060
rect 3712 51020 4620 51048
rect 3712 50921 3740 51020
rect 4614 51008 4620 51020
rect 4672 51008 4678 51060
rect 3970 50980 3976 50992
rect 3931 50952 3976 50980
rect 3970 50940 3976 50952
rect 4028 50940 4034 50992
rect 3697 50915 3755 50921
rect 3697 50881 3709 50915
rect 3743 50881 3755 50915
rect 3697 50875 3755 50881
rect 3878 50872 3884 50924
rect 3936 50912 3942 50924
rect 4117 50915 4175 50921
rect 3936 50884 4029 50912
rect 3936 50872 3942 50884
rect 4117 50881 4129 50915
rect 4163 50912 4175 50915
rect 7098 50912 7104 50924
rect 4163 50884 7104 50912
rect 4163 50881 4175 50884
rect 4117 50875 4175 50881
rect 7098 50872 7104 50884
rect 7156 50912 7162 50924
rect 7558 50912 7564 50924
rect 7156 50884 7564 50912
rect 7156 50872 7162 50884
rect 7558 50872 7564 50884
rect 7616 50872 7622 50924
rect 2590 50804 2596 50856
rect 2648 50844 2654 50856
rect 3896 50844 3924 50872
rect 2648 50816 3924 50844
rect 2648 50804 2654 50816
rect 4249 50711 4307 50717
rect 4249 50677 4261 50711
rect 4295 50708 4307 50711
rect 5902 50708 5908 50720
rect 4295 50680 5908 50708
rect 4295 50677 4307 50680
rect 4249 50671 4307 50677
rect 5902 50668 5908 50680
rect 5960 50668 5966 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 24210 50328 24216 50380
rect 24268 50368 24274 50380
rect 39298 50368 39304 50380
rect 24268 50340 39304 50368
rect 24268 50328 24274 50340
rect 39298 50328 39304 50340
rect 39356 50328 39362 50380
rect 45002 50260 45008 50312
rect 45060 50300 45066 50312
rect 57885 50303 57943 50309
rect 57885 50300 57897 50303
rect 45060 50272 57897 50300
rect 45060 50260 45066 50272
rect 57885 50269 57897 50272
rect 57931 50269 57943 50303
rect 57885 50263 57943 50269
rect 1670 50232 1676 50244
rect 1631 50204 1676 50232
rect 1670 50192 1676 50204
rect 1728 50192 1734 50244
rect 1857 50235 1915 50241
rect 1857 50201 1869 50235
rect 1903 50232 1915 50235
rect 2038 50232 2044 50244
rect 1903 50204 2044 50232
rect 1903 50201 1915 50204
rect 1857 50195 1915 50201
rect 2038 50192 2044 50204
rect 2096 50192 2102 50244
rect 58161 50235 58219 50241
rect 58161 50232 58173 50235
rect 57900 50204 58173 50232
rect 57900 50176 57928 50204
rect 58161 50201 58173 50204
rect 58207 50201 58219 50235
rect 58161 50195 58219 50201
rect 57882 50124 57888 50176
rect 57940 50124 57946 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1578 49824 1584 49836
rect 1539 49796 1584 49824
rect 1578 49784 1584 49796
rect 1636 49784 1642 49836
rect 22278 49756 22284 49768
rect 1780 49728 22284 49756
rect 1780 49697 1808 49728
rect 22278 49716 22284 49728
rect 22336 49716 22342 49768
rect 1765 49691 1823 49697
rect 1765 49657 1777 49691
rect 1811 49657 1823 49691
rect 1765 49651 1823 49657
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1670 49144 1676 49156
rect 1631 49116 1676 49144
rect 1670 49104 1676 49116
rect 1728 49104 1734 49156
rect 7834 49104 7840 49156
rect 7892 49144 7898 49156
rect 34790 49144 34796 49156
rect 7892 49116 34796 49144
rect 7892 49104 7898 49116
rect 34790 49104 34796 49116
rect 34848 49104 34854 49156
rect 41782 49104 41788 49156
rect 41840 49144 41846 49156
rect 54570 49144 54576 49156
rect 41840 49116 54576 49144
rect 41840 49104 41846 49116
rect 54570 49104 54576 49116
rect 54628 49104 54634 49156
rect 57974 49144 57980 49156
rect 57935 49116 57980 49144
rect 57974 49104 57980 49116
rect 58032 49104 58038 49156
rect 1765 49079 1823 49085
rect 1765 49045 1777 49079
rect 1811 49076 1823 49079
rect 15838 49076 15844 49088
rect 1811 49048 15844 49076
rect 1811 49045 1823 49048
rect 1765 49039 1823 49045
rect 15838 49036 15844 49048
rect 15896 49036 15902 49088
rect 51902 49036 51908 49088
rect 51960 49076 51966 49088
rect 58069 49079 58127 49085
rect 58069 49076 58081 49079
rect 51960 49048 58081 49076
rect 51960 49036 51966 49048
rect 58069 49045 58081 49048
rect 58115 49045 58127 49079
rect 58069 49039 58127 49045
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1670 48736 1676 48748
rect 1631 48708 1676 48736
rect 1670 48696 1676 48708
rect 1728 48696 1734 48748
rect 1857 48603 1915 48609
rect 1857 48569 1869 48603
rect 1903 48600 1915 48603
rect 1946 48600 1952 48612
rect 1903 48572 1952 48600
rect 1903 48569 1915 48572
rect 1857 48563 1915 48569
rect 1946 48560 1952 48572
rect 2004 48560 2010 48612
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 24762 48220 24768 48272
rect 24820 48260 24826 48272
rect 25406 48260 25412 48272
rect 24820 48232 25412 48260
rect 24820 48220 24826 48232
rect 25406 48220 25412 48232
rect 25464 48220 25470 48272
rect 56965 48127 57023 48133
rect 56965 48124 56977 48127
rect 56612 48096 56977 48124
rect 36262 47948 36268 48000
rect 36320 47988 36326 48000
rect 56612 47997 56640 48096
rect 56965 48093 56977 48096
rect 57011 48093 57023 48127
rect 56965 48087 57023 48093
rect 57238 48056 57244 48068
rect 57199 48028 57244 48056
rect 57238 48016 57244 48028
rect 57296 48016 57302 48068
rect 57974 48056 57980 48068
rect 57935 48028 57980 48056
rect 57974 48016 57980 48028
rect 58032 48016 58038 48068
rect 56597 47991 56655 47997
rect 56597 47988 56609 47991
rect 36320 47960 56609 47988
rect 36320 47948 36326 47960
rect 56597 47957 56609 47960
rect 56643 47957 56655 47991
rect 58066 47988 58072 48000
rect 58027 47960 58072 47988
rect 56597 47951 56655 47957
rect 58066 47948 58072 47960
rect 58124 47948 58130 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 46290 47744 46296 47796
rect 46348 47784 46354 47796
rect 58066 47784 58072 47796
rect 46348 47756 58072 47784
rect 46348 47744 46354 47756
rect 58066 47744 58072 47756
rect 58124 47744 58130 47796
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 3326 47540 3332 47592
rect 3384 47580 3390 47592
rect 20254 47580 20260 47592
rect 3384 47552 20260 47580
rect 3384 47540 3390 47552
rect 20254 47540 20260 47552
rect 20312 47540 20318 47592
rect 22186 47540 22192 47592
rect 22244 47580 22250 47592
rect 39390 47580 39396 47592
rect 22244 47552 39396 47580
rect 22244 47540 22250 47552
rect 39390 47540 39396 47552
rect 39448 47540 39454 47592
rect 1857 47515 1915 47521
rect 1857 47481 1869 47515
rect 1903 47512 1915 47515
rect 5442 47512 5448 47524
rect 1903 47484 5448 47512
rect 1903 47481 1915 47484
rect 1857 47475 1915 47481
rect 5442 47472 5448 47484
rect 5500 47472 5506 47524
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1578 47036 1584 47048
rect 1539 47008 1584 47036
rect 1578 46996 1584 47008
rect 1636 46996 1642 47048
rect 57514 46996 57520 47048
rect 57572 47036 57578 47048
rect 57885 47039 57943 47045
rect 57885 47036 57897 47039
rect 57572 47008 57897 47036
rect 57572 46996 57578 47008
rect 57885 47005 57897 47008
rect 57931 47005 57943 47039
rect 57885 46999 57943 47005
rect 24854 46968 24860 46980
rect 1780 46940 24860 46968
rect 1780 46909 1808 46940
rect 24854 46928 24860 46940
rect 24912 46928 24918 46980
rect 58161 46971 58219 46977
rect 58161 46968 58173 46971
rect 57900 46940 58173 46968
rect 57900 46912 57928 46940
rect 58161 46937 58173 46940
rect 58207 46937 58219 46971
rect 58161 46931 58219 46937
rect 1765 46903 1823 46909
rect 1765 46869 1777 46903
rect 1811 46869 1823 46903
rect 1765 46863 1823 46869
rect 57882 46860 57888 46912
rect 57940 46860 57946 46912
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1578 46560 1584 46572
rect 1539 46532 1584 46560
rect 1578 46520 1584 46532
rect 1636 46520 1642 46572
rect 19058 46384 19064 46436
rect 19116 46424 19122 46436
rect 39114 46424 39120 46436
rect 19116 46396 39120 46424
rect 19116 46384 19122 46396
rect 39114 46384 39120 46396
rect 39172 46384 39178 46436
rect 1765 46359 1823 46365
rect 1765 46325 1777 46359
rect 1811 46356 1823 46359
rect 20714 46356 20720 46368
rect 1811 46328 20720 46356
rect 1811 46325 1823 46328
rect 1765 46319 1823 46325
rect 20714 46316 20720 46328
rect 20772 46316 20778 46368
rect 34238 46316 34244 46368
rect 34296 46356 34302 46368
rect 54846 46356 54852 46368
rect 34296 46328 54852 46356
rect 34296 46316 34302 46328
rect 54846 46316 54852 46328
rect 54904 46316 54910 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1670 45880 1676 45892
rect 1631 45852 1676 45880
rect 1670 45840 1676 45852
rect 1728 45840 1734 45892
rect 57974 45880 57980 45892
rect 57935 45852 57980 45880
rect 57974 45840 57980 45852
rect 58032 45840 58038 45892
rect 1765 45815 1823 45821
rect 1765 45781 1777 45815
rect 1811 45812 1823 45815
rect 17678 45812 17684 45824
rect 1811 45784 17684 45812
rect 1811 45781 1823 45784
rect 1765 45775 1823 45781
rect 17678 45772 17684 45784
rect 17736 45772 17742 45824
rect 44910 45772 44916 45824
rect 44968 45812 44974 45824
rect 58069 45815 58127 45821
rect 58069 45812 58081 45815
rect 44968 45784 58081 45812
rect 44968 45772 44974 45784
rect 58069 45781 58081 45784
rect 58115 45781 58127 45815
rect 58069 45775 58127 45781
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 17862 45568 17868 45620
rect 17920 45608 17926 45620
rect 17920 45580 18000 45608
rect 17920 45568 17926 45580
rect 17770 45540 17776 45552
rect 17604 45512 17776 45540
rect 7558 45432 7564 45484
rect 7616 45472 7622 45484
rect 17604 45481 17632 45512
rect 17770 45500 17776 45512
rect 17828 45500 17834 45552
rect 17972 45549 18000 45580
rect 17957 45543 18015 45549
rect 17957 45509 17969 45543
rect 18003 45509 18015 45543
rect 17957 45503 18015 45509
rect 19720 45512 19932 45540
rect 17589 45475 17647 45481
rect 7616 45444 9674 45472
rect 7616 45432 7622 45444
rect 9646 45336 9674 45444
rect 17589 45441 17601 45475
rect 17635 45441 17647 45475
rect 17589 45435 17647 45441
rect 17678 45432 17684 45484
rect 17736 45472 17742 45484
rect 17865 45475 17923 45481
rect 17736 45444 17781 45472
rect 17736 45432 17742 45444
rect 17865 45441 17877 45475
rect 17911 45441 17923 45475
rect 17865 45435 17923 45441
rect 18095 45475 18153 45481
rect 18095 45441 18107 45475
rect 18141 45472 18153 45475
rect 18230 45472 18236 45484
rect 18141 45444 18236 45472
rect 18141 45441 18153 45444
rect 18095 45435 18153 45441
rect 17880 45336 17908 45435
rect 18230 45432 18236 45444
rect 18288 45432 18294 45484
rect 19720 45404 19748 45512
rect 19904 45472 19932 45512
rect 20714 45500 20720 45552
rect 20772 45540 20778 45552
rect 36541 45543 36599 45549
rect 20772 45512 26234 45540
rect 20772 45500 20778 45512
rect 24118 45472 24124 45484
rect 19904 45444 24124 45472
rect 24118 45432 24124 45444
rect 24176 45432 24182 45484
rect 26206 45472 26234 45512
rect 36541 45509 36553 45543
rect 36587 45540 36599 45543
rect 39850 45540 39856 45552
rect 36587 45512 39856 45540
rect 36587 45509 36599 45512
rect 36541 45503 36599 45509
rect 39850 45500 39856 45512
rect 39908 45500 39914 45552
rect 36265 45475 36323 45481
rect 36265 45472 36277 45475
rect 26206 45444 36277 45472
rect 36265 45441 36277 45444
rect 36311 45441 36323 45475
rect 36446 45472 36452 45484
rect 36407 45444 36452 45472
rect 36265 45435 36323 45441
rect 36446 45432 36452 45444
rect 36504 45432 36510 45484
rect 36685 45475 36743 45481
rect 36685 45441 36697 45475
rect 36731 45472 36743 45475
rect 37090 45472 37096 45484
rect 36731 45444 37096 45472
rect 36731 45441 36743 45444
rect 36685 45435 36743 45441
rect 37090 45432 37096 45444
rect 37148 45432 37154 45484
rect 19444 45376 19748 45404
rect 19444 45336 19472 45376
rect 9646 45308 19472 45336
rect 19794 45296 19800 45348
rect 19852 45336 19858 45348
rect 30558 45336 30564 45348
rect 19852 45308 30564 45336
rect 19852 45296 19858 45308
rect 30558 45296 30564 45308
rect 30616 45296 30622 45348
rect 36817 45339 36875 45345
rect 36817 45305 36829 45339
rect 36863 45336 36875 45339
rect 37550 45336 37556 45348
rect 36863 45308 37556 45336
rect 36863 45305 36875 45308
rect 36817 45299 36875 45305
rect 37550 45296 37556 45308
rect 37608 45296 37614 45348
rect 18230 45268 18236 45280
rect 18191 45240 18236 45268
rect 18230 45228 18236 45240
rect 18288 45228 18294 45280
rect 18322 45228 18328 45280
rect 18380 45268 18386 45280
rect 20806 45268 20812 45280
rect 18380 45240 20812 45268
rect 18380 45228 18386 45240
rect 20806 45228 20812 45240
rect 20864 45268 20870 45280
rect 21174 45268 21180 45280
rect 20864 45240 21180 45268
rect 20864 45228 20870 45240
rect 21174 45228 21180 45240
rect 21232 45228 21238 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 17770 45024 17776 45076
rect 17828 45064 17834 45076
rect 19794 45064 19800 45076
rect 17828 45036 19800 45064
rect 17828 45024 17834 45036
rect 19794 45024 19800 45036
rect 19852 45024 19858 45076
rect 30558 45024 30564 45076
rect 30616 45064 30622 45076
rect 38197 45067 38255 45073
rect 38197 45064 38209 45067
rect 30616 45036 38209 45064
rect 30616 45024 30622 45036
rect 38197 45033 38209 45036
rect 38243 45033 38255 45067
rect 38197 45027 38255 45033
rect 57054 44928 57060 44940
rect 37936 44900 57060 44928
rect 1578 44860 1584 44872
rect 1539 44832 1584 44860
rect 1578 44820 1584 44832
rect 1636 44820 1642 44872
rect 22830 44820 22836 44872
rect 22888 44860 22894 44872
rect 30742 44860 30748 44872
rect 22888 44832 30748 44860
rect 22888 44820 22894 44832
rect 30742 44820 30748 44832
rect 30800 44820 30806 44872
rect 37642 44860 37648 44872
rect 37603 44832 37648 44860
rect 37642 44820 37648 44832
rect 37700 44820 37706 44872
rect 37936 44869 37964 44900
rect 57054 44888 57060 44900
rect 57112 44888 57118 44940
rect 37921 44863 37979 44869
rect 37921 44829 37933 44863
rect 37967 44829 37979 44863
rect 37921 44823 37979 44829
rect 38018 44863 38076 44869
rect 38018 44829 38030 44863
rect 38064 44829 38076 44863
rect 38018 44823 38076 44829
rect 1857 44795 1915 44801
rect 1857 44761 1869 44795
rect 1903 44792 1915 44795
rect 31018 44792 31024 44804
rect 1903 44764 31024 44792
rect 1903 44761 1915 44764
rect 1857 44755 1915 44761
rect 31018 44752 31024 44764
rect 31076 44752 31082 44804
rect 37090 44752 37096 44804
rect 37148 44792 37154 44804
rect 37829 44795 37887 44801
rect 37829 44792 37841 44795
rect 37148 44764 37841 44792
rect 37148 44752 37154 44764
rect 37829 44761 37841 44764
rect 37875 44761 37887 44795
rect 37829 44755 37887 44761
rect 37366 44684 37372 44736
rect 37424 44724 37430 44736
rect 38028 44724 38056 44823
rect 50890 44820 50896 44872
rect 50948 44860 50954 44872
rect 56965 44863 57023 44869
rect 56965 44860 56977 44863
rect 50948 44832 56977 44860
rect 50948 44820 50954 44832
rect 56965 44829 56977 44832
rect 57011 44829 57023 44863
rect 56965 44823 57023 44829
rect 57238 44792 57244 44804
rect 57199 44764 57244 44792
rect 57238 44752 57244 44764
rect 57296 44752 57302 44804
rect 57882 44752 57888 44804
rect 57940 44792 57946 44804
rect 57977 44795 58035 44801
rect 57977 44792 57989 44795
rect 57940 44764 57989 44792
rect 57940 44752 57946 44764
rect 57977 44761 57989 44764
rect 58023 44761 58035 44795
rect 57977 44755 58035 44761
rect 58250 44724 58256 44736
rect 37424 44696 38056 44724
rect 58211 44696 58256 44724
rect 37424 44684 37430 44696
rect 58250 44684 58256 44696
rect 58308 44684 58314 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1670 44384 1676 44396
rect 1631 44356 1676 44384
rect 1670 44344 1676 44356
rect 1728 44344 1734 44396
rect 1765 44183 1823 44189
rect 1765 44149 1777 44183
rect 1811 44180 1823 44183
rect 17126 44180 17132 44192
rect 1811 44152 17132 44180
rect 1811 44149 1823 44152
rect 1765 44143 1823 44149
rect 17126 44140 17132 44152
rect 17184 44140 17190 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 35434 43908 35440 43920
rect 35395 43880 35440 43908
rect 35434 43868 35440 43880
rect 35492 43868 35498 43920
rect 17126 43800 17132 43852
rect 17184 43840 17190 43852
rect 35805 43843 35863 43849
rect 35805 43840 35817 43843
rect 17184 43812 35817 43840
rect 17184 43800 17190 43812
rect 34900 43781 34928 43812
rect 35805 43809 35817 43812
rect 35851 43809 35863 43843
rect 35805 43803 35863 43809
rect 34885 43775 34943 43781
rect 34885 43741 34897 43775
rect 34931 43741 34943 43775
rect 34885 43735 34943 43741
rect 35305 43775 35363 43781
rect 35305 43741 35317 43775
rect 35351 43772 35363 43775
rect 35351 43744 35894 43772
rect 35351 43741 35363 43744
rect 35305 43735 35363 43741
rect 1670 43704 1676 43716
rect 1631 43676 1676 43704
rect 1670 43664 1676 43676
rect 1728 43664 1734 43716
rect 34054 43664 34060 43716
rect 34112 43704 34118 43716
rect 35069 43707 35127 43713
rect 35069 43704 35081 43707
rect 34112 43676 35081 43704
rect 34112 43664 34118 43676
rect 35069 43673 35081 43676
rect 35115 43673 35127 43707
rect 35069 43667 35127 43673
rect 1765 43639 1823 43645
rect 1765 43605 1777 43639
rect 1811 43636 1823 43639
rect 33962 43636 33968 43648
rect 1811 43608 33968 43636
rect 1811 43605 1823 43608
rect 1765 43599 1823 43605
rect 33962 43596 33968 43608
rect 34020 43596 34026 43648
rect 35084 43636 35112 43667
rect 35158 43664 35164 43716
rect 35216 43704 35222 43716
rect 35866 43704 35894 43744
rect 50798 43732 50804 43784
rect 50856 43772 50862 43784
rect 57885 43775 57943 43781
rect 57885 43772 57897 43775
rect 50856 43744 57897 43772
rect 50856 43732 50862 43744
rect 57885 43741 57897 43744
rect 57931 43741 57943 43775
rect 57885 43735 57943 43741
rect 36170 43704 36176 43716
rect 35216 43676 35261 43704
rect 35866 43676 36176 43704
rect 35216 43664 35222 43676
rect 36170 43664 36176 43676
rect 36228 43664 36234 43716
rect 58158 43704 58164 43716
rect 58119 43676 58164 43704
rect 58158 43664 58164 43676
rect 58216 43664 58222 43716
rect 36446 43636 36452 43648
rect 35084 43608 36452 43636
rect 36446 43596 36452 43608
rect 36504 43596 36510 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 6730 43392 6736 43444
rect 6788 43432 6794 43444
rect 22002 43432 22008 43444
rect 6788 43404 22008 43432
rect 6788 43392 6794 43404
rect 22002 43392 22008 43404
rect 22060 43392 22066 43444
rect 37182 43392 37188 43444
rect 37240 43432 37246 43444
rect 54294 43432 54300 43444
rect 37240 43404 54300 43432
rect 37240 43392 37246 43404
rect 54294 43392 54300 43404
rect 54352 43392 54358 43444
rect 34238 43364 34244 43376
rect 34199 43336 34244 43364
rect 34238 43324 34244 43336
rect 34296 43324 34302 43376
rect 1578 43296 1584 43308
rect 1539 43268 1584 43296
rect 1578 43256 1584 43268
rect 1636 43256 1642 43308
rect 33962 43296 33968 43308
rect 33923 43268 33968 43296
rect 33962 43256 33968 43268
rect 34020 43256 34026 43308
rect 34054 43256 34060 43308
rect 34112 43296 34118 43308
rect 34149 43299 34207 43305
rect 34149 43296 34161 43299
rect 34112 43268 34161 43296
rect 34112 43256 34118 43268
rect 34149 43265 34161 43268
rect 34195 43265 34207 43299
rect 34149 43259 34207 43265
rect 34385 43299 34443 43305
rect 34385 43265 34397 43299
rect 34431 43296 34443 43299
rect 37366 43296 37372 43308
rect 34431 43268 37372 43296
rect 34431 43265 34443 43268
rect 34385 43259 34443 43265
rect 37366 43256 37372 43268
rect 37424 43256 37430 43308
rect 1762 43092 1768 43104
rect 1723 43064 1768 43092
rect 1762 43052 1768 43064
rect 1820 43052 1826 43104
rect 34514 43092 34520 43104
rect 34475 43064 34520 43092
rect 34514 43052 34520 43064
rect 34572 43052 34578 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 36170 42820 36176 42832
rect 33428 42792 36176 42820
rect 24302 42712 24308 42764
rect 24360 42752 24366 42764
rect 33428 42752 33456 42792
rect 36170 42780 36176 42792
rect 36228 42780 36234 42832
rect 37461 42823 37519 42829
rect 37461 42789 37473 42823
rect 37507 42789 37519 42823
rect 37461 42783 37519 42789
rect 24360 42724 33456 42752
rect 24360 42712 24366 42724
rect 1762 42644 1768 42696
rect 1820 42684 1826 42696
rect 33336 42693 33364 42724
rect 33502 42712 33508 42764
rect 33560 42712 33566 42764
rect 37476 42752 37504 42783
rect 33704 42724 37504 42752
rect 33321 42687 33379 42693
rect 1820 42656 33088 42684
rect 1820 42644 1826 42656
rect 32950 42548 32956 42560
rect 32911 42520 32956 42548
rect 32950 42508 32956 42520
rect 33008 42508 33014 42560
rect 33060 42548 33088 42656
rect 33321 42653 33333 42687
rect 33367 42653 33379 42687
rect 33321 42647 33379 42653
rect 33413 42687 33471 42693
rect 33413 42653 33425 42687
rect 33459 42684 33471 42687
rect 33520 42684 33548 42712
rect 33704 42693 33732 42724
rect 33459 42656 33548 42684
rect 33689 42687 33747 42693
rect 33459 42653 33471 42656
rect 33413 42647 33471 42653
rect 33689 42653 33701 42687
rect 33735 42653 33747 42687
rect 33962 42684 33968 42696
rect 33923 42656 33968 42684
rect 33689 42647 33747 42653
rect 33962 42644 33968 42656
rect 34020 42644 34026 42696
rect 34149 42687 34207 42693
rect 34149 42653 34161 42687
rect 34195 42653 34207 42687
rect 36906 42684 36912 42696
rect 36867 42656 36912 42684
rect 34149 42647 34207 42653
rect 34164 42548 34192 42647
rect 36906 42644 36912 42656
rect 36964 42644 36970 42696
rect 37182 42684 37188 42696
rect 37143 42656 37188 42684
rect 37182 42644 37188 42656
rect 37240 42644 37246 42696
rect 37277 42687 37335 42693
rect 37277 42653 37289 42687
rect 37323 42684 37335 42687
rect 37366 42684 37372 42696
rect 37323 42656 37372 42684
rect 37323 42653 37335 42656
rect 37277 42647 37335 42653
rect 37366 42644 37372 42656
rect 37424 42644 37430 42696
rect 37090 42616 37096 42628
rect 37051 42588 37096 42616
rect 37090 42576 37096 42588
rect 37148 42576 37154 42628
rect 57054 42616 57060 42628
rect 57015 42588 57060 42616
rect 57054 42576 57060 42588
rect 57112 42576 57118 42628
rect 57974 42616 57980 42628
rect 57935 42588 57980 42616
rect 57974 42576 57980 42588
rect 58032 42576 58038 42628
rect 58345 42619 58403 42625
rect 58345 42585 58357 42619
rect 58391 42616 58403 42619
rect 58618 42616 58624 42628
rect 58391 42588 58624 42616
rect 58391 42585 58403 42588
rect 58345 42579 58403 42585
rect 58618 42576 58624 42588
rect 58676 42576 58682 42628
rect 57146 42548 57152 42560
rect 33060 42520 34192 42548
rect 57107 42520 57152 42548
rect 57146 42508 57152 42520
rect 57204 42508 57210 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 23474 42304 23480 42356
rect 23532 42344 23538 42356
rect 37090 42344 37096 42356
rect 23532 42316 37096 42344
rect 23532 42304 23538 42316
rect 37090 42304 37096 42316
rect 37148 42304 37154 42356
rect 1670 42208 1676 42220
rect 1631 42180 1676 42208
rect 1670 42168 1676 42180
rect 1728 42168 1734 42220
rect 5442 42100 5448 42152
rect 5500 42140 5506 42152
rect 20898 42140 20904 42152
rect 5500 42112 20904 42140
rect 5500 42100 5506 42112
rect 20898 42100 20904 42112
rect 20956 42100 20962 42152
rect 1857 42075 1915 42081
rect 1857 42041 1869 42075
rect 1903 42072 1915 42075
rect 5534 42072 5540 42084
rect 1903 42044 5540 42072
rect 1903 42041 1915 42044
rect 1857 42035 1915 42041
rect 5534 42032 5540 42044
rect 5592 42032 5598 42084
rect 42886 42072 42892 42084
rect 6886 42044 42892 42072
rect 5626 41964 5632 42016
rect 5684 42004 5690 42016
rect 6886 42004 6914 42044
rect 42886 42032 42892 42044
rect 42944 42032 42950 42084
rect 5684 41976 6914 42004
rect 5684 41964 5690 41976
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 23750 41692 23756 41744
rect 23808 41732 23814 41744
rect 23808 41704 25636 41732
rect 23808 41692 23814 41704
rect 24118 41624 24124 41676
rect 24176 41664 24182 41676
rect 25133 41667 25191 41673
rect 25133 41664 25145 41667
rect 24176 41636 25145 41664
rect 24176 41624 24182 41636
rect 25133 41633 25145 41636
rect 25179 41633 25191 41667
rect 25133 41627 25191 41633
rect 24026 41556 24032 41608
rect 24084 41596 24090 41608
rect 25608 41605 25636 41704
rect 25225 41599 25283 41605
rect 25225 41596 25237 41599
rect 24084 41568 25237 41596
rect 24084 41556 24090 41568
rect 25225 41565 25237 41568
rect 25271 41565 25283 41599
rect 25225 41559 25283 41565
rect 25593 41599 25651 41605
rect 25593 41565 25605 41599
rect 25639 41565 25651 41599
rect 25593 41559 25651 41565
rect 25685 41599 25743 41605
rect 25685 41565 25697 41599
rect 25731 41565 25743 41599
rect 25685 41559 25743 41565
rect 1670 41528 1676 41540
rect 1631 41500 1676 41528
rect 1670 41488 1676 41500
rect 1728 41488 1734 41540
rect 24578 41528 24584 41540
rect 24539 41500 24584 41528
rect 24578 41488 24584 41500
rect 24636 41488 24642 41540
rect 1765 41463 1823 41469
rect 1765 41429 1777 41463
rect 1811 41460 1823 41463
rect 1854 41460 1860 41472
rect 1811 41432 1860 41460
rect 1811 41429 1823 41432
rect 1765 41423 1823 41429
rect 1854 41420 1860 41432
rect 1912 41420 1918 41472
rect 20806 41420 20812 41472
rect 20864 41460 20870 41472
rect 25700 41460 25728 41559
rect 51718 41556 51724 41608
rect 51776 41596 51782 41608
rect 56965 41599 57023 41605
rect 56965 41596 56977 41599
rect 51776 41568 56977 41596
rect 51776 41556 51782 41568
rect 56965 41565 56977 41568
rect 57011 41565 57023 41599
rect 56965 41559 57023 41565
rect 57238 41528 57244 41540
rect 57199 41500 57244 41528
rect 57238 41488 57244 41500
rect 57296 41488 57302 41540
rect 57882 41488 57888 41540
rect 57940 41528 57946 41540
rect 57977 41531 58035 41537
rect 57977 41528 57989 41531
rect 57940 41500 57989 41528
rect 57940 41488 57946 41500
rect 57977 41497 57989 41500
rect 58023 41497 58035 41531
rect 57977 41491 58035 41497
rect 20864 41432 25728 41460
rect 20864 41420 20870 41432
rect 38562 41420 38568 41472
rect 38620 41460 38626 41472
rect 58069 41463 58127 41469
rect 58069 41460 58081 41463
rect 38620 41432 58081 41460
rect 38620 41420 38626 41432
rect 58069 41429 58081 41432
rect 58115 41429 58127 41463
rect 58069 41423 58127 41429
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1670 41120 1676 41132
rect 1631 41092 1676 41120
rect 1670 41080 1676 41092
rect 1728 41080 1734 41132
rect 5534 40944 5540 40996
rect 5592 40984 5598 40996
rect 22370 40984 22376 40996
rect 5592 40956 22376 40984
rect 5592 40944 5598 40956
rect 22370 40944 22376 40956
rect 22428 40944 22434 40996
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 20530 40916 20536 40928
rect 1811 40888 20536 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 20530 40876 20536 40888
rect 20588 40876 20594 40928
rect 36814 40876 36820 40928
rect 36872 40916 36878 40928
rect 48958 40916 48964 40928
rect 36872 40888 48964 40916
rect 36872 40876 36878 40888
rect 48958 40876 48964 40888
rect 49016 40876 49022 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 20162 40672 20168 40724
rect 20220 40712 20226 40724
rect 41046 40712 41052 40724
rect 20220 40684 41052 40712
rect 20220 40672 20226 40684
rect 41046 40672 41052 40684
rect 41104 40672 41110 40724
rect 56962 40508 56968 40520
rect 56923 40480 56968 40508
rect 56962 40468 56968 40480
rect 57020 40468 57026 40520
rect 57790 40468 57796 40520
rect 57848 40508 57854 40520
rect 57885 40511 57943 40517
rect 57885 40508 57897 40511
rect 57848 40480 57897 40508
rect 57848 40468 57854 40480
rect 57885 40477 57897 40480
rect 57931 40477 57943 40511
rect 57885 40471 57943 40477
rect 1670 40440 1676 40452
rect 1631 40412 1676 40440
rect 1670 40400 1676 40412
rect 1728 40400 1734 40452
rect 44082 40400 44088 40452
rect 44140 40440 44146 40452
rect 57241 40443 57299 40449
rect 57241 40440 57253 40443
rect 44140 40412 57253 40440
rect 44140 40400 44146 40412
rect 57241 40409 57253 40412
rect 57287 40409 57299 40443
rect 58161 40443 58219 40449
rect 58161 40440 58173 40443
rect 57241 40403 57299 40409
rect 57900 40412 58173 40440
rect 57900 40384 57928 40412
rect 58161 40409 58173 40412
rect 58207 40409 58219 40443
rect 58161 40403 58219 40409
rect 1765 40375 1823 40381
rect 1765 40341 1777 40375
rect 1811 40372 1823 40375
rect 11054 40372 11060 40384
rect 1811 40344 11060 40372
rect 1811 40341 1823 40344
rect 1765 40335 1823 40341
rect 11054 40332 11060 40344
rect 11112 40332 11118 40384
rect 57882 40332 57888 40384
rect 57940 40332 57946 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 15838 40060 15844 40112
rect 15896 40100 15902 40112
rect 19334 40100 19340 40112
rect 15896 40072 19340 40100
rect 15896 40060 15902 40072
rect 19334 40060 19340 40072
rect 19392 40060 19398 40112
rect 26602 40060 26608 40112
rect 26660 40100 26666 40112
rect 30282 40100 30288 40112
rect 26660 40072 30288 40100
rect 26660 40060 26666 40072
rect 30282 40060 30288 40072
rect 30340 40060 30346 40112
rect 33318 40060 33324 40112
rect 33376 40100 33382 40112
rect 38562 40100 38568 40112
rect 33376 40072 38568 40100
rect 33376 40060 33382 40072
rect 38562 40060 38568 40072
rect 38620 40060 38626 40112
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2869 39559 2927 39565
rect 2869 39525 2881 39559
rect 2915 39556 2927 39559
rect 15838 39556 15844 39568
rect 2915 39528 15844 39556
rect 2915 39525 2927 39528
rect 2869 39519 2927 39525
rect 15838 39516 15844 39528
rect 15896 39516 15902 39568
rect 1857 39491 1915 39497
rect 1857 39457 1869 39491
rect 1903 39488 1915 39491
rect 1903 39460 2636 39488
rect 1903 39457 1915 39460
rect 1857 39451 1915 39457
rect 2314 39420 2320 39432
rect 2275 39392 2320 39420
rect 2314 39380 2320 39392
rect 2372 39380 2378 39432
rect 2608 39429 2636 39460
rect 2746 39460 21036 39488
rect 2746 39429 2774 39460
rect 2593 39423 2651 39429
rect 2593 39389 2605 39423
rect 2639 39389 2651 39423
rect 2593 39383 2651 39389
rect 2731 39423 2789 39429
rect 2731 39389 2743 39423
rect 2777 39389 2789 39423
rect 20622 39420 20628 39432
rect 20583 39392 20628 39420
rect 2731 39383 2789 39389
rect 20622 39380 20628 39392
rect 20680 39380 20686 39432
rect 21008 39429 21036 39460
rect 20901 39423 20959 39429
rect 20901 39420 20913 39423
rect 20732 39392 20913 39420
rect 1670 39352 1676 39364
rect 1631 39324 1676 39352
rect 1670 39312 1676 39324
rect 1728 39312 1734 39364
rect 2501 39355 2559 39361
rect 2501 39321 2513 39355
rect 2547 39321 2559 39355
rect 2501 39315 2559 39321
rect 2516 39284 2544 39315
rect 20530 39312 20536 39364
rect 20588 39352 20594 39364
rect 20732 39352 20760 39392
rect 20901 39389 20913 39392
rect 20947 39389 20959 39423
rect 20901 39383 20959 39389
rect 20993 39423 21051 39429
rect 20993 39389 21005 39423
rect 21039 39420 21051 39423
rect 22094 39420 22100 39432
rect 21039 39392 22100 39420
rect 21039 39389 21051 39392
rect 20993 39383 21051 39389
rect 22094 39380 22100 39392
rect 22152 39380 22158 39432
rect 20588 39324 20760 39352
rect 20588 39312 20594 39324
rect 20806 39312 20812 39364
rect 20864 39352 20870 39364
rect 57054 39352 57060 39364
rect 20864 39324 20909 39352
rect 57015 39324 57060 39352
rect 20864 39312 20870 39324
rect 57054 39312 57060 39324
rect 57112 39312 57118 39364
rect 57974 39352 57980 39364
rect 57935 39324 57980 39352
rect 57974 39312 57980 39324
rect 58032 39312 58038 39364
rect 2590 39284 2596 39296
rect 2516 39256 2596 39284
rect 2590 39244 2596 39256
rect 2648 39244 2654 39296
rect 21177 39287 21235 39293
rect 21177 39253 21189 39287
rect 21223 39284 21235 39287
rect 21358 39284 21364 39296
rect 21223 39256 21364 39284
rect 21223 39253 21235 39256
rect 21177 39247 21235 39253
rect 21358 39244 21364 39256
rect 21416 39244 21422 39296
rect 35526 39244 35532 39296
rect 35584 39284 35590 39296
rect 57149 39287 57207 39293
rect 57149 39284 57161 39287
rect 35584 39256 57161 39284
rect 35584 39244 35590 39256
rect 57149 39253 57161 39256
rect 57195 39253 57207 39287
rect 58066 39284 58072 39296
rect 58027 39256 58072 39284
rect 57149 39247 57207 39253
rect 58066 39244 58072 39256
rect 58124 39244 58130 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 34054 39040 34060 39092
rect 34112 39080 34118 39092
rect 34112 39052 35894 39080
rect 34112 39040 34118 39052
rect 9306 38972 9312 39024
rect 9364 39012 9370 39024
rect 34333 39015 34391 39021
rect 34333 39012 34345 39015
rect 9364 38984 34345 39012
rect 9364 38972 9370 38984
rect 34333 38981 34345 38984
rect 34379 38981 34391 39015
rect 34333 38975 34391 38981
rect 1670 38944 1676 38956
rect 1631 38916 1676 38944
rect 1670 38904 1676 38916
rect 1728 38904 1734 38956
rect 34054 38944 34060 38956
rect 34015 38916 34060 38944
rect 34054 38904 34060 38916
rect 34112 38904 34118 38956
rect 34241 38947 34299 38953
rect 34241 38944 34253 38947
rect 34164 38916 34253 38944
rect 26050 38836 26056 38888
rect 26108 38876 26114 38888
rect 34164 38876 34192 38916
rect 34241 38913 34253 38916
rect 34287 38913 34299 38947
rect 34241 38907 34299 38913
rect 34422 38904 34428 38956
rect 34480 38953 34486 38956
rect 34480 38944 34488 38953
rect 35866 38944 35894 39052
rect 47670 39040 47676 39092
rect 47728 39080 47734 39092
rect 58066 39080 58072 39092
rect 47728 39052 58072 39080
rect 47728 39040 47734 39052
rect 58066 39040 58072 39052
rect 58124 39040 58130 39092
rect 45830 38944 45836 38956
rect 34480 38916 34525 38944
rect 35866 38916 45836 38944
rect 34480 38907 34488 38916
rect 34480 38904 34486 38907
rect 45830 38904 45836 38916
rect 45888 38904 45894 38956
rect 26108 38848 34192 38876
rect 26108 38836 26114 38848
rect 1857 38811 1915 38817
rect 1857 38777 1869 38811
rect 1903 38808 1915 38811
rect 4798 38808 4804 38820
rect 1903 38780 4804 38808
rect 1903 38777 1915 38780
rect 1857 38771 1915 38777
rect 4798 38768 4804 38780
rect 4856 38768 4862 38820
rect 34164 38740 34192 38848
rect 34606 38808 34612 38820
rect 34567 38780 34612 38808
rect 34606 38768 34612 38780
rect 34664 38768 34670 38820
rect 38562 38740 38568 38752
rect 34164 38712 38568 38740
rect 38562 38700 38568 38712
rect 38620 38700 38626 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 23474 38400 23480 38412
rect 23032 38372 23480 38400
rect 22738 38332 22744 38344
rect 22699 38304 22744 38332
rect 22738 38292 22744 38304
rect 22796 38292 22802 38344
rect 22922 38341 22928 38344
rect 22889 38335 22928 38341
rect 22889 38301 22901 38335
rect 22889 38295 22928 38301
rect 22922 38292 22928 38295
rect 22980 38292 22986 38344
rect 23032 38276 23060 38372
rect 23474 38360 23480 38372
rect 23532 38360 23538 38412
rect 23198 38292 23204 38344
rect 23256 38341 23262 38344
rect 23256 38332 23264 38341
rect 23256 38304 23301 38332
rect 23256 38295 23264 38304
rect 23256 38292 23262 38295
rect 49050 38292 49056 38344
rect 49108 38332 49114 38344
rect 57885 38335 57943 38341
rect 57885 38332 57897 38335
rect 49108 38304 57897 38332
rect 49108 38292 49114 38304
rect 57885 38301 57897 38304
rect 57931 38301 57943 38335
rect 57885 38295 57943 38301
rect 1670 38264 1676 38276
rect 1631 38236 1676 38264
rect 1670 38224 1676 38236
rect 1728 38224 1734 38276
rect 11054 38224 11060 38276
rect 11112 38264 11118 38276
rect 23014 38264 23020 38276
rect 11112 38236 22094 38264
rect 22975 38236 23020 38264
rect 11112 38224 11118 38236
rect 1765 38199 1823 38205
rect 1765 38165 1777 38199
rect 1811 38196 1823 38199
rect 19426 38196 19432 38208
rect 1811 38168 19432 38196
rect 1811 38165 1823 38168
rect 1765 38159 1823 38165
rect 19426 38156 19432 38168
rect 19484 38156 19490 38208
rect 22066 38196 22094 38236
rect 23014 38224 23020 38236
rect 23072 38224 23078 38276
rect 23109 38267 23167 38273
rect 23109 38233 23121 38267
rect 23155 38233 23167 38267
rect 58158 38264 58164 38276
rect 58119 38236 58164 38264
rect 23109 38227 23167 38233
rect 23124 38196 23152 38227
rect 58158 38224 58164 38236
rect 58216 38224 58222 38276
rect 22066 38168 23152 38196
rect 23385 38199 23443 38205
rect 23385 38165 23397 38199
rect 23431 38196 23443 38199
rect 23658 38196 23664 38208
rect 23431 38168 23664 38196
rect 23431 38165 23443 38168
rect 23385 38159 23443 38165
rect 23658 38156 23664 38168
rect 23716 38156 23722 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 20898 37992 20904 38004
rect 19352 37964 20760 37992
rect 20859 37964 20904 37992
rect 1670 37856 1676 37868
rect 1631 37828 1676 37856
rect 1670 37816 1676 37828
rect 1728 37816 1734 37868
rect 4798 37856 4804 37868
rect 4759 37828 4804 37856
rect 4798 37816 4804 37828
rect 4856 37816 4862 37868
rect 4982 37816 4988 37868
rect 5040 37856 5046 37868
rect 19242 37856 19248 37868
rect 5040 37828 12434 37856
rect 19203 37828 19248 37856
rect 5040 37816 5046 37828
rect 1857 37723 1915 37729
rect 1857 37689 1869 37723
rect 1903 37720 1915 37723
rect 4062 37720 4068 37732
rect 1903 37692 4068 37720
rect 1903 37689 1915 37692
rect 1857 37683 1915 37689
rect 4062 37680 4068 37692
rect 4120 37680 4126 37732
rect 12406 37720 12434 37828
rect 19242 37816 19248 37828
rect 19300 37816 19306 37868
rect 19352 37865 19380 37964
rect 19426 37884 19432 37936
rect 19484 37924 19490 37936
rect 19613 37927 19671 37933
rect 19613 37924 19625 37927
rect 19484 37896 19625 37924
rect 19484 37884 19490 37896
rect 19613 37893 19625 37896
rect 19659 37893 19671 37927
rect 20732 37924 20760 37964
rect 20898 37952 20904 37964
rect 20956 37952 20962 38004
rect 22922 37952 22928 38004
rect 22980 37992 22986 38004
rect 38010 37992 38016 38004
rect 22980 37964 38016 37992
rect 22980 37952 22986 37964
rect 38010 37952 38016 37964
rect 38068 37952 38074 38004
rect 51994 37952 52000 38004
rect 52052 37992 52058 38004
rect 58250 37992 58256 38004
rect 52052 37964 58256 37992
rect 52052 37952 52058 37964
rect 58250 37952 58256 37964
rect 58308 37952 58314 38004
rect 20732 37896 35894 37924
rect 19613 37887 19671 37893
rect 19338 37859 19396 37865
rect 19338 37825 19350 37859
rect 19384 37825 19396 37859
rect 19518 37856 19524 37868
rect 19479 37828 19524 37856
rect 19338 37819 19396 37825
rect 19518 37816 19524 37828
rect 19576 37816 19582 37868
rect 19702 37816 19708 37868
rect 19760 37865 19766 37868
rect 19760 37859 19787 37865
rect 19775 37825 19787 37859
rect 19760 37819 19787 37825
rect 20717 37859 20775 37865
rect 20717 37825 20729 37859
rect 20763 37825 20775 37859
rect 20717 37819 20775 37825
rect 20993 37859 21051 37865
rect 20993 37825 21005 37859
rect 21039 37856 21051 37859
rect 24302 37856 24308 37868
rect 21039 37828 24308 37856
rect 21039 37825 21051 37828
rect 20993 37819 21051 37825
rect 19760 37816 19766 37819
rect 20257 37791 20315 37797
rect 20257 37757 20269 37791
rect 20303 37788 20315 37791
rect 20732 37788 20760 37819
rect 24302 37816 24308 37828
rect 24360 37816 24366 37868
rect 35866 37788 35894 37896
rect 58066 37856 58072 37868
rect 58027 37828 58072 37856
rect 58066 37816 58072 37828
rect 58124 37816 58130 37868
rect 47946 37788 47952 37800
rect 20303 37760 31754 37788
rect 35866 37760 47952 37788
rect 20303 37757 20315 37760
rect 20257 37751 20315 37757
rect 19702 37720 19708 37732
rect 12406 37692 19708 37720
rect 19702 37680 19708 37692
rect 19760 37720 19766 37732
rect 22554 37720 22560 37732
rect 19760 37692 22560 37720
rect 19760 37680 19766 37692
rect 22554 37680 22560 37692
rect 22612 37680 22618 37732
rect 31726 37720 31754 37760
rect 47946 37748 47952 37760
rect 48004 37748 48010 37800
rect 54018 37720 54024 37732
rect 31726 37692 54024 37720
rect 54018 37680 54024 37692
rect 54076 37680 54082 37732
rect 5169 37655 5227 37661
rect 5169 37621 5181 37655
rect 5215 37652 5227 37655
rect 6730 37652 6736 37664
rect 5215 37624 6736 37652
rect 5215 37621 5227 37624
rect 5169 37615 5227 37621
rect 6730 37612 6736 37624
rect 6788 37612 6794 37664
rect 19889 37655 19947 37661
rect 19889 37621 19901 37655
rect 19935 37652 19947 37655
rect 20070 37652 20076 37664
rect 19935 37624 20076 37652
rect 19935 37621 19947 37624
rect 19889 37615 19947 37621
rect 20070 37612 20076 37624
rect 20128 37612 20134 37664
rect 20530 37652 20536 37664
rect 20491 37624 20536 37652
rect 20530 37612 20536 37624
rect 20588 37612 20594 37664
rect 58250 37652 58256 37664
rect 58211 37624 58256 37652
rect 58250 37612 58256 37624
rect 58308 37612 58314 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 20349 37451 20407 37457
rect 20349 37417 20361 37451
rect 20395 37448 20407 37451
rect 22094 37448 22100 37460
rect 20395 37420 22100 37448
rect 20395 37417 20407 37420
rect 20349 37411 20407 37417
rect 22094 37408 22100 37420
rect 22152 37408 22158 37460
rect 20533 37383 20591 37389
rect 20533 37380 20545 37383
rect 15120 37352 20545 37380
rect 2038 37244 2044 37256
rect 1999 37216 2044 37244
rect 2038 37204 2044 37216
rect 2096 37204 2102 37256
rect 2409 37247 2467 37253
rect 2409 37213 2421 37247
rect 2455 37244 2467 37247
rect 6178 37244 6184 37256
rect 2455 37216 6184 37244
rect 2455 37213 2467 37216
rect 2409 37207 2467 37213
rect 6178 37204 6184 37216
rect 6236 37204 6242 37256
rect 2222 37176 2228 37188
rect 2135 37148 2228 37176
rect 2222 37136 2228 37148
rect 2280 37136 2286 37188
rect 2314 37136 2320 37188
rect 2372 37176 2378 37188
rect 7558 37176 7564 37188
rect 2372 37148 2417 37176
rect 2516 37148 7564 37176
rect 2372 37136 2378 37148
rect 2240 37108 2268 37136
rect 2516 37108 2544 37148
rect 7558 37136 7564 37148
rect 7616 37136 7622 37188
rect 2240 37080 2544 37108
rect 2593 37111 2651 37117
rect 2593 37077 2605 37111
rect 2639 37108 2651 37111
rect 15120 37108 15148 37352
rect 20533 37349 20545 37352
rect 20579 37349 20591 37383
rect 20533 37343 20591 37349
rect 20073 37315 20131 37321
rect 20073 37281 20085 37315
rect 20119 37312 20131 37315
rect 21082 37312 21088 37324
rect 20119 37284 21088 37312
rect 20119 37281 20131 37284
rect 20073 37275 20131 37281
rect 21082 37272 21088 37284
rect 21140 37272 21146 37324
rect 18414 37244 18420 37256
rect 18375 37216 18420 37244
rect 18414 37204 18420 37216
rect 18472 37204 18478 37256
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 20220 37216 20453 37244
rect 20220 37204 20226 37216
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 20625 37247 20683 37253
rect 20625 37213 20637 37247
rect 20671 37213 20683 37247
rect 20625 37207 20683 37213
rect 20809 37247 20867 37253
rect 20809 37213 20821 37247
rect 20855 37213 20867 37247
rect 20809 37207 20867 37213
rect 18690 37176 18696 37188
rect 18651 37148 18696 37176
rect 18690 37136 18696 37148
rect 18748 37176 18754 37188
rect 19242 37176 19248 37188
rect 18748 37148 19248 37176
rect 18748 37136 18754 37148
rect 19242 37136 19248 37148
rect 19300 37136 19306 37188
rect 20254 37136 20260 37188
rect 20312 37176 20318 37188
rect 20640 37176 20668 37207
rect 20312 37148 20668 37176
rect 20312 37136 20318 37148
rect 2639 37080 15148 37108
rect 2639 37077 2651 37080
rect 2593 37071 2651 37077
rect 16390 37068 16396 37120
rect 16448 37108 16454 37120
rect 20824 37108 20852 37207
rect 48958 37204 48964 37256
rect 49016 37244 49022 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 49016 37216 57897 37244
rect 49016 37204 49022 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 58158 37176 58164 37188
rect 58119 37148 58164 37176
rect 58158 37136 58164 37148
rect 58216 37136 58222 37188
rect 21634 37108 21640 37120
rect 16448 37080 21640 37108
rect 16448 37068 16454 37080
rect 21634 37068 21640 37080
rect 21692 37068 21698 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 53745 36907 53803 36913
rect 53745 36904 53757 36907
rect 6932 36876 53757 36904
rect 2130 36796 2136 36848
rect 2188 36836 2194 36848
rect 2317 36839 2375 36845
rect 2317 36836 2329 36839
rect 2188 36808 2329 36836
rect 2188 36796 2194 36808
rect 2317 36805 2329 36808
rect 2363 36805 2375 36839
rect 2317 36799 2375 36805
rect 2590 36796 2596 36848
rect 2648 36836 2654 36848
rect 6638 36836 6644 36848
rect 2648 36808 6500 36836
rect 6599 36808 6644 36836
rect 2648 36796 2654 36808
rect 1946 36728 1952 36780
rect 2004 36768 2010 36780
rect 2041 36771 2099 36777
rect 2041 36768 2053 36771
rect 2004 36740 2053 36768
rect 2004 36728 2010 36740
rect 2041 36737 2053 36740
rect 2087 36737 2099 36771
rect 2222 36768 2228 36780
rect 2183 36740 2228 36768
rect 2041 36731 2099 36737
rect 2222 36728 2228 36740
rect 2280 36728 2286 36780
rect 2409 36771 2467 36777
rect 2409 36737 2421 36771
rect 2455 36768 2467 36771
rect 2682 36768 2688 36780
rect 2455 36740 2688 36768
rect 2455 36737 2467 36740
rect 2409 36731 2467 36737
rect 2682 36728 2688 36740
rect 2740 36728 2746 36780
rect 3050 36768 3056 36780
rect 3011 36740 3056 36768
rect 3050 36728 3056 36740
rect 3108 36728 3114 36780
rect 6472 36768 6500 36808
rect 6638 36796 6644 36808
rect 6696 36796 6702 36848
rect 6932 36777 6960 36876
rect 53745 36873 53757 36876
rect 53791 36873 53803 36907
rect 53745 36867 53803 36873
rect 7006 36796 7012 36848
rect 7064 36836 7070 36848
rect 18690 36836 18696 36848
rect 7064 36808 18696 36836
rect 7064 36796 7070 36808
rect 18690 36796 18696 36808
rect 18748 36796 18754 36848
rect 19058 36796 19064 36848
rect 19116 36836 19122 36848
rect 33962 36836 33968 36848
rect 19116 36808 19161 36836
rect 19306 36808 22094 36836
rect 19116 36796 19122 36808
rect 19306 36780 19334 36808
rect 6917 36771 6975 36777
rect 6472 36740 6868 36768
rect 6730 36700 6736 36712
rect 6691 36672 6736 36700
rect 6730 36660 6736 36672
rect 6788 36660 6794 36712
rect 6840 36700 6868 36740
rect 6917 36737 6929 36771
rect 6963 36737 6975 36771
rect 17954 36768 17960 36780
rect 17915 36740 17960 36768
rect 6917 36731 6975 36737
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 18785 36771 18843 36777
rect 18785 36766 18797 36771
rect 18708 36738 18797 36766
rect 7834 36700 7840 36712
rect 6840 36672 7840 36700
rect 7834 36660 7840 36672
rect 7892 36660 7898 36712
rect 18046 36700 18052 36712
rect 18007 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 18138 36660 18144 36712
rect 18196 36700 18202 36712
rect 18708 36700 18736 36738
rect 18785 36737 18797 36738
rect 18831 36737 18843 36771
rect 18785 36731 18843 36737
rect 18874 36728 18880 36780
rect 18932 36768 18938 36780
rect 19242 36777 19248 36780
rect 18969 36771 19027 36777
rect 18969 36768 18981 36771
rect 18932 36740 18981 36768
rect 18932 36728 18938 36740
rect 18969 36737 18981 36740
rect 19015 36737 19027 36771
rect 19199 36771 19248 36777
rect 19199 36768 19211 36771
rect 19155 36740 19211 36768
rect 18969 36731 19027 36737
rect 19199 36737 19211 36740
rect 19245 36737 19248 36771
rect 19199 36731 19248 36737
rect 19242 36728 19248 36731
rect 19300 36740 19334 36780
rect 19981 36771 20039 36777
rect 19300 36728 19306 36740
rect 19981 36737 19993 36771
rect 20027 36737 20039 36771
rect 19981 36731 20039 36737
rect 19996 36700 20024 36731
rect 20070 36728 20076 36780
rect 20128 36768 20134 36780
rect 20257 36771 20315 36777
rect 20257 36768 20269 36771
rect 20128 36740 20269 36768
rect 20128 36728 20134 36740
rect 20257 36737 20269 36740
rect 20303 36737 20315 36771
rect 20257 36731 20315 36737
rect 20438 36700 20444 36712
rect 18196 36672 18736 36700
rect 18846 36672 20024 36700
rect 20399 36672 20444 36700
rect 18196 36660 18202 36672
rect 2593 36635 2651 36641
rect 2593 36601 2605 36635
rect 2639 36632 2651 36635
rect 18325 36635 18383 36641
rect 2639 36604 6684 36632
rect 2639 36601 2651 36604
rect 2593 36595 2651 36601
rect 3234 36564 3240 36576
rect 3195 36536 3240 36564
rect 3234 36524 3240 36536
rect 3292 36524 3298 36576
rect 6656 36573 6684 36604
rect 18325 36601 18337 36635
rect 18371 36632 18383 36635
rect 18846 36632 18874 36672
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 18371 36604 18874 36632
rect 18371 36601 18383 36604
rect 18325 36595 18383 36601
rect 19150 36592 19156 36644
rect 19208 36632 19214 36644
rect 19337 36635 19395 36641
rect 19337 36632 19349 36635
rect 19208 36604 19349 36632
rect 19208 36592 19214 36604
rect 19337 36601 19349 36604
rect 19383 36601 19395 36635
rect 19337 36595 19395 36601
rect 20073 36635 20131 36641
rect 20073 36601 20085 36635
rect 20119 36632 20131 36635
rect 20530 36632 20536 36644
rect 20119 36604 20536 36632
rect 20119 36601 20131 36604
rect 20073 36595 20131 36601
rect 20530 36592 20536 36604
rect 20588 36592 20594 36644
rect 22066 36632 22094 36808
rect 26988 36808 33968 36836
rect 23569 36771 23627 36777
rect 23569 36737 23581 36771
rect 23615 36768 23627 36771
rect 23750 36768 23756 36780
rect 23615 36740 23756 36768
rect 23615 36737 23627 36740
rect 23569 36731 23627 36737
rect 23750 36728 23756 36740
rect 23808 36768 23814 36780
rect 24302 36768 24308 36780
rect 23808 36740 24308 36768
rect 23808 36728 23814 36740
rect 24302 36728 24308 36740
rect 24360 36728 24366 36780
rect 22830 36660 22836 36712
rect 22888 36700 22894 36712
rect 24213 36703 24271 36709
rect 24213 36700 24225 36703
rect 22888 36672 24225 36700
rect 22888 36660 22894 36672
rect 24213 36669 24225 36672
rect 24259 36700 24271 36703
rect 26988 36700 27016 36808
rect 33962 36796 33968 36808
rect 34020 36796 34026 36848
rect 53650 36728 53656 36780
rect 53708 36768 53714 36780
rect 54297 36771 54355 36777
rect 54297 36768 54309 36771
rect 53708 36740 54309 36768
rect 53708 36728 53714 36740
rect 54297 36737 54309 36740
rect 54343 36737 54355 36771
rect 54297 36731 54355 36737
rect 54665 36771 54723 36777
rect 54665 36737 54677 36771
rect 54711 36768 54723 36771
rect 56594 36768 56600 36780
rect 54711 36740 56600 36768
rect 54711 36737 54723 36740
rect 54665 36731 54723 36737
rect 56594 36728 56600 36740
rect 56652 36728 56658 36780
rect 33134 36700 33140 36712
rect 24259 36672 27016 36700
rect 31726 36672 33140 36700
rect 24259 36669 24271 36672
rect 24213 36663 24271 36669
rect 31726 36632 31754 36672
rect 33134 36660 33140 36672
rect 33192 36660 33198 36712
rect 54389 36703 54447 36709
rect 54389 36669 54401 36703
rect 54435 36669 54447 36703
rect 54570 36700 54576 36712
rect 54531 36672 54576 36700
rect 54389 36663 54447 36669
rect 22066 36604 31754 36632
rect 54404 36632 54432 36663
rect 54570 36660 54576 36672
rect 54628 36660 54634 36712
rect 55122 36632 55128 36644
rect 54404 36604 55128 36632
rect 55122 36592 55128 36604
rect 55180 36592 55186 36644
rect 6641 36567 6699 36573
rect 6641 36533 6653 36567
rect 6687 36533 6699 36567
rect 6641 36527 6699 36533
rect 7101 36567 7159 36573
rect 7101 36533 7113 36567
rect 7147 36564 7159 36567
rect 16666 36564 16672 36576
rect 7147 36536 16672 36564
rect 7147 36533 7159 36536
rect 7101 36527 7159 36533
rect 16666 36524 16672 36536
rect 16724 36524 16730 36576
rect 18141 36567 18199 36573
rect 18141 36533 18153 36567
rect 18187 36564 18199 36567
rect 18874 36564 18880 36576
rect 18187 36536 18880 36564
rect 18187 36533 18199 36536
rect 18141 36527 18199 36533
rect 18874 36524 18880 36536
rect 18932 36524 18938 36576
rect 18966 36524 18972 36576
rect 19024 36564 19030 36576
rect 23842 36564 23848 36576
rect 19024 36536 23848 36564
rect 19024 36524 19030 36536
rect 23842 36524 23848 36536
rect 23900 36524 23906 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 3053 36363 3111 36369
rect 3053 36329 3065 36363
rect 3099 36360 3111 36363
rect 7190 36360 7196 36372
rect 3099 36332 7196 36360
rect 3099 36329 3111 36332
rect 3053 36323 3111 36329
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 7834 36320 7840 36372
rect 7892 36360 7898 36372
rect 16390 36360 16396 36372
rect 7892 36332 16396 36360
rect 7892 36320 7898 36332
rect 16390 36320 16396 36332
rect 16448 36320 16454 36372
rect 19058 36360 19064 36372
rect 18708 36332 19064 36360
rect 1857 36295 1915 36301
rect 1857 36261 1869 36295
rect 1903 36292 1915 36295
rect 18708 36292 18736 36332
rect 19058 36320 19064 36332
rect 19116 36360 19122 36372
rect 32122 36360 32128 36372
rect 19116 36332 19334 36360
rect 19116 36320 19122 36332
rect 18874 36292 18880 36304
rect 1903 36264 6408 36292
rect 1903 36261 1915 36264
rect 1857 36255 1915 36261
rect 2682 36184 2688 36236
rect 2740 36224 2746 36236
rect 2740 36196 2912 36224
rect 2740 36184 2746 36196
rect 2498 36156 2504 36168
rect 2459 36128 2504 36156
rect 2498 36116 2504 36128
rect 2556 36116 2562 36168
rect 2884 36165 2912 36196
rect 5552 36196 6040 36224
rect 5552 36165 5580 36196
rect 2869 36159 2927 36165
rect 2869 36125 2881 36159
rect 2915 36156 2927 36159
rect 5537 36159 5595 36165
rect 2915 36128 5396 36156
rect 2915 36125 2927 36128
rect 2869 36119 2927 36125
rect 1670 36088 1676 36100
rect 1631 36060 1676 36088
rect 1670 36048 1676 36060
rect 1728 36048 1734 36100
rect 2590 36048 2596 36100
rect 2648 36088 2654 36100
rect 2685 36091 2743 36097
rect 2685 36088 2697 36091
rect 2648 36060 2697 36088
rect 2648 36048 2654 36060
rect 2685 36057 2697 36060
rect 2731 36057 2743 36091
rect 2685 36051 2743 36057
rect 2774 36048 2780 36100
rect 2832 36088 2838 36100
rect 2832 36060 2877 36088
rect 2832 36048 2838 36060
rect 5166 36020 5172 36032
rect 5127 35992 5172 36020
rect 5166 35980 5172 35992
rect 5224 35980 5230 36032
rect 5368 36020 5396 36128
rect 5537 36125 5549 36159
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 5626 36116 5632 36168
rect 5684 36156 5690 36168
rect 5902 36156 5908 36168
rect 5684 36128 5729 36156
rect 5863 36128 5908 36156
rect 5684 36116 5690 36128
rect 5902 36116 5908 36128
rect 5960 36116 5966 36168
rect 6012 36088 6040 36196
rect 6178 36156 6184 36168
rect 6139 36128 6184 36156
rect 6178 36116 6184 36128
rect 6236 36116 6242 36168
rect 6380 36165 6408 36264
rect 9646 36264 18736 36292
rect 18835 36264 18880 36292
rect 9646 36224 9674 36264
rect 18874 36252 18880 36264
rect 18932 36252 18938 36304
rect 19306 36292 19334 36332
rect 21192 36332 32128 36360
rect 19426 36292 19432 36304
rect 19306 36264 19432 36292
rect 19426 36252 19432 36264
rect 19484 36252 19490 36304
rect 21192 36301 21220 36332
rect 32122 36320 32128 36332
rect 32180 36320 32186 36372
rect 46198 36360 46204 36372
rect 35866 36332 46204 36360
rect 21177 36295 21235 36301
rect 21177 36261 21189 36295
rect 21223 36261 21235 36295
rect 21177 36255 21235 36261
rect 22462 36252 22468 36304
rect 22520 36292 22526 36304
rect 23290 36292 23296 36304
rect 22520 36264 23296 36292
rect 22520 36252 22526 36264
rect 23290 36252 23296 36264
rect 23348 36252 23354 36304
rect 35866 36224 35894 36332
rect 46198 36320 46204 36332
rect 46256 36320 46262 36372
rect 54018 36360 54024 36372
rect 53979 36332 54024 36360
rect 54018 36320 54024 36332
rect 54076 36320 54082 36372
rect 40770 36224 40776 36236
rect 7116 36196 9674 36224
rect 12406 36196 18828 36224
rect 6365 36159 6423 36165
rect 6365 36125 6377 36159
rect 6411 36125 6423 36159
rect 6365 36119 6423 36125
rect 7006 36088 7012 36100
rect 6012 36060 7012 36088
rect 7006 36048 7012 36060
rect 7064 36048 7070 36100
rect 7116 36020 7144 36196
rect 7190 36116 7196 36168
rect 7248 36156 7254 36168
rect 12406 36156 12434 36196
rect 18800 36168 18828 36196
rect 20180 36196 35894 36224
rect 40328 36196 40776 36224
rect 7248 36128 12434 36156
rect 18049 36159 18107 36165
rect 7248 36116 7254 36128
rect 18049 36125 18061 36159
rect 18095 36156 18107 36159
rect 18322 36156 18328 36168
rect 18095 36128 18328 36156
rect 18095 36125 18107 36128
rect 18049 36119 18107 36125
rect 18322 36116 18328 36128
rect 18380 36116 18386 36168
rect 18598 36156 18604 36168
rect 18559 36128 18604 36156
rect 18598 36116 18604 36128
rect 18656 36116 18662 36168
rect 18693 36159 18751 36165
rect 18693 36125 18705 36159
rect 18739 36125 18751 36159
rect 18693 36119 18751 36125
rect 18509 36091 18567 36097
rect 18509 36057 18521 36091
rect 18555 36057 18567 36091
rect 18708 36088 18736 36119
rect 18782 36116 18788 36168
rect 18840 36116 18846 36168
rect 19978 36156 19984 36168
rect 19939 36128 19984 36156
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 20180 36165 20208 36196
rect 20129 36159 20208 36165
rect 20129 36125 20141 36159
rect 20175 36128 20208 36159
rect 20346 36156 20352 36168
rect 20307 36128 20352 36156
rect 20175 36125 20187 36128
rect 20129 36119 20187 36125
rect 20346 36116 20352 36128
rect 20404 36116 20410 36168
rect 20530 36165 20536 36168
rect 20487 36159 20536 36165
rect 20487 36125 20499 36159
rect 20533 36125 20536 36159
rect 20487 36119 20536 36125
rect 20530 36116 20536 36119
rect 20588 36156 20594 36168
rect 20714 36156 20720 36168
rect 20588 36128 20720 36156
rect 20588 36116 20594 36128
rect 20714 36116 20720 36128
rect 20772 36116 20778 36168
rect 21082 36156 21088 36168
rect 21043 36128 21088 36156
rect 21082 36116 21088 36128
rect 21140 36116 21146 36168
rect 21358 36156 21364 36168
rect 21319 36128 21364 36156
rect 21358 36116 21364 36128
rect 21416 36116 21422 36168
rect 22462 36156 22468 36168
rect 22423 36128 22468 36156
rect 22462 36116 22468 36128
rect 22520 36116 22526 36168
rect 22741 36159 22799 36165
rect 22741 36156 22753 36159
rect 22572 36128 22753 36156
rect 19886 36088 19892 36100
rect 18708 36060 19892 36088
rect 18509 36051 18567 36057
rect 5368 35992 7144 36020
rect 18524 36020 18552 36051
rect 19886 36048 19892 36060
rect 19944 36048 19950 36100
rect 20257 36091 20315 36097
rect 20257 36057 20269 36091
rect 20303 36088 20315 36091
rect 20806 36088 20812 36100
rect 20303 36060 20812 36088
rect 20303 36057 20315 36060
rect 20257 36051 20315 36057
rect 20806 36048 20812 36060
rect 20864 36048 20870 36100
rect 22278 36048 22284 36100
rect 22336 36088 22342 36100
rect 22572 36088 22600 36128
rect 22741 36125 22753 36128
rect 22787 36125 22799 36159
rect 22741 36119 22799 36125
rect 22830 36116 22836 36168
rect 22888 36156 22894 36168
rect 23658 36156 23664 36168
rect 22888 36128 22933 36156
rect 23619 36128 23664 36156
rect 22888 36116 22894 36128
rect 23658 36116 23664 36128
rect 23716 36116 23722 36168
rect 40328 36165 40356 36196
rect 40770 36184 40776 36196
rect 40828 36184 40834 36236
rect 40313 36159 40371 36165
rect 40313 36125 40325 36159
rect 40359 36125 40371 36159
rect 40678 36156 40684 36168
rect 40639 36128 40684 36156
rect 40313 36119 40371 36125
rect 40678 36116 40684 36128
rect 40736 36116 40742 36168
rect 53466 36156 53472 36168
rect 53427 36128 53472 36156
rect 53466 36116 53472 36128
rect 53524 36116 53530 36168
rect 53742 36156 53748 36168
rect 53703 36128 53748 36156
rect 53742 36116 53748 36128
rect 53800 36116 53806 36168
rect 53889 36159 53947 36165
rect 53889 36125 53901 36159
rect 53935 36156 53947 36159
rect 54570 36156 54576 36168
rect 53935 36128 54576 36156
rect 53935 36125 53947 36128
rect 53889 36119 53947 36125
rect 54570 36116 54576 36128
rect 54628 36116 54634 36168
rect 22336 36060 22600 36088
rect 22336 36048 22342 36060
rect 22646 36048 22652 36100
rect 22704 36088 22710 36100
rect 23474 36088 23480 36100
rect 22704 36060 22749 36088
rect 23435 36060 23480 36088
rect 22704 36048 22710 36060
rect 23474 36048 23480 36060
rect 23532 36048 23538 36100
rect 24026 36088 24032 36100
rect 23987 36060 24032 36088
rect 24026 36048 24032 36060
rect 24084 36048 24090 36100
rect 38562 36048 38568 36100
rect 38620 36088 38626 36100
rect 40497 36091 40555 36097
rect 40497 36088 40509 36091
rect 38620 36060 40509 36088
rect 38620 36048 38626 36060
rect 40497 36057 40509 36060
rect 40543 36057 40555 36091
rect 40497 36051 40555 36057
rect 40589 36091 40647 36097
rect 40589 36057 40601 36091
rect 40635 36088 40647 36091
rect 41690 36088 41696 36100
rect 40635 36060 41696 36088
rect 40635 36057 40647 36060
rect 40589 36051 40647 36057
rect 41690 36048 41696 36060
rect 41748 36048 41754 36100
rect 52822 36048 52828 36100
rect 52880 36088 52886 36100
rect 53650 36088 53656 36100
rect 52880 36060 53656 36088
rect 52880 36048 52886 36060
rect 53650 36048 53656 36060
rect 53708 36048 53714 36100
rect 57974 36088 57980 36100
rect 57935 36060 57980 36088
rect 57974 36048 57980 36060
rect 58032 36048 58038 36100
rect 58342 36088 58348 36100
rect 58303 36060 58348 36088
rect 58342 36048 58348 36060
rect 58400 36048 58406 36100
rect 20162 36020 20168 36032
rect 18524 35992 20168 36020
rect 20162 35980 20168 35992
rect 20220 35980 20226 36032
rect 20625 36023 20683 36029
rect 20625 35989 20637 36023
rect 20671 36020 20683 36023
rect 20714 36020 20720 36032
rect 20671 35992 20720 36020
rect 20671 35989 20683 35992
rect 20625 35983 20683 35989
rect 20714 35980 20720 35992
rect 20772 35980 20778 36032
rect 21542 36020 21548 36032
rect 21503 35992 21548 36020
rect 21542 35980 21548 35992
rect 21600 35980 21606 36032
rect 23017 36023 23075 36029
rect 23017 35989 23029 36023
rect 23063 36020 23075 36023
rect 23658 36020 23664 36032
rect 23063 35992 23664 36020
rect 23063 35989 23075 35992
rect 23017 35983 23075 35989
rect 23658 35980 23664 35992
rect 23716 35980 23722 36032
rect 37274 35980 37280 36032
rect 37332 36020 37338 36032
rect 40865 36023 40923 36029
rect 40865 36020 40877 36023
rect 37332 35992 40877 36020
rect 37332 35980 37338 35992
rect 40865 35989 40877 35992
rect 40911 35989 40923 36023
rect 40865 35983 40923 35989
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 20254 35816 20260 35828
rect 19536 35788 20260 35816
rect 1857 35751 1915 35757
rect 1857 35717 1869 35751
rect 1903 35748 1915 35751
rect 2314 35748 2320 35760
rect 1903 35720 2320 35748
rect 1903 35717 1915 35720
rect 1857 35711 1915 35717
rect 2314 35708 2320 35720
rect 2372 35708 2378 35760
rect 1670 35680 1676 35692
rect 1631 35652 1676 35680
rect 1670 35640 1676 35652
rect 1728 35640 1734 35692
rect 19536 35689 19564 35788
rect 20254 35776 20260 35788
rect 20312 35776 20318 35828
rect 23474 35776 23480 35828
rect 23532 35816 23538 35828
rect 24305 35819 24363 35825
rect 24305 35816 24317 35819
rect 23532 35788 24317 35816
rect 23532 35776 23538 35788
rect 24305 35785 24317 35788
rect 24351 35785 24363 35819
rect 24305 35779 24363 35785
rect 26142 35776 26148 35828
rect 26200 35816 26206 35828
rect 34422 35816 34428 35828
rect 26200 35788 34428 35816
rect 26200 35776 26206 35788
rect 34422 35776 34428 35788
rect 34480 35776 34486 35828
rect 19797 35751 19855 35757
rect 19797 35748 19809 35751
rect 19628 35720 19809 35748
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 19521 35643 19579 35649
rect 19334 35572 19340 35624
rect 19392 35612 19398 35624
rect 19628 35612 19656 35720
rect 19797 35717 19809 35720
rect 19843 35717 19855 35751
rect 23201 35751 23259 35757
rect 23201 35748 23213 35751
rect 19797 35711 19855 35717
rect 19904 35720 23213 35748
rect 19904 35689 19932 35720
rect 23201 35717 23213 35720
rect 23247 35748 23259 35751
rect 23750 35748 23756 35760
rect 23247 35720 23756 35748
rect 23247 35717 23259 35720
rect 23201 35711 23259 35717
rect 23750 35708 23756 35720
rect 23808 35708 23814 35760
rect 23845 35751 23903 35757
rect 23845 35717 23857 35751
rect 23891 35748 23903 35751
rect 37274 35748 37280 35760
rect 23891 35720 37280 35748
rect 23891 35717 23903 35720
rect 23845 35711 23903 35717
rect 37274 35708 37280 35720
rect 37332 35708 37338 35760
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35649 19763 35683
rect 19705 35643 19763 35649
rect 19889 35683 19947 35689
rect 19889 35649 19901 35683
rect 19935 35649 19947 35683
rect 19889 35643 19947 35649
rect 20625 35683 20683 35689
rect 20625 35649 20637 35683
rect 20671 35680 20683 35683
rect 22186 35680 22192 35692
rect 20671 35652 22094 35680
rect 22147 35652 22192 35680
rect 20671 35649 20683 35652
rect 20625 35643 20683 35649
rect 19392 35584 19656 35612
rect 19392 35572 19398 35584
rect 19720 35544 19748 35643
rect 20070 35572 20076 35624
rect 20128 35612 20134 35624
rect 20530 35612 20536 35624
rect 20128 35584 20536 35612
rect 20128 35572 20134 35584
rect 20530 35572 20536 35584
rect 20588 35612 20594 35624
rect 21177 35615 21235 35621
rect 21177 35612 21189 35615
rect 20588 35584 21189 35612
rect 20588 35572 20594 35584
rect 21177 35581 21189 35584
rect 21223 35612 21235 35615
rect 21223 35584 21956 35612
rect 21223 35581 21235 35584
rect 21177 35575 21235 35581
rect 19886 35544 19892 35556
rect 19720 35516 19892 35544
rect 19886 35504 19892 35516
rect 19944 35504 19950 35556
rect 21358 35544 21364 35556
rect 19996 35516 21364 35544
rect 15838 35436 15844 35488
rect 15896 35476 15902 35488
rect 19996 35476 20024 35516
rect 21358 35504 21364 35516
rect 21416 35504 21422 35556
rect 15896 35448 20024 35476
rect 20073 35479 20131 35485
rect 15896 35436 15902 35448
rect 20073 35445 20085 35479
rect 20119 35476 20131 35479
rect 21818 35476 21824 35488
rect 20119 35448 21824 35476
rect 20119 35445 20131 35448
rect 20073 35439 20131 35445
rect 21818 35436 21824 35448
rect 21876 35436 21882 35488
rect 21928 35476 21956 35584
rect 22066 35544 22094 35652
rect 22186 35640 22192 35652
rect 22244 35640 22250 35692
rect 24118 35680 24124 35692
rect 24079 35652 24124 35680
rect 24118 35640 24124 35652
rect 24176 35640 24182 35692
rect 33134 35640 33140 35692
rect 33192 35680 33198 35692
rect 35989 35683 36047 35689
rect 35989 35680 36001 35683
rect 33192 35652 36001 35680
rect 33192 35640 33198 35652
rect 35989 35649 36001 35652
rect 36035 35649 36047 35683
rect 35989 35643 36047 35649
rect 23658 35572 23664 35624
rect 23716 35612 23722 35624
rect 23937 35615 23995 35621
rect 23937 35612 23949 35615
rect 23716 35584 23949 35612
rect 23716 35572 23722 35584
rect 23937 35581 23949 35584
rect 23983 35581 23995 35615
rect 23937 35575 23995 35581
rect 36170 35572 36176 35624
rect 36228 35612 36234 35624
rect 36265 35615 36323 35621
rect 36265 35612 36277 35615
rect 36228 35584 36277 35612
rect 36228 35572 36234 35584
rect 36265 35581 36277 35584
rect 36311 35612 36323 35615
rect 40678 35612 40684 35624
rect 36311 35584 40684 35612
rect 36311 35581 36323 35584
rect 36265 35575 36323 35581
rect 40678 35572 40684 35584
rect 40736 35572 40742 35624
rect 22066 35516 23980 35544
rect 23952 35488 23980 35516
rect 35986 35504 35992 35556
rect 36044 35544 36050 35556
rect 36188 35544 36216 35572
rect 36044 35516 36216 35544
rect 36044 35504 36050 35516
rect 22738 35476 22744 35488
rect 21928 35448 22744 35476
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 23842 35476 23848 35488
rect 23803 35448 23848 35476
rect 23842 35436 23848 35448
rect 23900 35436 23906 35488
rect 23934 35436 23940 35488
rect 23992 35436 23998 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 19978 35232 19984 35284
rect 20036 35272 20042 35284
rect 20073 35275 20131 35281
rect 20073 35272 20085 35275
rect 20036 35244 20085 35272
rect 20036 35232 20042 35244
rect 20073 35241 20085 35244
rect 20119 35241 20131 35275
rect 21818 35272 21824 35284
rect 21779 35244 21824 35272
rect 20073 35235 20131 35241
rect 21818 35232 21824 35244
rect 21876 35232 21882 35284
rect 43438 35232 43444 35284
rect 43496 35272 43502 35284
rect 50154 35272 50160 35284
rect 43496 35244 50160 35272
rect 43496 35232 43502 35244
rect 50154 35232 50160 35244
rect 50212 35232 50218 35284
rect 1857 35207 1915 35213
rect 1857 35173 1869 35207
rect 1903 35204 1915 35207
rect 2774 35204 2780 35216
rect 1903 35176 2780 35204
rect 1903 35173 1915 35176
rect 1857 35167 1915 35173
rect 2774 35164 2780 35176
rect 2832 35164 2838 35216
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 20714 35204 20720 35216
rect 16724 35176 20484 35204
rect 20675 35176 20720 35204
rect 16724 35164 16730 35176
rect 20349 35139 20407 35145
rect 20349 35136 20361 35139
rect 19536 35108 20361 35136
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 19536 35077 19564 35108
rect 20349 35105 20361 35108
rect 20395 35105 20407 35139
rect 20349 35099 20407 35105
rect 19521 35071 19579 35077
rect 19521 35068 19533 35071
rect 19392 35040 19533 35068
rect 19392 35028 19398 35040
rect 19521 35037 19533 35040
rect 19567 35037 19579 35071
rect 19797 35071 19855 35077
rect 19797 35068 19809 35071
rect 19521 35031 19579 35037
rect 19628 35040 19809 35068
rect 1670 35000 1676 35012
rect 1631 34972 1676 35000
rect 1670 34960 1676 34972
rect 1728 34960 1734 35012
rect 12158 34960 12164 35012
rect 12216 35000 12222 35012
rect 19628 35000 19656 35040
rect 19797 35037 19809 35040
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 19889 35071 19947 35077
rect 19889 35037 19901 35071
rect 19935 35037 19947 35071
rect 20456 35068 20484 35176
rect 20714 35164 20720 35176
rect 20772 35164 20778 35216
rect 23658 35204 23664 35216
rect 20916 35176 23664 35204
rect 20916 35077 20944 35176
rect 23658 35164 23664 35176
rect 23716 35204 23722 35216
rect 24762 35204 24768 35216
rect 23716 35176 24768 35204
rect 23716 35164 23722 35176
rect 24762 35164 24768 35176
rect 24820 35164 24826 35216
rect 35621 35207 35679 35213
rect 35621 35173 35633 35207
rect 35667 35204 35679 35207
rect 36998 35204 37004 35216
rect 35667 35176 37004 35204
rect 35667 35173 35679 35176
rect 35621 35167 35679 35173
rect 36998 35164 37004 35176
rect 37056 35164 37062 35216
rect 40589 35207 40647 35213
rect 40589 35173 40601 35207
rect 40635 35173 40647 35207
rect 40589 35167 40647 35173
rect 22005 35139 22063 35145
rect 22005 35105 22017 35139
rect 22051 35136 22063 35139
rect 40604 35136 40632 35167
rect 44818 35164 44824 35216
rect 44876 35204 44882 35216
rect 58618 35204 58624 35216
rect 44876 35176 58624 35204
rect 44876 35164 44882 35176
rect 58618 35164 58624 35176
rect 58676 35164 58682 35216
rect 22051 35108 40632 35136
rect 22051 35105 22063 35108
rect 22005 35099 22063 35105
rect 20625 35071 20683 35077
rect 20625 35068 20637 35071
rect 20456 35040 20637 35068
rect 19889 35031 19947 35037
rect 20625 35037 20637 35040
rect 20671 35037 20683 35071
rect 20625 35031 20683 35037
rect 20901 35071 20959 35077
rect 20901 35037 20913 35071
rect 20947 35037 20959 35071
rect 20901 35031 20959 35037
rect 12216 34972 19656 35000
rect 12216 34960 12222 34972
rect 19702 34960 19708 35012
rect 19760 35000 19766 35012
rect 19904 35000 19932 35031
rect 21358 35028 21364 35080
rect 21416 35068 21422 35080
rect 21821 35071 21879 35077
rect 21821 35068 21833 35071
rect 21416 35040 21833 35068
rect 21416 35028 21422 35040
rect 21821 35037 21833 35040
rect 21867 35037 21879 35071
rect 21821 35031 21879 35037
rect 22094 35028 22100 35080
rect 22152 35068 22158 35080
rect 22646 35068 22652 35080
rect 22152 35040 22652 35068
rect 22152 35028 22158 35040
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 24762 35028 24768 35080
rect 24820 35068 24826 35080
rect 35986 35068 35992 35080
rect 24820 35040 35756 35068
rect 35947 35040 35992 35068
rect 24820 35028 24826 35040
rect 26142 35000 26148 35012
rect 19760 34972 19805 35000
rect 19904 34972 21220 35000
rect 19760 34960 19766 34972
rect 21082 34932 21088 34944
rect 21043 34904 21088 34932
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 21192 34932 21220 34972
rect 22066 34972 26148 35000
rect 22066 34932 22094 34972
rect 26142 34960 26148 34972
rect 26200 34960 26206 35012
rect 21192 34904 22094 34932
rect 22281 34935 22339 34941
rect 22281 34901 22293 34935
rect 22327 34932 22339 34935
rect 22462 34932 22468 34944
rect 22327 34904 22468 34932
rect 22327 34901 22339 34904
rect 22281 34895 22339 34901
rect 22462 34892 22468 34904
rect 22520 34892 22526 34944
rect 35728 34932 35756 35040
rect 35986 35028 35992 35040
rect 36044 35028 36050 35080
rect 36078 35028 36084 35080
rect 36136 35068 36142 35080
rect 36357 35071 36415 35077
rect 36136 35040 36181 35068
rect 36136 35028 36142 35040
rect 36357 35037 36369 35071
rect 36403 35037 36415 35071
rect 36357 35031 36415 35037
rect 36633 35071 36691 35077
rect 36633 35037 36645 35071
rect 36679 35037 36691 35071
rect 36814 35068 36820 35080
rect 36775 35040 36820 35068
rect 36633 35031 36691 35037
rect 36372 34932 36400 35031
rect 36648 35000 36676 35031
rect 36814 35028 36820 35040
rect 36872 35028 36878 35080
rect 40037 35071 40095 35077
rect 40037 35037 40049 35071
rect 40083 35037 40095 35071
rect 40310 35068 40316 35080
rect 40271 35040 40316 35068
rect 40037 35031 40095 35037
rect 37366 35000 37372 35012
rect 36648 34972 37372 35000
rect 37366 34960 37372 34972
rect 37424 34960 37430 35012
rect 35728 34904 36400 34932
rect 40052 34932 40080 35031
rect 40310 35028 40316 35040
rect 40368 35028 40374 35080
rect 40405 35071 40463 35077
rect 40405 35037 40417 35071
rect 40451 35068 40463 35071
rect 40678 35068 40684 35080
rect 40451 35040 40684 35068
rect 40451 35037 40463 35040
rect 40405 35031 40463 35037
rect 40678 35028 40684 35040
rect 40736 35028 40742 35080
rect 47762 35028 47768 35080
rect 47820 35068 47826 35080
rect 57885 35071 57943 35077
rect 57885 35068 57897 35071
rect 47820 35040 57897 35068
rect 47820 35028 47826 35040
rect 57885 35037 57897 35040
rect 57931 35037 57943 35071
rect 57885 35031 57943 35037
rect 40218 35000 40224 35012
rect 40179 34972 40224 35000
rect 40218 34960 40224 34972
rect 40276 34960 40282 35012
rect 58158 35000 58164 35012
rect 58119 34972 58164 35000
rect 58158 34960 58164 34972
rect 58216 34960 58222 35012
rect 45094 34932 45100 34944
rect 40052 34904 45100 34932
rect 45094 34892 45100 34904
rect 45152 34892 45158 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 22370 34688 22376 34740
rect 22428 34728 22434 34740
rect 22428 34700 22508 34728
rect 22428 34688 22434 34700
rect 22480 34669 22508 34700
rect 23842 34688 23848 34740
rect 23900 34728 23906 34740
rect 23937 34731 23995 34737
rect 23937 34728 23949 34731
rect 23900 34700 23949 34728
rect 23900 34688 23906 34700
rect 23937 34697 23949 34700
rect 23983 34697 23995 34731
rect 37366 34728 37372 34740
rect 23937 34691 23995 34697
rect 24044 34700 26469 34728
rect 22465 34663 22523 34669
rect 22465 34629 22477 34663
rect 22511 34629 22523 34663
rect 22465 34623 22523 34629
rect 22738 34620 22744 34672
rect 22796 34660 22802 34672
rect 22796 34632 23796 34660
rect 22796 34620 22802 34632
rect 22094 34592 22100 34604
rect 22055 34564 22100 34592
rect 22094 34552 22100 34564
rect 22152 34552 22158 34604
rect 22278 34601 22284 34604
rect 22245 34595 22284 34601
rect 22245 34561 22257 34595
rect 22245 34555 22284 34561
rect 22278 34552 22284 34555
rect 22336 34552 22342 34604
rect 22373 34595 22431 34601
rect 22373 34561 22385 34595
rect 22419 34561 22431 34595
rect 22554 34592 22560 34604
rect 22513 34564 22560 34592
rect 22373 34555 22431 34561
rect 20806 34416 20812 34468
rect 20864 34456 20870 34468
rect 22388 34456 22416 34555
rect 22554 34552 22560 34564
rect 22612 34601 22618 34604
rect 22612 34595 22661 34601
rect 22612 34561 22615 34595
rect 22649 34592 22661 34595
rect 22830 34592 22836 34604
rect 22649 34564 22836 34592
rect 22649 34561 22661 34564
rect 22612 34555 22661 34561
rect 22612 34552 22618 34555
rect 22830 34552 22836 34564
rect 22888 34552 22894 34604
rect 23385 34595 23443 34601
rect 23385 34561 23397 34595
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 22738 34484 22744 34536
rect 22796 34524 22802 34536
rect 23017 34527 23075 34533
rect 23017 34524 23029 34527
rect 22796 34496 23029 34524
rect 22796 34484 22802 34496
rect 23017 34493 23029 34496
rect 23063 34524 23075 34527
rect 23400 34524 23428 34555
rect 23474 34552 23480 34604
rect 23532 34592 23538 34604
rect 23768 34601 23796 34632
rect 23569 34595 23627 34601
rect 23569 34592 23581 34595
rect 23532 34564 23581 34592
rect 23532 34552 23538 34564
rect 23569 34561 23581 34564
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 23661 34595 23719 34601
rect 23661 34561 23673 34595
rect 23707 34561 23719 34595
rect 23661 34555 23719 34561
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 24044 34592 24072 34700
rect 26326 34660 26332 34672
rect 26287 34632 26332 34660
rect 26326 34620 26332 34632
rect 26384 34620 26390 34672
rect 25958 34592 25964 34604
rect 23799 34564 24072 34592
rect 25919 34564 25964 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 23063 34496 23428 34524
rect 23676 34524 23704 34555
rect 25958 34552 25964 34564
rect 26016 34552 26022 34604
rect 26142 34601 26148 34604
rect 26109 34595 26148 34601
rect 26109 34561 26121 34595
rect 26109 34555 26148 34561
rect 26142 34552 26148 34555
rect 26200 34552 26206 34604
rect 26441 34601 26469 34700
rect 26528 34700 37372 34728
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34561 26295 34595
rect 26237 34555 26295 34561
rect 26426 34595 26484 34601
rect 26426 34561 26438 34595
rect 26472 34561 26484 34595
rect 26426 34555 26484 34561
rect 24486 34524 24492 34536
rect 23676 34496 24492 34524
rect 23063 34493 23075 34496
rect 23017 34487 23075 34493
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 24670 34484 24676 34536
rect 24728 34524 24734 34536
rect 26252 34524 26280 34555
rect 26528 34524 26556 34700
rect 37366 34688 37372 34700
rect 37424 34688 37430 34740
rect 50706 34688 50712 34740
rect 50764 34728 50770 34740
rect 57790 34728 57796 34740
rect 50764 34700 57796 34728
rect 50764 34688 50770 34700
rect 57790 34688 57796 34700
rect 57848 34688 57854 34740
rect 57974 34688 57980 34740
rect 58032 34728 58038 34740
rect 58253 34731 58311 34737
rect 58253 34728 58265 34731
rect 58032 34700 58265 34728
rect 58032 34688 58038 34700
rect 58253 34697 58265 34700
rect 58299 34697 58311 34731
rect 58253 34691 58311 34697
rect 26878 34620 26884 34672
rect 26936 34660 26942 34672
rect 40218 34660 40224 34672
rect 26936 34632 40224 34660
rect 26936 34620 26942 34632
rect 40218 34620 40224 34632
rect 40276 34620 40282 34672
rect 57882 34552 57888 34604
rect 57940 34592 57946 34604
rect 58069 34595 58127 34601
rect 58069 34592 58081 34595
rect 57940 34564 58081 34592
rect 57940 34552 57946 34564
rect 58069 34561 58081 34564
rect 58115 34561 58127 34595
rect 58069 34555 58127 34561
rect 24728 34496 26280 34524
rect 26344 34496 26556 34524
rect 24728 34484 24734 34496
rect 23198 34456 23204 34468
rect 20864 34428 23204 34456
rect 20864 34416 20870 34428
rect 23198 34416 23204 34428
rect 23256 34416 23262 34468
rect 26050 34416 26056 34468
rect 26108 34456 26114 34468
rect 26344 34456 26372 34496
rect 33594 34484 33600 34536
rect 33652 34524 33658 34536
rect 34422 34524 34428 34536
rect 33652 34496 34428 34524
rect 33652 34484 33658 34496
rect 34422 34484 34428 34496
rect 34480 34484 34486 34536
rect 26108 34428 26372 34456
rect 26108 34416 26114 34428
rect 19426 34348 19432 34400
rect 19484 34388 19490 34400
rect 20346 34388 20352 34400
rect 19484 34360 20352 34388
rect 19484 34348 19490 34360
rect 20346 34348 20352 34360
rect 20404 34388 20410 34400
rect 21266 34388 21272 34400
rect 20404 34360 21272 34388
rect 20404 34348 20410 34360
rect 21266 34348 21272 34360
rect 21324 34348 21330 34400
rect 22094 34348 22100 34400
rect 22152 34388 22158 34400
rect 22741 34391 22799 34397
rect 22741 34388 22753 34391
rect 22152 34360 22753 34388
rect 22152 34348 22158 34360
rect 22741 34357 22753 34360
rect 22787 34357 22799 34391
rect 26602 34388 26608 34400
rect 26563 34360 26608 34388
rect 22741 34351 22799 34357
rect 26602 34348 26608 34360
rect 26660 34348 26666 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 31754 34184 31760 34196
rect 21192 34156 31760 34184
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20680 33952 20821 33980
rect 20680 33940 20686 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 20957 33983 21015 33989
rect 20957 33949 20969 33983
rect 21003 33980 21015 33983
rect 21192 33980 21220 34156
rect 31754 34144 31760 34156
rect 31812 34144 31818 34196
rect 21453 34119 21511 34125
rect 21453 34085 21465 34119
rect 21499 34085 21511 34119
rect 21453 34079 21511 34085
rect 21003 33952 21220 33980
rect 21003 33949 21015 33952
rect 20957 33943 21015 33949
rect 21266 33940 21272 33992
rect 21324 33989 21330 33992
rect 21324 33980 21332 33989
rect 21468 33980 21496 34079
rect 22554 34048 22560 34060
rect 22515 34020 22560 34048
rect 22554 34008 22560 34020
rect 22612 34008 22618 34060
rect 22005 33983 22063 33989
rect 22005 33980 22017 33983
rect 21324 33952 21369 33980
rect 21468 33952 22017 33980
rect 21324 33943 21332 33952
rect 22005 33949 22017 33952
rect 22051 33949 22063 33983
rect 22462 33980 22468 33992
rect 22423 33952 22468 33980
rect 22005 33943 22063 33949
rect 21324 33940 21330 33943
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 35342 33940 35348 33992
rect 35400 33980 35406 33992
rect 35400 33952 45554 33980
rect 35400 33940 35406 33952
rect 1670 33912 1676 33924
rect 1631 33884 1676 33912
rect 1670 33872 1676 33884
rect 1728 33872 1734 33924
rect 20714 33872 20720 33924
rect 20772 33912 20778 33924
rect 21085 33915 21143 33921
rect 21085 33912 21097 33915
rect 20772 33884 21097 33912
rect 20772 33872 20778 33884
rect 21085 33881 21097 33884
rect 21131 33881 21143 33915
rect 21085 33875 21143 33881
rect 21177 33915 21235 33921
rect 21177 33881 21189 33915
rect 21223 33881 21235 33915
rect 21177 33875 21235 33881
rect 1765 33847 1823 33853
rect 1765 33813 1777 33847
rect 1811 33844 1823 33847
rect 21192 33844 21220 33875
rect 35434 33872 35440 33924
rect 35492 33912 35498 33924
rect 35894 33912 35900 33924
rect 35492 33884 35900 33912
rect 35492 33872 35498 33884
rect 35894 33872 35900 33884
rect 35952 33872 35958 33924
rect 45526 33912 45554 33952
rect 57146 33912 57152 33924
rect 45526 33884 57152 33912
rect 57146 33872 57152 33884
rect 57204 33872 57210 33924
rect 1811 33816 21220 33844
rect 1811 33813 1823 33816
rect 1765 33807 1823 33813
rect 22278 33804 22284 33856
rect 22336 33844 22342 33856
rect 49326 33844 49332 33856
rect 22336 33816 49332 33844
rect 22336 33804 22342 33816
rect 49326 33804 49332 33816
rect 49384 33804 49390 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1857 33575 1915 33581
rect 1857 33541 1869 33575
rect 1903 33572 1915 33575
rect 2130 33572 2136 33584
rect 1903 33544 2136 33572
rect 1903 33541 1915 33544
rect 1857 33535 1915 33541
rect 2130 33532 2136 33544
rect 2188 33532 2194 33584
rect 1670 33504 1676 33516
rect 1631 33476 1676 33504
rect 1670 33464 1676 33476
rect 1728 33464 1734 33516
rect 22002 33504 22008 33516
rect 21963 33476 22008 33504
rect 22002 33464 22008 33476
rect 22060 33464 22066 33516
rect 22094 33464 22100 33516
rect 22152 33504 22158 33516
rect 22281 33507 22339 33513
rect 22152 33476 22197 33504
rect 22152 33464 22158 33476
rect 22281 33473 22293 33507
rect 22327 33504 22339 33507
rect 23658 33504 23664 33516
rect 22327 33476 23664 33504
rect 22327 33473 22339 33476
rect 22281 33467 22339 33473
rect 23658 33464 23664 33476
rect 23716 33504 23722 33516
rect 24762 33504 24768 33516
rect 23716 33476 24768 33504
rect 23716 33464 23722 33476
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 22741 33439 22799 33445
rect 22741 33405 22753 33439
rect 22787 33436 22799 33439
rect 27430 33436 27436 33448
rect 22787 33408 27436 33436
rect 22787 33405 22799 33408
rect 22741 33399 22799 33405
rect 27430 33396 27436 33408
rect 27488 33396 27494 33448
rect 38838 33260 38844 33312
rect 38896 33300 38902 33312
rect 45002 33300 45008 33312
rect 38896 33272 45008 33300
rect 38896 33260 38902 33272
rect 45002 33260 45008 33272
rect 45060 33260 45066 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 19426 33056 19432 33108
rect 19484 33096 19490 33108
rect 28350 33096 28356 33108
rect 19484 33068 28356 33096
rect 19484 33056 19490 33068
rect 28350 33056 28356 33068
rect 28408 33056 28414 33108
rect 26602 32988 26608 33040
rect 26660 33028 26666 33040
rect 26789 33031 26847 33037
rect 26789 33028 26801 33031
rect 26660 33000 26801 33028
rect 26660 32988 26666 33000
rect 26789 32997 26801 33000
rect 26835 32997 26847 33031
rect 26789 32991 26847 32997
rect 16942 32920 16948 32972
rect 17000 32960 17006 32972
rect 21082 32960 21088 32972
rect 17000 32932 21088 32960
rect 17000 32920 17006 32932
rect 21082 32920 21088 32932
rect 21140 32920 21146 32972
rect 21634 32920 21640 32972
rect 21692 32960 21698 32972
rect 22833 32963 22891 32969
rect 22833 32960 22845 32963
rect 21692 32932 22845 32960
rect 21692 32920 21698 32932
rect 22833 32929 22845 32932
rect 22879 32929 22891 32963
rect 58158 32960 58164 32972
rect 58119 32932 58164 32960
rect 22833 32923 22891 32929
rect 58158 32920 58164 32932
rect 58216 32920 58222 32972
rect 22557 32895 22615 32901
rect 22557 32861 22569 32895
rect 22603 32892 22615 32895
rect 23658 32892 23664 32904
rect 22603 32864 23664 32892
rect 22603 32861 22615 32864
rect 22557 32855 22615 32861
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 26694 32892 26700 32904
rect 26655 32864 26700 32892
rect 26694 32852 26700 32864
rect 26752 32852 26758 32904
rect 26970 32892 26976 32904
rect 26931 32864 26976 32892
rect 26970 32852 26976 32864
rect 27028 32852 27034 32904
rect 57698 32852 57704 32904
rect 57756 32892 57762 32904
rect 57885 32895 57943 32901
rect 57885 32892 57897 32895
rect 57756 32864 57897 32892
rect 57756 32852 57762 32864
rect 57885 32861 57897 32864
rect 57931 32861 57943 32895
rect 57885 32855 57943 32861
rect 1670 32824 1676 32836
rect 1631 32796 1676 32824
rect 1670 32784 1676 32796
rect 1728 32784 1734 32836
rect 57054 32824 57060 32836
rect 57015 32796 57060 32824
rect 57054 32784 57060 32796
rect 57112 32784 57118 32836
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 18138 32756 18144 32768
rect 1811 32728 18144 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 18138 32716 18144 32728
rect 18196 32716 18202 32768
rect 27154 32756 27160 32768
rect 27115 32728 27160 32756
rect 27154 32716 27160 32728
rect 27212 32716 27218 32768
rect 57146 32756 57152 32768
rect 57107 32728 57152 32756
rect 57146 32716 57152 32728
rect 57204 32716 57210 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 29914 32512 29920 32564
rect 29972 32552 29978 32564
rect 41598 32552 41604 32564
rect 29972 32524 41604 32552
rect 29972 32512 29978 32524
rect 41598 32512 41604 32524
rect 41656 32512 41662 32564
rect 31754 32444 31760 32496
rect 31812 32484 31818 32496
rect 47394 32484 47400 32496
rect 31812 32456 47400 32484
rect 31812 32444 31818 32456
rect 47394 32444 47400 32456
rect 47452 32444 47458 32496
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 15654 32376 15660 32428
rect 15712 32416 15718 32428
rect 24026 32416 24032 32428
rect 15712 32388 24032 32416
rect 15712 32376 15718 32388
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 26142 32376 26148 32428
rect 26200 32416 26206 32428
rect 53834 32416 53840 32428
rect 26200 32388 53840 32416
rect 26200 32376 26206 32388
rect 53834 32376 53840 32388
rect 53892 32376 53898 32428
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 25314 32212 25320 32224
rect 1811 32184 25320 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 21818 31968 21824 32020
rect 21876 32008 21882 32020
rect 21876 31980 22094 32008
rect 21876 31968 21882 31980
rect 22066 31940 22094 31980
rect 23014 31968 23020 32020
rect 23072 32008 23078 32020
rect 26050 32008 26056 32020
rect 23072 31980 26056 32008
rect 23072 31968 23078 31980
rect 26050 31968 26056 31980
rect 26108 31968 26114 32020
rect 25498 31940 25504 31952
rect 22066 31912 25504 31940
rect 25498 31900 25504 31912
rect 25556 31900 25562 31952
rect 25869 31943 25927 31949
rect 25869 31909 25881 31943
rect 25915 31940 25927 31943
rect 25958 31940 25964 31952
rect 25915 31912 25964 31940
rect 25915 31909 25927 31912
rect 25869 31903 25927 31909
rect 25958 31900 25964 31912
rect 26016 31900 26022 31952
rect 58434 31940 58440 31952
rect 31726 31912 58440 31940
rect 25041 31875 25099 31881
rect 25041 31841 25053 31875
rect 25087 31872 25099 31875
rect 31726 31872 31754 31912
rect 58434 31900 58440 31912
rect 58492 31900 58498 31952
rect 25087 31844 31754 31872
rect 25087 31841 25099 31844
rect 25041 31835 25099 31841
rect 25314 31804 25320 31816
rect 25275 31776 25320 31804
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 25608 31813 25636 31844
rect 44358 31832 44364 31884
rect 44416 31872 44422 31884
rect 44416 31844 45554 31872
rect 44416 31832 44422 31844
rect 25593 31807 25651 31813
rect 25593 31773 25605 31807
rect 25639 31773 25651 31807
rect 25593 31767 25651 31773
rect 25685 31807 25743 31813
rect 25685 31773 25697 31807
rect 25731 31804 25743 31807
rect 26050 31804 26056 31816
rect 25731 31776 26056 31804
rect 25731 31773 25743 31776
rect 25685 31767 25743 31773
rect 26050 31764 26056 31776
rect 26108 31764 26114 31816
rect 45526 31804 45554 31844
rect 57790 31832 57796 31884
rect 57848 31872 57854 31884
rect 58069 31875 58127 31881
rect 58069 31872 58081 31875
rect 57848 31844 58081 31872
rect 57848 31832 57854 31844
rect 58069 31841 58081 31844
rect 58115 31841 58127 31875
rect 58069 31835 58127 31841
rect 57885 31807 57943 31813
rect 57885 31804 57897 31807
rect 45526 31776 57897 31804
rect 57885 31773 57897 31776
rect 57931 31773 57943 31807
rect 57885 31767 57943 31773
rect 22922 31696 22928 31748
rect 22980 31736 22986 31748
rect 25501 31739 25559 31745
rect 25501 31736 25513 31739
rect 22980 31708 25513 31736
rect 22980 31696 22986 31708
rect 25501 31705 25513 31708
rect 25547 31736 25559 31739
rect 25774 31736 25780 31748
rect 25547 31708 25780 31736
rect 25547 31705 25559 31708
rect 25501 31699 25559 31705
rect 25774 31696 25780 31708
rect 25832 31696 25838 31748
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 25961 31467 26019 31473
rect 22066 31436 25728 31464
rect 19518 31356 19524 31408
rect 19576 31396 19582 31408
rect 22066 31396 22094 31436
rect 25590 31396 25596 31408
rect 19576 31368 22094 31396
rect 25551 31368 25596 31396
rect 19576 31356 19582 31368
rect 25590 31356 25596 31368
rect 25648 31356 25654 31408
rect 25700 31405 25728 31436
rect 25961 31433 25973 31467
rect 26007 31464 26019 31467
rect 26694 31464 26700 31476
rect 26007 31436 26700 31464
rect 26007 31433 26019 31436
rect 25961 31427 26019 31433
rect 26694 31424 26700 31436
rect 26752 31424 26758 31476
rect 25685 31399 25743 31405
rect 25685 31365 25697 31399
rect 25731 31365 25743 31399
rect 25685 31359 25743 31365
rect 1670 31328 1676 31340
rect 1631 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19613 31331 19671 31337
rect 19613 31328 19625 31331
rect 19484 31300 19625 31328
rect 19484 31288 19490 31300
rect 19613 31297 19625 31300
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31297 19947 31331
rect 19889 31291 19947 31297
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 19904 31260 19932 31291
rect 22646 31288 22652 31340
rect 22704 31328 22710 31340
rect 25222 31328 25228 31340
rect 22704 31300 25228 31328
rect 22704 31288 22710 31300
rect 25222 31288 25228 31300
rect 25280 31328 25286 31340
rect 25317 31331 25375 31337
rect 25317 31328 25329 31331
rect 25280 31300 25329 31328
rect 25280 31288 25286 31300
rect 25317 31297 25329 31300
rect 25363 31297 25375 31331
rect 25317 31291 25375 31297
rect 25465 31331 25523 31337
rect 25465 31297 25477 31331
rect 25511 31328 25523 31331
rect 25511 31297 25544 31328
rect 25465 31291 25544 31297
rect 20070 31260 20076 31272
rect 18288 31232 19932 31260
rect 20031 31232 20076 31260
rect 18288 31220 18294 31232
rect 20070 31220 20076 31232
rect 20128 31220 20134 31272
rect 25516 31260 25544 31291
rect 25774 31288 25780 31340
rect 25832 31337 25838 31340
rect 25832 31328 25840 31337
rect 46934 31328 46940 31340
rect 25832 31300 25877 31328
rect 31726 31300 46940 31328
rect 25832 31291 25840 31300
rect 25832 31288 25838 31291
rect 31726 31260 31754 31300
rect 46934 31288 46940 31300
rect 46992 31288 46998 31340
rect 58066 31328 58072 31340
rect 58027 31300 58072 31328
rect 58066 31288 58072 31300
rect 58124 31288 58130 31340
rect 25516 31232 31754 31260
rect 19702 31192 19708 31204
rect 19663 31164 19708 31192
rect 19702 31152 19708 31164
rect 19760 31152 19766 31204
rect 27706 31152 27712 31204
rect 27764 31192 27770 31204
rect 57146 31192 57152 31204
rect 27764 31164 57152 31192
rect 27764 31152 27770 31164
rect 57146 31152 57152 31164
rect 57204 31152 57210 31204
rect 1762 31124 1768 31136
rect 1723 31096 1768 31124
rect 1762 31084 1768 31096
rect 1820 31084 1826 31136
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 22646 31124 22652 31136
rect 19484 31096 22652 31124
rect 19484 31084 19490 31096
rect 22646 31084 22652 31096
rect 22704 31084 22710 31136
rect 28258 31084 28264 31136
rect 28316 31124 28322 31136
rect 40954 31124 40960 31136
rect 28316 31096 40960 31124
rect 28316 31084 28322 31096
rect 40954 31084 40960 31096
rect 41012 31084 41018 31136
rect 46474 31084 46480 31136
rect 46532 31124 46538 31136
rect 58253 31127 58311 31133
rect 58253 31124 58265 31127
rect 46532 31096 58265 31124
rect 46532 31084 46538 31096
rect 58253 31093 58265 31096
rect 58299 31093 58311 31127
rect 58253 31087 58311 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1762 30880 1768 30932
rect 1820 30920 1826 30932
rect 19518 30920 19524 30932
rect 1820 30892 19524 30920
rect 1820 30880 1826 30892
rect 19518 30880 19524 30892
rect 19576 30880 19582 30932
rect 19702 30880 19708 30932
rect 19760 30920 19766 30932
rect 20073 30923 20131 30929
rect 20073 30920 20085 30923
rect 19760 30892 20085 30920
rect 19760 30880 19766 30892
rect 20073 30889 20085 30892
rect 20119 30889 20131 30923
rect 20073 30883 20131 30889
rect 25314 30880 25320 30932
rect 25372 30920 25378 30932
rect 25590 30920 25596 30932
rect 25372 30892 25596 30920
rect 25372 30880 25378 30892
rect 25590 30880 25596 30892
rect 25648 30880 25654 30932
rect 19978 30852 19984 30864
rect 19720 30824 19984 30852
rect 19426 30716 19432 30728
rect 19387 30688 19432 30716
rect 19426 30676 19432 30688
rect 19484 30676 19490 30728
rect 19610 30725 19616 30728
rect 19577 30719 19616 30725
rect 19577 30685 19589 30719
rect 19577 30679 19616 30685
rect 19610 30676 19616 30679
rect 19668 30676 19674 30728
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 19720 30657 19748 30824
rect 19978 30812 19984 30824
rect 20036 30852 20042 30864
rect 20162 30852 20168 30864
rect 20036 30824 20168 30852
rect 20036 30812 20042 30824
rect 20162 30812 20168 30824
rect 20220 30812 20226 30864
rect 19935 30719 19993 30725
rect 19935 30685 19947 30719
rect 19981 30716 19993 30719
rect 20346 30716 20352 30728
rect 19981 30688 20352 30716
rect 19981 30685 19993 30688
rect 19935 30679 19993 30685
rect 20346 30676 20352 30688
rect 20404 30716 20410 30728
rect 22922 30716 22928 30728
rect 20404 30688 22928 30716
rect 20404 30676 20410 30688
rect 22922 30676 22928 30688
rect 22980 30676 22986 30728
rect 19705 30651 19763 30657
rect 19705 30617 19717 30651
rect 19751 30617 19763 30651
rect 19705 30611 19763 30617
rect 19797 30651 19855 30657
rect 19797 30617 19809 30651
rect 19843 30617 19855 30651
rect 19797 30611 19855 30617
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 19812 30580 19840 30611
rect 1811 30552 19840 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 22830 30336 22836 30388
rect 22888 30376 22894 30388
rect 24210 30376 24216 30388
rect 22888 30348 24216 30376
rect 22888 30336 22894 30348
rect 24210 30336 24216 30348
rect 24268 30376 24274 30388
rect 24268 30348 25636 30376
rect 24268 30336 24274 30348
rect 5718 30268 5724 30320
rect 5776 30308 5782 30320
rect 23661 30311 23719 30317
rect 5776 30280 22094 30308
rect 5776 30268 5782 30280
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30240 1639 30243
rect 17954 30240 17960 30252
rect 1627 30212 17960 30240
rect 1627 30209 1639 30212
rect 1581 30203 1639 30209
rect 17954 30200 17960 30212
rect 18012 30200 18018 30252
rect 22066 30240 22094 30280
rect 23661 30277 23673 30311
rect 23707 30277 23719 30311
rect 23661 30271 23719 30277
rect 23753 30311 23811 30317
rect 23753 30277 23765 30311
rect 23799 30308 23811 30311
rect 23934 30308 23940 30320
rect 23799 30280 23940 30308
rect 23799 30277 23811 30280
rect 23753 30271 23811 30277
rect 23477 30243 23535 30249
rect 23477 30240 23489 30243
rect 22066 30212 23489 30240
rect 23477 30209 23489 30212
rect 23523 30209 23535 30243
rect 23477 30203 23535 30209
rect 23676 30184 23704 30271
rect 23934 30268 23940 30280
rect 23992 30268 23998 30320
rect 24026 30268 24032 30320
rect 24084 30308 24090 30320
rect 24670 30308 24676 30320
rect 24084 30280 24676 30308
rect 24084 30268 24090 30280
rect 24670 30268 24676 30280
rect 24728 30268 24734 30320
rect 25314 30308 25320 30320
rect 25275 30280 25320 30308
rect 25314 30268 25320 30280
rect 25372 30268 25378 30320
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30240 23903 30243
rect 24486 30240 24492 30252
rect 23891 30212 24492 30240
rect 23891 30209 23903 30212
rect 23845 30203 23903 30209
rect 24486 30200 24492 30212
rect 24544 30200 24550 30252
rect 25130 30200 25136 30252
rect 25188 30240 25194 30252
rect 25409 30243 25467 30249
rect 25188 30212 25233 30240
rect 25188 30200 25194 30212
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 25409 30203 25467 30209
rect 25501 30243 25559 30249
rect 25501 30209 25513 30243
rect 25547 30240 25559 30243
rect 25608 30240 25636 30348
rect 46382 30240 46388 30252
rect 25547 30212 25636 30240
rect 31726 30212 46388 30240
rect 25547 30209 25559 30212
rect 25501 30203 25559 30209
rect 1762 30172 1768 30184
rect 1723 30144 1768 30172
rect 1762 30132 1768 30144
rect 1820 30132 1826 30184
rect 4062 30132 4068 30184
rect 4120 30172 4126 30184
rect 4120 30144 19334 30172
rect 4120 30132 4126 30144
rect 19306 30104 19334 30144
rect 23658 30132 23664 30184
rect 23716 30132 23722 30184
rect 25424 30172 25452 30203
rect 25240 30144 25452 30172
rect 25240 30104 25268 30144
rect 25682 30132 25688 30184
rect 25740 30172 25746 30184
rect 31726 30172 31754 30212
rect 46382 30200 46388 30212
rect 46440 30200 46446 30252
rect 44726 30172 44732 30184
rect 25740 30144 31754 30172
rect 35866 30144 44732 30172
rect 25740 30132 25746 30144
rect 19306 30076 25268 30104
rect 26326 30064 26332 30116
rect 26384 30104 26390 30116
rect 35866 30104 35894 30144
rect 44726 30132 44732 30144
rect 44784 30132 44790 30184
rect 26384 30076 35894 30104
rect 26384 30064 26390 30076
rect 24029 30039 24087 30045
rect 24029 30005 24041 30039
rect 24075 30036 24087 30039
rect 24302 30036 24308 30048
rect 24075 30008 24308 30036
rect 24075 30005 24087 30008
rect 24029 29999 24087 30005
rect 24302 29996 24308 30008
rect 24360 29996 24366 30048
rect 24762 29996 24768 30048
rect 24820 30036 24826 30048
rect 25130 30036 25136 30048
rect 24820 30008 25136 30036
rect 24820 29996 24826 30008
rect 25130 29996 25136 30008
rect 25188 29996 25194 30048
rect 25685 30039 25743 30045
rect 25685 30005 25697 30039
rect 25731 30036 25743 30039
rect 25866 30036 25872 30048
rect 25731 30008 25872 30036
rect 25731 30005 25743 30008
rect 25685 29999 25743 30005
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 22646 29792 22652 29844
rect 22704 29832 22710 29844
rect 23474 29832 23480 29844
rect 22704 29804 23480 29832
rect 22704 29792 22710 29804
rect 23474 29792 23480 29804
rect 23532 29832 23538 29844
rect 25866 29832 25872 29844
rect 23532 29804 24532 29832
rect 25827 29804 25872 29832
rect 23532 29792 23538 29804
rect 24504 29776 24532 29804
rect 25866 29792 25872 29804
rect 25924 29792 25930 29844
rect 25958 29792 25964 29844
rect 26016 29832 26022 29844
rect 26016 29804 26061 29832
rect 26016 29792 26022 29804
rect 20162 29724 20168 29776
rect 20220 29764 20226 29776
rect 23934 29764 23940 29776
rect 20220 29736 23940 29764
rect 20220 29724 20226 29736
rect 23934 29724 23940 29736
rect 23992 29724 23998 29776
rect 24026 29724 24032 29776
rect 24084 29764 24090 29776
rect 24084 29736 24129 29764
rect 24084 29724 24090 29736
rect 24486 29724 24492 29776
rect 24544 29764 24550 29776
rect 24544 29736 26372 29764
rect 24544 29724 24550 29736
rect 18690 29656 18696 29708
rect 18748 29696 18754 29708
rect 18748 29668 24992 29696
rect 18748 29656 18754 29668
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 16390 29628 16396 29640
rect 1627 29600 16396 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 16390 29588 16396 29600
rect 16448 29588 16454 29640
rect 23474 29628 23480 29640
rect 23435 29600 23480 29628
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 23842 29628 23848 29640
rect 23803 29600 23848 29628
rect 23842 29588 23848 29600
rect 23900 29588 23906 29640
rect 24578 29628 24584 29640
rect 24539 29600 24584 29628
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 24854 29628 24860 29640
rect 24815 29600 24860 29628
rect 24854 29588 24860 29600
rect 24912 29588 24918 29640
rect 24964 29637 24992 29668
rect 25130 29656 25136 29708
rect 25188 29696 25194 29708
rect 25188 29668 26004 29696
rect 25188 29656 25194 29668
rect 25976 29640 26004 29668
rect 24949 29631 25007 29637
rect 24949 29597 24961 29631
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 25958 29588 25964 29640
rect 26016 29628 26022 29640
rect 26053 29631 26111 29637
rect 26053 29628 26065 29631
rect 26016 29600 26065 29628
rect 26016 29588 26022 29600
rect 26053 29597 26065 29600
rect 26099 29597 26111 29631
rect 26053 29591 26111 29597
rect 26142 29588 26148 29640
rect 26200 29628 26206 29640
rect 26344 29637 26372 29736
rect 58158 29696 58164 29708
rect 58119 29668 58164 29696
rect 58158 29656 58164 29668
rect 58216 29656 58222 29708
rect 26329 29631 26387 29637
rect 26200 29600 26245 29628
rect 26200 29588 26206 29600
rect 26329 29597 26341 29631
rect 26375 29597 26387 29631
rect 26329 29591 26387 29597
rect 57790 29588 57796 29640
rect 57848 29628 57854 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 57848 29600 57897 29628
rect 57848 29588 57854 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 1854 29560 1860 29572
rect 1815 29532 1860 29560
rect 1854 29520 1860 29532
rect 1912 29520 1918 29572
rect 23198 29520 23204 29572
rect 23256 29560 23262 29572
rect 23661 29563 23719 29569
rect 23661 29560 23673 29563
rect 23256 29532 23673 29560
rect 23256 29520 23262 29532
rect 23661 29529 23673 29532
rect 23707 29529 23719 29563
rect 23661 29523 23719 29529
rect 23753 29563 23811 29569
rect 23753 29529 23765 29563
rect 23799 29560 23811 29563
rect 24394 29560 24400 29572
rect 23799 29532 24400 29560
rect 23799 29529 23811 29532
rect 23753 29523 23811 29529
rect 24394 29520 24400 29532
rect 24452 29520 24458 29572
rect 24670 29520 24676 29572
rect 24728 29560 24734 29572
rect 24765 29563 24823 29569
rect 24765 29560 24777 29563
rect 24728 29532 24777 29560
rect 24728 29520 24734 29532
rect 24765 29529 24777 29532
rect 24811 29529 24823 29563
rect 25314 29560 25320 29572
rect 24765 29523 24823 29529
rect 24872 29532 25320 29560
rect 20070 29452 20076 29504
rect 20128 29492 20134 29504
rect 24872 29492 24900 29532
rect 25314 29520 25320 29532
rect 25372 29520 25378 29572
rect 57054 29560 57060 29572
rect 57015 29532 57060 29560
rect 57054 29520 57060 29532
rect 57112 29520 57118 29572
rect 25130 29492 25136 29504
rect 20128 29464 24900 29492
rect 25091 29464 25136 29492
rect 20128 29452 20134 29464
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 25590 29492 25596 29504
rect 25551 29464 25596 29492
rect 25590 29452 25596 29464
rect 25648 29452 25654 29504
rect 30926 29452 30932 29504
rect 30984 29492 30990 29504
rect 57149 29495 57207 29501
rect 57149 29492 57161 29495
rect 30984 29464 57161 29492
rect 30984 29452 30990 29464
rect 57149 29461 57161 29464
rect 57195 29461 57207 29495
rect 57149 29455 57207 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 23474 29248 23480 29300
rect 23532 29288 23538 29300
rect 48774 29288 48780 29300
rect 23532 29260 48780 29288
rect 23532 29248 23538 29260
rect 48774 29248 48780 29260
rect 48832 29248 48838 29300
rect 17954 29220 17960 29232
rect 17915 29192 17960 29220
rect 17954 29180 17960 29192
rect 18012 29180 18018 29232
rect 24302 29220 24308 29232
rect 24263 29192 24308 29220
rect 24302 29180 24308 29192
rect 24360 29180 24366 29232
rect 25130 29180 25136 29232
rect 25188 29220 25194 29232
rect 25188 29192 25912 29220
rect 25188 29180 25194 29192
rect 17678 29112 17684 29164
rect 17736 29152 17742 29164
rect 17773 29155 17831 29161
rect 17773 29152 17785 29155
rect 17736 29124 17785 29152
rect 17736 29112 17742 29124
rect 17773 29121 17785 29124
rect 17819 29121 17831 29155
rect 17773 29115 17831 29121
rect 18138 29112 18144 29164
rect 18196 29152 18202 29164
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 18196 29124 18245 29152
rect 18196 29112 18202 29124
rect 18233 29121 18245 29124
rect 18279 29152 18291 29155
rect 20162 29152 20168 29164
rect 18279 29124 20168 29152
rect 18279 29121 18291 29124
rect 18233 29115 18291 29121
rect 20162 29112 20168 29124
rect 20220 29112 20226 29164
rect 23566 29112 23572 29164
rect 23624 29152 23630 29164
rect 24535 29155 24593 29161
rect 24535 29152 24547 29155
rect 23624 29124 24547 29152
rect 23624 29112 23630 29124
rect 24535 29121 24547 29124
rect 24581 29121 24593 29155
rect 25590 29152 25596 29164
rect 25551 29124 25596 29152
rect 24535 29115 24593 29121
rect 25590 29112 25596 29124
rect 25648 29112 25654 29164
rect 25884 29161 25912 29192
rect 25869 29155 25927 29161
rect 25869 29121 25881 29155
rect 25915 29121 25927 29155
rect 25869 29115 25927 29121
rect 24026 29044 24032 29096
rect 24084 29084 24090 29096
rect 24452 29087 24510 29093
rect 24452 29084 24464 29087
rect 24084 29056 24464 29084
rect 24084 29044 24090 29056
rect 24452 29053 24464 29056
rect 24498 29053 24510 29087
rect 24452 29047 24510 29053
rect 24673 29087 24731 29093
rect 24673 29053 24685 29087
rect 24719 29084 24731 29087
rect 25314 29084 25320 29096
rect 24719 29056 25320 29084
rect 24719 29053 24731 29056
rect 24673 29047 24731 29053
rect 25314 29044 25320 29056
rect 25372 29044 25378 29096
rect 25406 29044 25412 29096
rect 25464 29084 25470 29096
rect 25685 29087 25743 29093
rect 25685 29084 25697 29087
rect 25464 29056 25697 29084
rect 25464 29044 25470 29056
rect 25685 29053 25697 29056
rect 25731 29053 25743 29087
rect 25685 29047 25743 29053
rect 26329 29087 26387 29093
rect 26329 29053 26341 29087
rect 26375 29084 26387 29087
rect 26970 29084 26976 29096
rect 26375 29056 26976 29084
rect 26375 29053 26387 29056
rect 26329 29047 26387 29053
rect 26970 29044 26976 29056
rect 27028 29044 27034 29096
rect 24765 29019 24823 29025
rect 24765 29016 24777 29019
rect 24504 28988 24777 29016
rect 24504 28960 24532 28988
rect 24765 28985 24777 28988
rect 24811 28985 24823 29019
rect 24765 28979 24823 28985
rect 24486 28908 24492 28960
rect 24544 28908 24550 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 50982 28500 50988 28552
rect 51040 28540 51046 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 51040 28512 57897 28540
rect 51040 28500 51046 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 18322 28432 18328 28484
rect 18380 28472 18386 28484
rect 39482 28472 39488 28484
rect 18380 28444 39488 28472
rect 18380 28432 18386 28444
rect 39482 28432 39488 28444
rect 39540 28432 39546 28484
rect 58158 28472 58164 28484
rect 58119 28444 58164 28472
rect 58158 28432 58164 28444
rect 58216 28432 58222 28484
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 20162 28404 20168 28416
rect 7708 28376 20168 28404
rect 7708 28364 7714 28376
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 24578 28364 24584 28416
rect 24636 28404 24642 28416
rect 54754 28404 54760 28416
rect 24636 28376 54760 28404
rect 24636 28364 24642 28376
rect 54754 28364 54760 28376
rect 54812 28364 54818 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1578 28160 1584 28212
rect 1636 28200 1642 28212
rect 2869 28203 2927 28209
rect 2869 28200 2881 28203
rect 1636 28172 2881 28200
rect 1636 28160 1642 28172
rect 2869 28169 2881 28172
rect 2915 28169 2927 28203
rect 2869 28163 2927 28169
rect 1581 28067 1639 28073
rect 1581 28033 1593 28067
rect 1627 28033 1639 28067
rect 2498 28064 2504 28076
rect 2459 28036 2504 28064
rect 1581 28027 1639 28033
rect 1596 27928 1624 28027
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2655 28067 2713 28073
rect 2655 28033 2667 28067
rect 2701 28064 2713 28067
rect 4982 28064 4988 28076
rect 2701 28036 4988 28064
rect 2701 28033 2713 28036
rect 2655 28027 2713 28033
rect 4982 28024 4988 28036
rect 5040 28024 5046 28076
rect 58066 28064 58072 28076
rect 58027 28036 58072 28064
rect 58066 28024 58072 28036
rect 58124 28024 58130 28076
rect 1762 27996 1768 28008
rect 1723 27968 1768 27996
rect 1762 27956 1768 27968
rect 1820 27956 1826 28008
rect 14458 27928 14464 27940
rect 1596 27900 2774 27928
rect 2746 27860 2774 27900
rect 12406 27900 14464 27928
rect 12406 27860 12434 27900
rect 14458 27888 14464 27900
rect 14516 27888 14522 27940
rect 2746 27832 12434 27860
rect 32766 27820 32772 27872
rect 32824 27860 32830 27872
rect 58253 27863 58311 27869
rect 58253 27860 58265 27863
rect 32824 27832 58265 27860
rect 32824 27820 32830 27832
rect 58253 27829 58265 27832
rect 58299 27829 58311 27863
rect 58253 27823 58311 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 1854 27384 1860 27396
rect 1815 27356 1860 27384
rect 1854 27344 1860 27356
rect 1912 27344 1918 27396
rect 3234 27344 3240 27396
rect 3292 27384 3298 27396
rect 9582 27384 9588 27396
rect 3292 27356 9588 27384
rect 3292 27344 3298 27356
rect 9582 27344 9588 27356
rect 9640 27344 9646 27396
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 25406 27316 25412 27328
rect 24176 27288 25412 27316
rect 24176 27276 24182 27288
rect 25406 27276 25412 27288
rect 25464 27276 25470 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1578 27072 1584 27124
rect 1636 27112 1642 27124
rect 2869 27115 2927 27121
rect 2869 27112 2881 27115
rect 1636 27084 2881 27112
rect 1636 27072 1642 27084
rect 2869 27081 2881 27084
rect 2915 27081 2927 27115
rect 2869 27075 2927 27081
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26945 1639 26979
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 1581 26939 1639 26945
rect 1596 26840 1624 26939
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2682 26985 2688 26988
rect 2655 26979 2688 26985
rect 2655 26945 2667 26979
rect 2655 26939 2688 26945
rect 2682 26936 2688 26939
rect 2740 26936 2746 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 29546 26976 29552 26988
rect 18104 26948 29552 26976
rect 18104 26936 18110 26948
rect 29546 26936 29552 26948
rect 29604 26936 29610 26988
rect 1762 26908 1768 26920
rect 1723 26880 1768 26908
rect 1762 26868 1768 26880
rect 1820 26868 1826 26920
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 20990 26908 20996 26920
rect 6236 26880 20996 26908
rect 6236 26868 6242 26880
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 23290 26868 23296 26920
rect 23348 26908 23354 26920
rect 55674 26908 55680 26920
rect 23348 26880 55680 26908
rect 23348 26868 23354 26880
rect 55674 26868 55680 26880
rect 55732 26868 55738 26920
rect 15194 26840 15200 26852
rect 1596 26812 2774 26840
rect 2746 26772 2774 26812
rect 12406 26812 15200 26840
rect 12406 26772 12434 26812
rect 15194 26800 15200 26812
rect 15252 26800 15258 26852
rect 2746 26744 12434 26772
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 58158 26432 58164 26444
rect 58119 26404 58164 26432
rect 58158 26392 58164 26404
rect 58216 26392 58222 26444
rect 45646 26324 45652 26376
rect 45704 26364 45710 26376
rect 57885 26367 57943 26373
rect 57885 26364 57897 26367
rect 45704 26336 57897 26364
rect 45704 26324 45710 26336
rect 57885 26333 57897 26336
rect 57931 26333 57943 26367
rect 57885 26327 57943 26333
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 57054 26296 57060 26308
rect 26384 26268 56916 26296
rect 57015 26268 57060 26296
rect 26384 26256 26390 26268
rect 56888 26234 56916 26268
rect 57054 26256 57060 26268
rect 57112 26256 57118 26308
rect 56888 26228 57008 26234
rect 57149 26231 57207 26237
rect 57149 26228 57161 26231
rect 56888 26206 57161 26228
rect 56980 26200 57161 26206
rect 57149 26197 57161 26200
rect 57195 26197 57207 26231
rect 57149 26191 57207 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 18141 25959 18199 25965
rect 18141 25956 18153 25959
rect 2746 25928 18153 25956
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 2746 25888 2774 25928
rect 18141 25925 18153 25928
rect 18187 25925 18199 25959
rect 18141 25919 18199 25925
rect 1627 25860 2774 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 17957 25891 18015 25897
rect 17957 25888 17969 25891
rect 17736 25860 17969 25888
rect 17736 25848 17742 25860
rect 17957 25857 17969 25860
rect 18003 25857 18015 25891
rect 17957 25851 18015 25857
rect 20438 25848 20444 25900
rect 20496 25888 20502 25900
rect 32490 25888 32496 25900
rect 20496 25860 32496 25888
rect 20496 25848 20502 25860
rect 32490 25848 32496 25860
rect 32548 25848 32554 25900
rect 1762 25820 1768 25832
rect 1723 25792 1768 25820
rect 1762 25780 1768 25792
rect 1820 25780 1826 25832
rect 18233 25823 18291 25829
rect 18233 25789 18245 25823
rect 18279 25820 18291 25823
rect 21818 25820 21824 25832
rect 18279 25792 21824 25820
rect 18279 25789 18291 25792
rect 18233 25783 18291 25789
rect 21818 25780 21824 25792
rect 21876 25780 21882 25832
rect 29822 25712 29828 25764
rect 29880 25752 29886 25764
rect 42426 25752 42432 25764
rect 29880 25724 42432 25752
rect 29880 25712 29886 25724
rect 42426 25712 42432 25724
rect 42484 25712 42490 25764
rect 5166 25644 5172 25696
rect 5224 25684 5230 25696
rect 18506 25684 18512 25696
rect 5224 25656 18512 25684
rect 5224 25644 5230 25656
rect 18506 25644 18512 25656
rect 18564 25644 18570 25696
rect 26142 25644 26148 25696
rect 26200 25684 26206 25696
rect 43530 25684 43536 25696
rect 26200 25656 43536 25684
rect 26200 25644 26206 25656
rect 43530 25644 43536 25656
rect 43588 25644 43594 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 2869 25347 2927 25353
rect 2869 25344 2881 25347
rect 1596 25316 2881 25344
rect 1596 25285 1624 25316
rect 2869 25313 2881 25316
rect 2915 25313 2927 25347
rect 2869 25307 2927 25313
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25245 1639 25279
rect 2498 25276 2504 25288
rect 2459 25248 2504 25276
rect 1581 25239 1639 25245
rect 2498 25236 2504 25248
rect 2556 25236 2562 25288
rect 2682 25285 2688 25288
rect 2655 25279 2688 25285
rect 2655 25245 2667 25279
rect 2655 25239 2688 25245
rect 2682 25236 2688 25239
rect 2740 25236 2746 25288
rect 39942 25236 39948 25288
rect 40000 25276 40006 25288
rect 57885 25279 57943 25285
rect 57885 25276 57897 25279
rect 40000 25248 57897 25276
rect 40000 25236 40006 25248
rect 57885 25245 57897 25248
rect 57931 25245 57943 25279
rect 57885 25239 57943 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 58158 25208 58164 25220
rect 58119 25180 58164 25208
rect 58158 25168 58164 25180
rect 58216 25168 58222 25220
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 46750 24828 46756 24880
rect 46808 24868 46814 24880
rect 49050 24868 49056 24880
rect 46808 24840 49056 24868
rect 46808 24828 46814 24840
rect 49050 24828 49056 24840
rect 49108 24828 49114 24880
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 58066 24800 58072 24812
rect 58027 24772 58072 24800
rect 58066 24760 58072 24772
rect 58124 24760 58130 24812
rect 1762 24732 1768 24744
rect 1723 24704 1768 24732
rect 1762 24692 1768 24704
rect 1820 24692 1826 24744
rect 2682 24692 2688 24744
rect 2740 24732 2746 24744
rect 18690 24732 18696 24744
rect 2740 24704 18696 24732
rect 2740 24692 2746 24704
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 37918 24556 37924 24608
rect 37976 24596 37982 24608
rect 58253 24599 58311 24605
rect 58253 24596 58265 24599
rect 37976 24568 58265 24596
rect 37976 24556 37982 24568
rect 58253 24565 58265 24568
rect 58299 24565 58311 24599
rect 58253 24559 58311 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1578 24352 1584 24404
rect 1636 24392 1642 24404
rect 4157 24395 4215 24401
rect 4157 24392 4169 24395
rect 1636 24364 4169 24392
rect 1636 24352 1642 24364
rect 4157 24361 4169 24364
rect 4203 24361 4215 24395
rect 4157 24355 4215 24361
rect 6914 24284 6920 24336
rect 6972 24324 6978 24336
rect 6972 24296 12434 24324
rect 6972 24284 6978 24296
rect 12406 24256 12434 24296
rect 40770 24284 40776 24336
rect 40828 24324 40834 24336
rect 50154 24324 50160 24336
rect 40828 24296 50160 24324
rect 40828 24284 40834 24296
rect 50154 24284 50160 24296
rect 50212 24284 50218 24336
rect 18414 24256 18420 24268
rect 1596 24228 7052 24256
rect 12406 24228 18420 24256
rect 1596 24197 1624 24228
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 1581 24151 1639 24157
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4127 24191 4185 24197
rect 4127 24157 4139 24191
rect 4173 24188 4185 24191
rect 6914 24188 6920 24200
rect 4173 24160 6920 24188
rect 4173 24157 4185 24160
rect 4127 24151 4185 24157
rect 1854 24120 1860 24132
rect 1815 24092 1860 24120
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 3988 24052 4016 24151
rect 6914 24148 6920 24160
rect 6972 24148 6978 24200
rect 7024 24120 7052 24228
rect 18414 24216 18420 24228
rect 18472 24216 18478 24268
rect 24946 24216 24952 24268
rect 25004 24256 25010 24268
rect 47578 24256 47584 24268
rect 25004 24228 47584 24256
rect 25004 24216 25010 24228
rect 47578 24216 47584 24228
rect 47636 24216 47642 24268
rect 17218 24188 17224 24200
rect 12406 24160 17224 24188
rect 12406 24120 12434 24160
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 54018 24188 54024 24200
rect 20036 24160 54024 24188
rect 20036 24148 20042 24160
rect 54018 24148 54024 24160
rect 54076 24148 54082 24200
rect 16850 24120 16856 24132
rect 7024 24092 12434 24120
rect 16546 24092 16856 24120
rect 16546 24052 16574 24092
rect 16850 24080 16856 24092
rect 16908 24080 16914 24132
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 55214 24120 55220 24132
rect 20312 24092 55220 24120
rect 20312 24080 20318 24092
rect 55214 24080 55220 24092
rect 55272 24080 55278 24132
rect 3988 24024 16574 24052
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 17218 23848 17224 23860
rect 17179 23820 17224 23848
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 16850 23712 16856 23724
rect 16763 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 17007 23715 17065 23721
rect 17007 23681 17019 23715
rect 17053 23712 17065 23715
rect 18966 23712 18972 23724
rect 17053 23684 18972 23712
rect 17053 23681 17065 23684
rect 17007 23675 17065 23681
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 16868 23644 16896 23672
rect 17678 23644 17684 23656
rect 16868 23616 17684 23644
rect 17678 23604 17684 23616
rect 17736 23604 17742 23656
rect 15194 23536 15200 23588
rect 15252 23576 15258 23588
rect 18322 23576 18328 23588
rect 15252 23548 18328 23576
rect 15252 23536 15258 23548
rect 18322 23536 18328 23548
rect 18380 23536 18386 23588
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 20530 23508 20536 23520
rect 18472 23480 20536 23508
rect 18472 23468 18478 23480
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 22278 23264 22284 23316
rect 22336 23304 22342 23316
rect 26789 23307 26847 23313
rect 26789 23304 26801 23307
rect 22336 23276 26801 23304
rect 22336 23264 22342 23276
rect 26789 23273 26801 23276
rect 26835 23273 26847 23307
rect 26789 23267 26847 23273
rect 41138 23264 41144 23316
rect 41196 23304 41202 23316
rect 46474 23304 46480 23316
rect 41196 23276 46480 23304
rect 41196 23264 41202 23276
rect 46474 23264 46480 23276
rect 46532 23264 46538 23316
rect 23014 23196 23020 23248
rect 23072 23236 23078 23248
rect 23290 23236 23296 23248
rect 23072 23208 23296 23236
rect 23072 23196 23078 23208
rect 23290 23196 23296 23208
rect 23348 23196 23354 23248
rect 23385 23239 23443 23245
rect 23385 23205 23397 23239
rect 23431 23236 23443 23239
rect 24394 23236 24400 23248
rect 23431 23208 24400 23236
rect 23431 23205 23443 23208
rect 23385 23199 23443 23205
rect 24394 23196 24400 23208
rect 24452 23196 24458 23248
rect 18509 23171 18567 23177
rect 18509 23168 18521 23171
rect 2746 23140 18521 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 2746 23100 2774 23140
rect 18509 23137 18521 23140
rect 18555 23137 18567 23171
rect 18509 23131 18567 23137
rect 26421 23171 26479 23177
rect 26421 23137 26433 23171
rect 26467 23168 26479 23171
rect 27614 23168 27620 23180
rect 26467 23140 27620 23168
rect 26467 23137 26479 23140
rect 26421 23131 26479 23137
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 58158 23168 58164 23180
rect 58119 23140 58164 23168
rect 58158 23128 58164 23140
rect 58216 23128 58222 23180
rect 1627 23072 2774 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 17678 23060 17684 23112
rect 17736 23100 17742 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17736 23072 18153 23100
rect 17736 23060 17742 23072
rect 18141 23069 18153 23072
rect 18187 23069 18199 23103
rect 18141 23063 18199 23069
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 19334 23100 19340 23112
rect 18647 23072 19340 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 20070 23100 20076 23112
rect 19392 23072 20076 23100
rect 19392 23060 19398 23072
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24670 23100 24676 23112
rect 24627 23072 24676 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 26602 23100 26608 23112
rect 26563 23072 26608 23100
rect 26602 23060 26608 23072
rect 26660 23060 26666 23112
rect 57606 23060 57612 23112
rect 57664 23100 57670 23112
rect 57885 23103 57943 23109
rect 57885 23100 57897 23103
rect 57664 23072 57897 23100
rect 57664 23060 57670 23072
rect 57885 23069 57897 23072
rect 57931 23069 57943 23103
rect 57885 23063 57943 23069
rect 1854 23032 1860 23044
rect 1815 23004 1860 23032
rect 1854 22992 1860 23004
rect 1912 22992 1918 23044
rect 22462 22992 22468 23044
rect 22520 23032 22526 23044
rect 23017 23035 23075 23041
rect 23017 23032 23029 23035
rect 22520 23004 23029 23032
rect 22520 22992 22526 23004
rect 23017 23001 23029 23004
rect 23063 23001 23075 23035
rect 23017 22995 23075 23001
rect 24848 23035 24906 23041
rect 24848 23001 24860 23035
rect 24894 23032 24906 23035
rect 25498 23032 25504 23044
rect 24894 23004 25504 23032
rect 24894 23001 24906 23004
rect 24848 22995 24906 23001
rect 25498 22992 25504 23004
rect 25556 22992 25562 23044
rect 25976 23004 31754 23032
rect 23477 22967 23535 22973
rect 23477 22933 23489 22967
rect 23523 22964 23535 22967
rect 24578 22964 24584 22976
rect 23523 22936 24584 22964
rect 23523 22933 23535 22936
rect 23477 22927 23535 22933
rect 24578 22924 24584 22936
rect 24636 22924 24642 22976
rect 25976 22973 26004 23004
rect 25961 22967 26019 22973
rect 25961 22933 25973 22967
rect 26007 22933 26019 22967
rect 31726 22964 31754 23004
rect 32582 22964 32588 22976
rect 31726 22936 32588 22964
rect 25961 22927 26019 22933
rect 32582 22924 32588 22936
rect 32640 22924 32646 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 30650 22720 30656 22772
rect 30708 22760 30714 22772
rect 42518 22760 42524 22772
rect 30708 22732 42524 22760
rect 30708 22720 30714 22732
rect 42518 22720 42524 22732
rect 42576 22720 42582 22772
rect 17681 22695 17739 22701
rect 17681 22692 17693 22695
rect 2746 22664 17693 22692
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 2746 22624 2774 22664
rect 17681 22661 17693 22664
rect 17727 22661 17739 22695
rect 17681 22655 17739 22661
rect 25593 22695 25651 22701
rect 25593 22661 25605 22695
rect 25639 22692 25651 22695
rect 27798 22692 27804 22704
rect 25639 22664 27804 22692
rect 25639 22661 25651 22664
rect 25593 22655 25651 22661
rect 27798 22652 27804 22664
rect 27856 22652 27862 22704
rect 1627 22596 2774 22624
rect 17497 22627 17555 22633
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 17497 22593 17509 22627
rect 17543 22624 17555 22627
rect 22830 22624 22836 22636
rect 17543 22596 17724 22624
rect 22791 22596 22836 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 17696 22568 17724 22596
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 25774 22584 25780 22636
rect 25832 22624 25838 22636
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 25832 22596 27353 22624
rect 25832 22584 25838 22596
rect 27341 22593 27353 22596
rect 27387 22593 27399 22627
rect 58066 22624 58072 22636
rect 58027 22596 58072 22624
rect 27341 22587 27399 22593
rect 58066 22584 58072 22596
rect 58124 22584 58130 22636
rect 1762 22556 1768 22568
rect 1723 22528 1768 22556
rect 1762 22516 1768 22528
rect 1820 22516 1826 22568
rect 17678 22516 17684 22568
rect 17736 22516 17742 22568
rect 17773 22559 17831 22565
rect 17773 22525 17785 22559
rect 17819 22556 17831 22559
rect 23290 22556 23296 22568
rect 17819 22528 23296 22556
rect 17819 22525 17831 22528
rect 17773 22519 17831 22525
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 27157 22559 27215 22565
rect 27157 22525 27169 22559
rect 27203 22556 27215 22559
rect 27614 22556 27620 22568
rect 27203 22528 27620 22556
rect 27203 22525 27215 22528
rect 27157 22519 27215 22525
rect 27614 22516 27620 22528
rect 27672 22556 27678 22568
rect 28442 22556 28448 22568
rect 27672 22528 28448 22556
rect 27672 22516 27678 22528
rect 28442 22516 28448 22528
rect 28500 22516 28506 22568
rect 25866 22488 25872 22500
rect 25827 22460 25872 22488
rect 25866 22448 25872 22460
rect 25924 22448 25930 22500
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 24029 22423 24087 22429
rect 24029 22420 24041 22423
rect 22152 22392 24041 22420
rect 22152 22380 22158 22392
rect 24029 22389 24041 22392
rect 24075 22389 24087 22423
rect 26050 22420 26056 22432
rect 26011 22392 26056 22420
rect 24029 22383 24087 22389
rect 26050 22380 26056 22392
rect 26108 22380 26114 22432
rect 27522 22420 27528 22432
rect 27483 22392 27528 22420
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 32950 22380 32956 22432
rect 33008 22420 33014 22432
rect 34422 22420 34428 22432
rect 33008 22392 34428 22420
rect 33008 22380 33014 22392
rect 34422 22380 34428 22392
rect 34480 22380 34486 22432
rect 38470 22380 38476 22432
rect 38528 22420 38534 22432
rect 58253 22423 58311 22429
rect 58253 22420 58265 22423
rect 38528 22392 58265 22420
rect 38528 22380 38534 22392
rect 58253 22389 58265 22392
rect 58299 22389 58311 22423
rect 58253 22383 58311 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 23566 22176 23572 22228
rect 23624 22216 23630 22228
rect 23937 22219 23995 22225
rect 23937 22216 23949 22219
rect 23624 22188 23949 22216
rect 23624 22176 23630 22188
rect 23937 22185 23949 22188
rect 23983 22185 23995 22219
rect 23937 22179 23995 22185
rect 26510 22176 26516 22228
rect 26568 22216 26574 22228
rect 26568 22188 28580 22216
rect 26568 22176 26574 22188
rect 17681 22151 17739 22157
rect 17681 22148 17693 22151
rect 13832 22120 17693 22148
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 13832 22012 13860 22120
rect 17681 22117 17693 22120
rect 17727 22117 17739 22151
rect 17681 22111 17739 22117
rect 21726 22108 21732 22160
rect 21784 22148 21790 22160
rect 22741 22151 22799 22157
rect 22741 22148 22753 22151
rect 21784 22120 22753 22148
rect 21784 22108 21790 22120
rect 22741 22117 22753 22120
rect 22787 22117 22799 22151
rect 22741 22111 22799 22117
rect 27430 22108 27436 22160
rect 27488 22148 27494 22160
rect 27488 22120 27568 22148
rect 27488 22108 27494 22120
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 17773 22083 17831 22089
rect 17773 22080 17785 22083
rect 16172 22052 17785 22080
rect 16172 22040 16178 22052
rect 17773 22049 17785 22052
rect 17819 22049 17831 22083
rect 22462 22080 22468 22092
rect 22423 22052 22468 22080
rect 17773 22043 17831 22049
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 23753 22083 23811 22089
rect 23753 22049 23765 22083
rect 23799 22080 23811 22083
rect 26418 22080 26424 22092
rect 23799 22052 26424 22080
rect 23799 22049 23811 22052
rect 23753 22043 23811 22049
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 1627 21984 13860 22012
rect 17497 22015 17555 22021
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 17497 21981 17509 22015
rect 17543 22012 17555 22015
rect 17678 22012 17684 22024
rect 17543 21984 17684 22012
rect 17543 21981 17555 21984
rect 17497 21975 17555 21981
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 23661 22015 23719 22021
rect 23661 21981 23673 22015
rect 23707 21981 23719 22015
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 23661 21975 23719 21981
rect 1854 21944 1860 21956
rect 1815 21916 1860 21944
rect 1854 21904 1860 21916
rect 1912 21904 1918 21956
rect 22388 21944 22416 21975
rect 23014 21944 23020 21956
rect 22388 21916 23020 21944
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 23676 21944 23704 21975
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 27341 22015 27399 22021
rect 27341 22014 27353 22015
rect 27264 21986 27353 22014
rect 23750 21944 23756 21956
rect 23676 21916 23756 21944
rect 23750 21904 23756 21916
rect 23808 21904 23814 21956
rect 23934 21904 23940 21956
rect 23992 21944 23998 21956
rect 27264 21944 27292 21986
rect 27341 21981 27353 21986
rect 27387 21981 27399 22015
rect 27341 21975 27399 21981
rect 27540 21953 27568 22120
rect 27709 22015 27767 22021
rect 27709 21981 27721 22015
rect 27755 22012 27767 22015
rect 27890 22012 27896 22024
rect 27755 21984 27896 22012
rect 27755 21981 27767 21984
rect 27709 21975 27767 21981
rect 27890 21972 27896 21984
rect 27948 21972 27954 22024
rect 28442 22012 28448 22024
rect 28403 21984 28448 22012
rect 28442 21972 28448 21984
rect 28500 21972 28506 22024
rect 28552 22021 28580 22188
rect 28537 22015 28595 22021
rect 28537 21981 28549 22015
rect 28583 21981 28595 22015
rect 28537 21975 28595 21981
rect 55858 21972 55864 22024
rect 55916 22012 55922 22024
rect 57885 22015 57943 22021
rect 57885 22012 57897 22015
rect 55916 21984 57897 22012
rect 55916 21972 55922 21984
rect 57885 21981 57897 21984
rect 57931 21981 57943 22015
rect 57885 21975 57943 21981
rect 23992 21916 27292 21944
rect 27525 21947 27583 21953
rect 23992 21904 23998 21916
rect 27525 21913 27537 21947
rect 27571 21913 27583 21947
rect 27525 21907 27583 21913
rect 27617 21947 27675 21953
rect 27617 21913 27629 21947
rect 27663 21913 27675 21947
rect 41322 21944 41328 21956
rect 27617 21907 27675 21913
rect 27908 21916 41328 21944
rect 20346 21836 20352 21888
rect 20404 21876 20410 21888
rect 25777 21879 25835 21885
rect 25777 21876 25789 21879
rect 20404 21848 25789 21876
rect 20404 21836 20410 21848
rect 25777 21845 25789 21848
rect 25823 21845 25835 21879
rect 27632 21876 27660 21907
rect 27706 21876 27712 21888
rect 27632 21848 27712 21876
rect 25777 21839 25835 21845
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 27908 21885 27936 21916
rect 41322 21904 41328 21916
rect 41380 21904 41386 21956
rect 58158 21944 58164 21956
rect 58119 21916 58164 21944
rect 58158 21904 58164 21916
rect 58216 21904 58222 21956
rect 27893 21879 27951 21885
rect 27893 21845 27905 21879
rect 27939 21845 27951 21879
rect 28718 21876 28724 21888
rect 28679 21848 28724 21876
rect 27893 21839 27951 21845
rect 28718 21836 28724 21848
rect 28776 21836 28782 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 22741 21675 22799 21681
rect 22741 21641 22753 21675
rect 22787 21672 22799 21675
rect 22830 21672 22836 21684
rect 22787 21644 22836 21672
rect 22787 21641 22799 21644
rect 22741 21635 22799 21641
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 23293 21675 23351 21681
rect 23293 21641 23305 21675
rect 23339 21641 23351 21675
rect 23293 21635 23351 21641
rect 25685 21675 25743 21681
rect 25685 21641 25697 21675
rect 25731 21672 25743 21675
rect 25866 21672 25872 21684
rect 25731 21644 25872 21672
rect 25731 21641 25743 21644
rect 25685 21635 25743 21641
rect 20898 21604 20904 21616
rect 20859 21576 20904 21604
rect 20898 21564 20904 21576
rect 20956 21564 20962 21616
rect 21174 21613 21180 21616
rect 21117 21607 21180 21613
rect 21117 21573 21129 21607
rect 21163 21573 21180 21607
rect 21117 21567 21180 21573
rect 21174 21564 21180 21567
rect 21232 21564 21238 21616
rect 23308 21604 23336 21635
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 27706 21632 27712 21684
rect 27764 21672 27770 21684
rect 28166 21672 28172 21684
rect 27764 21644 28172 21672
rect 27764 21632 27770 21644
rect 28166 21632 28172 21644
rect 28224 21672 28230 21684
rect 28537 21675 28595 21681
rect 28537 21672 28549 21675
rect 28224 21644 28549 21672
rect 28224 21632 28230 21644
rect 28537 21641 28549 21644
rect 28583 21641 28595 21675
rect 28537 21635 28595 21641
rect 27424 21607 27482 21613
rect 23308 21576 24348 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 8202 21536 8208 21548
rect 1719 21508 8208 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22646 21536 22652 21548
rect 22419 21508 22652 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 23569 21539 23627 21545
rect 23569 21536 23581 21539
rect 23072 21508 23581 21536
rect 23072 21496 23078 21508
rect 23569 21505 23581 21508
rect 23615 21536 23627 21539
rect 24118 21536 24124 21548
rect 23615 21508 24124 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24320 21545 24348 21576
rect 27424 21573 27436 21607
rect 27470 21604 27482 21607
rect 27522 21604 27528 21616
rect 27470 21576 27528 21604
rect 27470 21573 27482 21576
rect 27424 21567 27482 21573
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 25590 21496 25596 21548
rect 25648 21536 25654 21548
rect 28718 21536 28724 21548
rect 25648 21508 28724 21536
rect 25648 21496 25654 21508
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 29178 21536 29184 21548
rect 29139 21508 29184 21536
rect 29178 21496 29184 21508
rect 29236 21496 29242 21548
rect 58066 21536 58072 21548
rect 58027 21508 58072 21536
rect 58066 21496 58072 21508
rect 58124 21496 58130 21548
rect 20622 21428 20628 21480
rect 20680 21468 20686 21480
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 20680 21440 22293 21468
rect 20680 21428 20686 21440
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22281 21431 22339 21437
rect 22462 21428 22468 21480
rect 22520 21468 22526 21480
rect 23106 21468 23112 21480
rect 22520 21440 23112 21468
rect 22520 21428 22526 21440
rect 23106 21428 23112 21440
rect 23164 21468 23170 21480
rect 23477 21471 23535 21477
rect 23477 21468 23489 21471
rect 23164 21440 23489 21468
rect 23164 21428 23170 21440
rect 23477 21437 23489 21440
rect 23523 21437 23535 21471
rect 23477 21431 23535 21437
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23753 21471 23811 21477
rect 23753 21437 23765 21471
rect 23799 21468 23811 21471
rect 26234 21468 26240 21480
rect 23799 21440 26240 21468
rect 23799 21437 23811 21440
rect 23753 21431 23811 21437
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 21082 21332 21088 21344
rect 21043 21304 21088 21332
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 21266 21332 21272 21344
rect 21227 21304 21272 21332
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 23676 21332 23704 21431
rect 26234 21428 26240 21440
rect 26292 21428 26298 21480
rect 27157 21471 27215 21477
rect 27157 21437 27169 21471
rect 27203 21437 27215 21471
rect 27157 21431 27215 21437
rect 23750 21332 23756 21344
rect 23663 21304 23756 21332
rect 23750 21292 23756 21304
rect 23808 21332 23814 21344
rect 26694 21332 26700 21344
rect 23808 21304 26700 21332
rect 23808 21292 23814 21304
rect 26694 21292 26700 21304
rect 26752 21292 26758 21344
rect 27172 21332 27200 21431
rect 28442 21428 28448 21480
rect 28500 21468 28506 21480
rect 28810 21468 28816 21480
rect 28500 21440 28816 21468
rect 28500 21428 28506 21440
rect 28810 21428 28816 21440
rect 28868 21468 28874 21480
rect 28997 21471 29055 21477
rect 28997 21468 29009 21471
rect 28868 21440 29009 21468
rect 28868 21428 28874 21440
rect 28997 21437 29009 21440
rect 29043 21437 29055 21471
rect 28997 21431 29055 21437
rect 28534 21360 28540 21412
rect 28592 21400 28598 21412
rect 28592 21372 31754 21400
rect 28592 21360 28598 21372
rect 28442 21332 28448 21344
rect 27172 21304 28448 21332
rect 28442 21292 28448 21304
rect 28500 21292 28506 21344
rect 28994 21292 29000 21344
rect 29052 21332 29058 21344
rect 29365 21335 29423 21341
rect 29365 21332 29377 21335
rect 29052 21304 29377 21332
rect 29052 21292 29058 21304
rect 29365 21301 29377 21304
rect 29411 21301 29423 21335
rect 31726 21332 31754 21372
rect 40034 21360 40040 21412
rect 40092 21400 40098 21412
rect 42058 21400 42064 21412
rect 40092 21372 42064 21400
rect 40092 21360 40098 21372
rect 42058 21360 42064 21372
rect 42116 21360 42122 21412
rect 58253 21335 58311 21341
rect 58253 21332 58265 21335
rect 31726 21304 58265 21332
rect 29365 21295 29423 21301
rect 58253 21301 58265 21304
rect 58299 21301 58311 21335
rect 58253 21295 58311 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 21085 21131 21143 21137
rect 21085 21097 21097 21131
rect 21131 21128 21143 21131
rect 22002 21128 22008 21140
rect 21131 21100 22008 21128
rect 21131 21097 21143 21100
rect 21085 21091 21143 21097
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 27338 21088 27344 21140
rect 27396 21128 27402 21140
rect 29733 21131 29791 21137
rect 29733 21128 29745 21131
rect 27396 21100 29745 21128
rect 27396 21088 27402 21100
rect 29733 21097 29745 21100
rect 29779 21097 29791 21131
rect 29733 21091 29791 21097
rect 19242 21020 19248 21072
rect 19300 21060 19306 21072
rect 21269 21063 21327 21069
rect 21269 21060 21281 21063
rect 19300 21032 21281 21060
rect 19300 21020 19306 21032
rect 21269 21029 21281 21032
rect 21315 21060 21327 21063
rect 27154 21060 27160 21072
rect 21315 21032 27160 21060
rect 21315 21029 21327 21032
rect 21269 21023 21327 21029
rect 27154 21020 27160 21032
rect 27212 21020 27218 21072
rect 23382 20952 23388 21004
rect 23440 20992 23446 21004
rect 24670 20992 24676 21004
rect 23440 20964 24676 20992
rect 23440 20952 23446 20964
rect 24670 20952 24676 20964
rect 24728 20992 24734 21004
rect 27525 20995 27583 21001
rect 27525 20992 27537 20995
rect 24728 20964 27537 20992
rect 24728 20952 24734 20964
rect 27525 20961 27537 20964
rect 27571 20961 27583 20995
rect 27525 20955 27583 20961
rect 28902 20952 28908 21004
rect 28960 20992 28966 21004
rect 30285 20995 30343 21001
rect 30285 20992 30297 20995
rect 28960 20964 30297 20992
rect 28960 20952 28966 20964
rect 30285 20961 30297 20964
rect 30331 20961 30343 20995
rect 30285 20955 30343 20961
rect 20070 20924 20076 20936
rect 20031 20896 20076 20924
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20924 20315 20927
rect 21266 20924 21272 20936
rect 20303 20896 21272 20924
rect 20303 20893 20315 20896
rect 20257 20887 20315 20893
rect 16666 20816 16672 20868
rect 16724 20856 16730 20868
rect 20272 20856 20300 20887
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 21729 20927 21787 20933
rect 21729 20893 21741 20927
rect 21775 20924 21787 20927
rect 22094 20924 22100 20936
rect 21775 20896 22100 20924
rect 21775 20893 21787 20896
rect 21729 20887 21787 20893
rect 22094 20884 22100 20896
rect 22152 20884 22158 20936
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 26050 20924 26056 20936
rect 24811 20896 26056 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 45094 20884 45100 20936
rect 45152 20924 45158 20936
rect 46014 20924 46020 20936
rect 45152 20896 46020 20924
rect 45152 20884 45158 20896
rect 46014 20884 46020 20896
rect 46072 20884 46078 20936
rect 16724 20828 20300 20856
rect 16724 20816 16730 20828
rect 20714 20816 20720 20868
rect 20772 20856 20778 20868
rect 20901 20859 20959 20865
rect 20901 20856 20913 20859
rect 20772 20828 20913 20856
rect 20772 20816 20778 20828
rect 20901 20825 20913 20828
rect 20947 20825 20959 20859
rect 20901 20819 20959 20825
rect 27065 20859 27123 20865
rect 27065 20825 27077 20859
rect 27111 20856 27123 20859
rect 27770 20859 27828 20865
rect 27770 20856 27782 20859
rect 27111 20828 27782 20856
rect 27111 20825 27123 20828
rect 27065 20819 27123 20825
rect 27770 20825 27782 20828
rect 27816 20825 27828 20859
rect 27770 20819 27828 20825
rect 32398 20816 32404 20868
rect 32456 20856 32462 20868
rect 33778 20856 33784 20868
rect 32456 20828 33784 20856
rect 32456 20816 32462 20828
rect 33778 20816 33784 20828
rect 33836 20816 33842 20868
rect 44266 20816 44272 20868
rect 44324 20856 44330 20868
rect 47762 20856 47768 20868
rect 44324 20828 47768 20856
rect 44324 20816 44330 20828
rect 47762 20816 47768 20828
rect 47820 20816 47826 20868
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 20530 20788 20536 20800
rect 20487 20760 20536 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21101 20791 21159 20797
rect 21101 20788 21113 20791
rect 20864 20760 21113 20788
rect 20864 20748 20870 20760
rect 21101 20757 21113 20760
rect 21147 20788 21159 20791
rect 21266 20788 21272 20800
rect 21147 20760 21272 20788
rect 21147 20757 21159 20760
rect 21101 20751 21159 20757
rect 21266 20748 21272 20760
rect 21324 20748 21330 20800
rect 22922 20788 22928 20800
rect 22883 20760 22928 20788
rect 22922 20748 22928 20760
rect 22980 20748 22986 20800
rect 27246 20748 27252 20800
rect 27304 20788 27310 20800
rect 27890 20788 27896 20800
rect 27304 20760 27896 20788
rect 27304 20748 27310 20760
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 28258 20748 28264 20800
rect 28316 20788 28322 20800
rect 28905 20791 28963 20797
rect 28905 20788 28917 20791
rect 28316 20760 28917 20788
rect 28316 20748 28322 20760
rect 28905 20757 28917 20760
rect 28951 20757 28963 20791
rect 30098 20788 30104 20800
rect 30059 20760 30104 20788
rect 28905 20751 28963 20757
rect 30098 20748 30104 20760
rect 30156 20748 30162 20800
rect 30193 20791 30251 20797
rect 30193 20757 30205 20791
rect 30239 20788 30251 20791
rect 30837 20791 30895 20797
rect 30837 20788 30849 20791
rect 30239 20760 30849 20788
rect 30239 20757 30251 20760
rect 30193 20751 30251 20757
rect 30837 20757 30849 20760
rect 30883 20788 30895 20791
rect 31386 20788 31392 20800
rect 30883 20760 31392 20788
rect 30883 20757 30895 20760
rect 30837 20751 30895 20757
rect 31386 20748 31392 20760
rect 31444 20788 31450 20800
rect 58342 20788 58348 20800
rect 31444 20760 58348 20788
rect 31444 20748 31450 20760
rect 58342 20748 58348 20760
rect 58400 20748 58406 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 19521 20587 19579 20593
rect 19521 20553 19533 20587
rect 19567 20584 19579 20587
rect 20622 20584 20628 20596
rect 19567 20556 20628 20584
rect 19567 20553 19579 20556
rect 19521 20547 19579 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20772 20556 21128 20584
rect 20772 20544 20778 20556
rect 19978 20516 19984 20528
rect 19352 20488 19984 20516
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 14274 20448 14280 20460
rect 1627 20420 14280 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18782 20448 18788 20460
rect 18739 20420 18788 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 19352 20457 19380 20488
rect 19978 20476 19984 20488
rect 20036 20516 20042 20528
rect 20036 20488 21036 20516
rect 20036 20476 20042 20488
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20417 19395 20451
rect 19518 20448 19524 20460
rect 19479 20420 19524 20448
rect 19337 20411 19395 20417
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 18892 20312 18920 20411
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 20254 20457 20260 20460
rect 20248 20448 20260 20457
rect 20215 20420 20260 20448
rect 20248 20411 20260 20420
rect 20254 20408 20260 20411
rect 20312 20408 20318 20460
rect 19426 20340 19432 20392
rect 19484 20380 19490 20392
rect 19981 20383 20039 20389
rect 19981 20380 19993 20383
rect 19484 20352 19993 20380
rect 19484 20340 19490 20352
rect 19981 20349 19993 20352
rect 20027 20349 20039 20383
rect 21008 20380 21036 20488
rect 21100 20448 21128 20556
rect 21266 20544 21272 20596
rect 21324 20584 21330 20596
rect 22833 20587 22891 20593
rect 22833 20584 22845 20587
rect 21324 20556 22845 20584
rect 21324 20544 21330 20556
rect 22833 20553 22845 20556
rect 22879 20553 22891 20587
rect 26418 20584 26424 20596
rect 26379 20556 26424 20584
rect 22833 20547 22891 20553
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 27433 20587 27491 20593
rect 27433 20553 27445 20587
rect 27479 20584 27491 20587
rect 33502 20584 33508 20596
rect 27479 20556 33508 20584
rect 27479 20553 27491 20556
rect 27433 20547 27491 20553
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 22152 20488 22753 20516
rect 22152 20476 22158 20488
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 24118 20476 24124 20528
rect 24176 20516 24182 20528
rect 27448 20516 27476 20547
rect 33502 20544 33508 20556
rect 33560 20544 33566 20596
rect 29730 20516 29736 20528
rect 24176 20488 27476 20516
rect 28460 20488 29736 20516
rect 24176 20476 24182 20488
rect 21910 20448 21916 20460
rect 21100 20420 21916 20448
rect 21910 20408 21916 20420
rect 21968 20448 21974 20460
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 21968 20420 22661 20448
rect 21968 20408 21974 20420
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 23566 20448 23572 20460
rect 23527 20420 23572 20448
rect 22649 20411 22707 20417
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 26528 20457 26556 20488
rect 28460 20460 28488 20488
rect 29730 20476 29736 20488
rect 29788 20516 29794 20528
rect 29788 20488 30420 20516
rect 29788 20476 29794 20488
rect 26329 20451 26387 20457
rect 26329 20448 26341 20451
rect 24636 20420 26341 20448
rect 24636 20408 24642 20420
rect 26329 20417 26341 20420
rect 26375 20417 26387 20451
rect 26329 20411 26387 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20417 26571 20451
rect 26513 20411 26571 20417
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 21008 20352 23029 20380
rect 19981 20343 20039 20349
rect 23017 20349 23029 20352
rect 23063 20380 23075 20383
rect 23474 20380 23480 20392
rect 23063 20352 23480 20380
rect 23063 20349 23075 20352
rect 23017 20343 23075 20349
rect 23474 20340 23480 20352
rect 23532 20380 23538 20392
rect 25130 20380 25136 20392
rect 23532 20352 25136 20380
rect 23532 20340 23538 20352
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 26344 20380 26372 20411
rect 26694 20408 26700 20460
rect 26752 20448 26758 20460
rect 27341 20451 27399 20457
rect 27341 20448 27353 20451
rect 26752 20420 27353 20448
rect 26752 20408 26758 20420
rect 27341 20417 27353 20420
rect 27387 20448 27399 20451
rect 27430 20448 27436 20460
rect 27387 20420 27436 20448
rect 27387 20417 27399 20420
rect 27341 20411 27399 20417
rect 27430 20408 27436 20420
rect 27488 20408 27494 20460
rect 27525 20451 27583 20457
rect 27525 20417 27537 20451
rect 27571 20417 27583 20451
rect 28442 20448 28448 20460
rect 28403 20420 28448 20448
rect 27525 20411 27583 20417
rect 27540 20380 27568 20411
rect 28442 20408 28448 20420
rect 28500 20408 28506 20460
rect 28712 20451 28770 20457
rect 28712 20417 28724 20451
rect 28758 20448 28770 20451
rect 28994 20448 29000 20460
rect 28758 20420 29000 20448
rect 28758 20417 28770 20420
rect 28712 20411 28770 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 30392 20457 30420 20488
rect 30484 20488 31754 20516
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 30484 20380 30512 20488
rect 30650 20457 30656 20460
rect 30633 20451 30656 20457
rect 30633 20417 30645 20451
rect 30633 20411 30656 20417
rect 30650 20408 30656 20411
rect 30708 20408 30714 20460
rect 31726 20448 31754 20488
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 31726 20420 32321 20448
rect 32309 20417 32321 20420
rect 32355 20417 32367 20451
rect 32490 20448 32496 20460
rect 32451 20420 32496 20448
rect 32309 20411 32367 20417
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 38746 20448 38752 20460
rect 38707 20420 38752 20448
rect 38746 20408 38752 20420
rect 38804 20408 38810 20460
rect 26344 20352 27568 20380
rect 29656 20352 30512 20380
rect 18966 20312 18972 20324
rect 18879 20284 18972 20312
rect 18966 20272 18972 20284
rect 19024 20312 19030 20324
rect 19886 20312 19892 20324
rect 19024 20284 19892 20312
rect 19024 20272 19030 20284
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 22370 20272 22376 20324
rect 22428 20312 22434 20324
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 22428 20284 22477 20312
rect 22428 20272 22434 20284
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 23032 20284 26188 20312
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 16632 20216 18705 20244
rect 16632 20204 16638 20216
rect 18693 20213 18705 20216
rect 18739 20213 18751 20247
rect 18693 20207 18751 20213
rect 19702 20204 19708 20256
rect 19760 20244 19766 20256
rect 20714 20244 20720 20256
rect 19760 20216 20720 20244
rect 19760 20204 19766 20216
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 23032 20244 23060 20284
rect 21407 20216 23060 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 23106 20204 23112 20256
rect 23164 20244 23170 20256
rect 24578 20244 24584 20256
rect 23164 20216 24584 20244
rect 23164 20204 23170 20216
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 24762 20244 24768 20256
rect 24723 20216 24768 20244
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 26160 20244 26188 20284
rect 26234 20272 26240 20324
rect 26292 20312 26298 20324
rect 27157 20315 27215 20321
rect 27157 20312 27169 20315
rect 26292 20284 27169 20312
rect 26292 20272 26298 20284
rect 27157 20281 27169 20284
rect 27203 20312 27215 20315
rect 27890 20312 27896 20324
rect 27203 20284 27896 20312
rect 27203 20281 27215 20284
rect 27157 20275 27215 20281
rect 27890 20272 27896 20284
rect 27948 20272 27954 20324
rect 26878 20244 26884 20256
rect 26160 20216 26884 20244
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 27709 20247 27767 20253
rect 27709 20213 27721 20247
rect 27755 20244 27767 20247
rect 27798 20244 27804 20256
rect 27755 20216 27804 20244
rect 27755 20213 27767 20216
rect 27709 20207 27767 20213
rect 27798 20204 27804 20216
rect 27856 20204 27862 20256
rect 28718 20204 28724 20256
rect 28776 20244 28782 20256
rect 29656 20244 29684 20352
rect 38378 20340 38384 20392
rect 38436 20380 38442 20392
rect 38565 20383 38623 20389
rect 38565 20380 38577 20383
rect 38436 20352 38577 20380
rect 38436 20340 38442 20352
rect 38565 20349 38577 20352
rect 38611 20349 38623 20383
rect 38565 20343 38623 20349
rect 39206 20340 39212 20392
rect 39264 20380 39270 20392
rect 57974 20380 57980 20392
rect 39264 20352 57980 20380
rect 39264 20340 39270 20352
rect 57974 20340 57980 20352
rect 58032 20340 58038 20392
rect 36262 20272 36268 20324
rect 36320 20312 36326 20324
rect 39114 20312 39120 20324
rect 36320 20284 39120 20312
rect 36320 20272 36326 20284
rect 39114 20272 39120 20284
rect 39172 20312 39178 20324
rect 39758 20312 39764 20324
rect 39172 20284 39764 20312
rect 39172 20272 39178 20284
rect 39758 20272 39764 20284
rect 39816 20272 39822 20324
rect 29822 20244 29828 20256
rect 28776 20216 29684 20244
rect 29783 20216 29828 20244
rect 28776 20204 28782 20216
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30098 20204 30104 20256
rect 30156 20244 30162 20256
rect 31757 20247 31815 20253
rect 31757 20244 31769 20247
rect 30156 20216 31769 20244
rect 30156 20204 30162 20216
rect 31757 20213 31769 20216
rect 31803 20213 31815 20247
rect 31757 20207 31815 20213
rect 31846 20204 31852 20256
rect 31904 20244 31910 20256
rect 32677 20247 32735 20253
rect 32677 20244 32689 20247
rect 31904 20216 32689 20244
rect 31904 20204 31910 20216
rect 32677 20213 32689 20216
rect 32723 20213 32735 20247
rect 32677 20207 32735 20213
rect 38933 20247 38991 20253
rect 38933 20213 38945 20247
rect 38979 20244 38991 20247
rect 39022 20244 39028 20256
rect 38979 20216 39028 20244
rect 38979 20213 38991 20216
rect 38933 20207 38991 20213
rect 39022 20204 39028 20216
rect 39080 20204 39086 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 19702 20040 19708 20052
rect 18156 20012 19708 20040
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19836 1639 19839
rect 4062 19836 4068 19848
rect 1627 19808 4068 19836
rect 1627 19805 1639 19808
rect 1581 19799 1639 19805
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 15068 19808 17969 19836
rect 15068 19796 15074 19808
rect 17957 19805 17969 19808
rect 18003 19836 18015 19839
rect 18046 19836 18052 19848
rect 18003 19808 18052 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 18046 19796 18052 19808
rect 18104 19796 18110 19848
rect 18156 19845 18184 20012
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 20898 20040 20904 20052
rect 19812 20012 20904 20040
rect 18598 19972 18604 19984
rect 18559 19944 18604 19972
rect 18598 19932 18604 19944
rect 18656 19932 18662 19984
rect 19812 19904 19840 20012
rect 20898 20000 20904 20012
rect 20956 20040 20962 20052
rect 24118 20040 24124 20052
rect 20956 20012 24124 20040
rect 20956 20000 20962 20012
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 24578 20000 24584 20052
rect 24636 20040 24642 20052
rect 25133 20043 25191 20049
rect 25133 20040 25145 20043
rect 24636 20012 25145 20040
rect 24636 20000 24642 20012
rect 25133 20009 25145 20012
rect 25179 20009 25191 20043
rect 25133 20003 25191 20009
rect 25222 20000 25228 20052
rect 25280 20040 25286 20052
rect 30374 20040 30380 20052
rect 25280 20012 30380 20040
rect 25280 20000 25286 20012
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 38565 20043 38623 20049
rect 30484 20012 31754 20040
rect 21177 19975 21235 19981
rect 21177 19941 21189 19975
rect 21223 19972 21235 19975
rect 29825 19975 29883 19981
rect 21223 19944 28994 19972
rect 21223 19941 21235 19944
rect 21177 19935 21235 19941
rect 18616 19876 19840 19904
rect 24029 19907 24087 19913
rect 18616 19845 18644 19876
rect 24029 19873 24041 19907
rect 24075 19904 24087 19907
rect 24854 19904 24860 19916
rect 24075 19876 24860 19904
rect 24075 19873 24087 19876
rect 24029 19867 24087 19873
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 25130 19904 25136 19916
rect 24964 19876 25136 19904
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 18966 19836 18972 19848
rect 18923 19808 18972 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19426 19796 19432 19848
rect 19484 19836 19490 19848
rect 19797 19839 19855 19845
rect 19797 19836 19809 19839
rect 19484 19808 19809 19836
rect 19484 19796 19490 19808
rect 19797 19805 19809 19808
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 21174 19836 21180 19848
rect 19944 19808 21180 19836
rect 19944 19796 19950 19808
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19836 21787 19839
rect 24670 19836 24676 19848
rect 21775 19808 24676 19836
rect 21775 19805 21787 19808
rect 21729 19799 21787 19805
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 24964 19845 24992 19876
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 27341 19907 27399 19913
rect 27341 19904 27353 19907
rect 25740 19876 27353 19904
rect 25740 19864 25746 19876
rect 27341 19873 27353 19876
rect 27387 19873 27399 19907
rect 28966 19904 28994 19944
rect 29825 19941 29837 19975
rect 29871 19972 29883 19975
rect 30484 19972 30512 20012
rect 29871 19944 30512 19972
rect 31726 19972 31754 20012
rect 38565 20009 38577 20043
rect 38611 20040 38623 20043
rect 38746 20040 38752 20052
rect 38611 20012 38752 20040
rect 38611 20009 38623 20012
rect 38565 20003 38623 20009
rect 38746 20000 38752 20012
rect 38804 20000 38810 20052
rect 40218 20000 40224 20052
rect 40276 20040 40282 20052
rect 41138 20040 41144 20052
rect 40276 20012 41144 20040
rect 40276 20000 40282 20012
rect 41138 20000 41144 20012
rect 41196 20000 41202 20052
rect 48130 20000 48136 20052
rect 48188 20040 48194 20052
rect 48958 20040 48964 20052
rect 48188 20012 48964 20040
rect 48188 20000 48194 20012
rect 48958 20000 48964 20012
rect 49016 20000 49022 20052
rect 47854 19972 47860 19984
rect 31726 19944 47860 19972
rect 29871 19941 29883 19944
rect 29825 19935 29883 19941
rect 47854 19932 47860 19944
rect 47912 19932 47918 19984
rect 28966 19876 30512 19904
rect 27341 19867 27399 19873
rect 24949 19839 25007 19845
rect 24820 19808 24865 19836
rect 24820 19796 24826 19808
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 26050 19796 26056 19848
rect 26108 19836 26114 19848
rect 26237 19839 26295 19845
rect 26237 19836 26249 19839
rect 26108 19808 26249 19836
rect 26108 19796 26114 19808
rect 26237 19805 26249 19808
rect 26283 19836 26295 19839
rect 30098 19836 30104 19848
rect 26283 19808 30104 19836
rect 26283 19805 26295 19808
rect 26237 19799 26295 19805
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 17310 19728 17316 19780
rect 17368 19768 17374 19780
rect 17368 19740 18460 19768
rect 17368 19728 17374 19740
rect 18046 19700 18052 19712
rect 18007 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 18432 19700 18460 19740
rect 18506 19728 18512 19780
rect 18564 19768 18570 19780
rect 20064 19771 20122 19777
rect 18564 19740 19564 19768
rect 18564 19728 18570 19740
rect 19536 19712 19564 19740
rect 20064 19737 20076 19771
rect 20110 19768 20122 19771
rect 22462 19768 22468 19780
rect 20110 19740 22468 19768
rect 20110 19737 20122 19740
rect 20064 19731 20122 19737
rect 22462 19728 22468 19740
rect 22520 19728 22526 19780
rect 24578 19768 24584 19780
rect 24539 19740 24584 19768
rect 24578 19728 24584 19740
rect 24636 19728 24642 19780
rect 30377 19771 30435 19777
rect 30377 19737 30389 19771
rect 30423 19737 30435 19771
rect 30484 19768 30512 19876
rect 30558 19864 30564 19916
rect 30616 19904 30622 19916
rect 32401 19907 32459 19913
rect 32401 19904 32413 19907
rect 30616 19876 32413 19904
rect 30616 19864 30622 19876
rect 32401 19873 32413 19876
rect 32447 19873 32459 19907
rect 32401 19867 32459 19873
rect 39117 19907 39175 19913
rect 39117 19873 39129 19907
rect 39163 19904 39175 19907
rect 39163 19876 39344 19904
rect 39163 19873 39175 19876
rect 39117 19867 39175 19873
rect 31297 19839 31355 19845
rect 31297 19805 31309 19839
rect 31343 19836 31355 19839
rect 33042 19836 33048 19848
rect 31343 19808 33048 19836
rect 31343 19805 31355 19808
rect 31297 19799 31355 19805
rect 33042 19796 33048 19808
rect 33100 19796 33106 19848
rect 36262 19796 36268 19848
rect 36320 19836 36326 19848
rect 36449 19839 36507 19845
rect 36449 19836 36461 19839
rect 36320 19808 36461 19836
rect 36320 19796 36326 19808
rect 36449 19805 36461 19808
rect 36495 19805 36507 19839
rect 36449 19799 36507 19805
rect 36633 19839 36691 19845
rect 36633 19805 36645 19839
rect 36679 19836 36691 19839
rect 37458 19836 37464 19848
rect 36679 19808 37464 19836
rect 36679 19805 36691 19808
rect 36633 19799 36691 19805
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 38289 19839 38347 19845
rect 38289 19805 38301 19839
rect 38335 19836 38347 19839
rect 39025 19839 39083 19845
rect 39025 19836 39037 19839
rect 38335 19808 39037 19836
rect 38335 19805 38347 19808
rect 38289 19799 38347 19805
rect 39025 19805 39037 19808
rect 39071 19836 39083 19839
rect 39206 19836 39212 19848
rect 39071 19808 39212 19836
rect 39071 19805 39083 19808
rect 39025 19799 39083 19805
rect 39206 19796 39212 19808
rect 39264 19796 39270 19848
rect 39316 19836 39344 19876
rect 39758 19864 39764 19916
rect 39816 19904 39822 19916
rect 40497 19907 40555 19913
rect 40497 19904 40509 19907
rect 39816 19876 40509 19904
rect 39816 19864 39822 19876
rect 40497 19873 40509 19876
rect 40543 19873 40555 19907
rect 41414 19904 41420 19916
rect 40497 19867 40555 19873
rect 40604 19876 41420 19904
rect 40310 19836 40316 19848
rect 39316 19808 40316 19836
rect 40310 19796 40316 19808
rect 40368 19836 40374 19848
rect 40604 19836 40632 19876
rect 41414 19864 41420 19876
rect 41472 19864 41478 19916
rect 48133 19907 48191 19913
rect 48133 19873 48145 19907
rect 48179 19904 48191 19907
rect 48866 19904 48872 19916
rect 48179 19876 48872 19904
rect 48179 19873 48191 19876
rect 48133 19867 48191 19873
rect 48866 19864 48872 19876
rect 48924 19864 48930 19916
rect 58158 19904 58164 19916
rect 58119 19876 58164 19904
rect 58158 19864 58164 19876
rect 58216 19864 58222 19916
rect 40368 19808 40632 19836
rect 40701 19839 40759 19845
rect 40368 19796 40374 19808
rect 40701 19805 40713 19839
rect 40747 19836 40759 19839
rect 40862 19836 40868 19848
rect 40747 19808 40868 19836
rect 40747 19805 40759 19808
rect 40701 19799 40759 19805
rect 40862 19796 40868 19808
rect 40920 19796 40926 19848
rect 48317 19839 48375 19845
rect 48317 19805 48329 19839
rect 48363 19836 48375 19839
rect 48590 19836 48596 19848
rect 48363 19808 48596 19836
rect 48363 19805 48375 19808
rect 48317 19799 48375 19805
rect 48590 19796 48596 19808
rect 48648 19796 48654 19848
rect 57885 19839 57943 19845
rect 57885 19836 57897 19839
rect 55186 19808 57897 19836
rect 37366 19768 37372 19780
rect 30484 19740 37372 19768
rect 30377 19731 30435 19737
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18432 19672 18797 19700
rect 18785 19669 18797 19672
rect 18831 19700 18843 19703
rect 19058 19700 19064 19712
rect 18831 19672 19064 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 19058 19660 19064 19672
rect 19116 19660 19122 19712
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 24857 19703 24915 19709
rect 24857 19700 24869 19703
rect 19576 19672 24869 19700
rect 19576 19660 19582 19672
rect 24857 19669 24869 19672
rect 24903 19700 24915 19703
rect 26786 19700 26792 19712
rect 24903 19672 26792 19700
rect 24903 19669 24915 19672
rect 24857 19663 24915 19669
rect 26786 19660 26792 19672
rect 26844 19660 26850 19712
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 28810 19700 28816 19712
rect 27672 19672 28816 19700
rect 27672 19660 27678 19672
rect 28810 19660 28816 19672
rect 28868 19660 28874 19712
rect 30282 19700 30288 19712
rect 30243 19672 30288 19700
rect 30282 19660 30288 19672
rect 30340 19660 30346 19712
rect 30392 19700 30420 19731
rect 37366 19728 37372 19740
rect 37424 19728 37430 19780
rect 37734 19728 37740 19780
rect 37792 19768 37798 19780
rect 55186 19768 55214 19808
rect 57885 19805 57897 19808
rect 57931 19805 57943 19839
rect 57885 19799 57943 19805
rect 37792 19740 55214 19768
rect 37792 19728 37798 19740
rect 30834 19700 30840 19712
rect 30392 19672 30840 19700
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 35526 19660 35532 19712
rect 35584 19700 35590 19712
rect 36446 19700 36452 19712
rect 35584 19672 36452 19700
rect 35584 19660 35590 19672
rect 36446 19660 36452 19672
rect 36504 19660 36510 19712
rect 36814 19700 36820 19712
rect 36775 19672 36820 19700
rect 36814 19660 36820 19672
rect 36872 19660 36878 19712
rect 38838 19660 38844 19712
rect 38896 19700 38902 19712
rect 38933 19703 38991 19709
rect 38933 19700 38945 19703
rect 38896 19672 38945 19700
rect 38896 19660 38902 19672
rect 38933 19669 38945 19672
rect 38979 19669 38991 19703
rect 38933 19663 38991 19669
rect 40770 19660 40776 19712
rect 40828 19700 40834 19712
rect 40865 19703 40923 19709
rect 40865 19700 40877 19703
rect 40828 19672 40877 19700
rect 40828 19660 40834 19672
rect 40865 19669 40877 19672
rect 40911 19669 40923 19703
rect 48498 19700 48504 19712
rect 48459 19672 48504 19700
rect 40865 19663 40923 19669
rect 48498 19660 48504 19672
rect 48556 19660 48562 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 19242 19496 19248 19508
rect 17512 19468 19248 19496
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19329 1639 19363
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1581 19323 1639 19329
rect 1596 19292 1624 19323
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 17512 19369 17540 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 20349 19499 20407 19505
rect 20349 19496 20361 19499
rect 20312 19468 20361 19496
rect 20312 19456 20318 19468
rect 20349 19465 20361 19468
rect 20395 19465 20407 19499
rect 23750 19496 23756 19508
rect 20349 19459 20407 19465
rect 21928 19468 22232 19496
rect 23711 19468 23756 19496
rect 21928 19428 21956 19468
rect 17696 19400 21956 19428
rect 17696 19369 17724 19400
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18506 19360 18512 19372
rect 18371 19332 18512 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 18708 19332 19165 19360
rect 18708 19301 18736 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 21082 19360 21088 19372
rect 19153 19323 19211 19329
rect 19260 19332 21088 19360
rect 18417 19295 18475 19301
rect 1596 19264 2452 19292
rect 2424 19165 2452 19264
rect 18417 19261 18429 19295
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 18432 19224 18460 19255
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19260 19292 19288 19332
rect 21082 19320 21088 19332
rect 21140 19360 21146 19372
rect 21450 19360 21456 19372
rect 21140 19332 21456 19360
rect 21140 19320 21146 19332
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 21836 19360 21956 19363
rect 21692 19335 22094 19360
rect 21692 19332 21864 19335
rect 21928 19332 22094 19335
rect 21692 19320 21698 19332
rect 19116 19264 19288 19292
rect 19116 19252 19122 19264
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 22066 19292 22094 19332
rect 19484 19264 22094 19292
rect 22204 19292 22232 19468
rect 23750 19456 23756 19468
rect 23808 19456 23814 19508
rect 25498 19496 25504 19508
rect 25459 19468 25504 19496
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 27249 19499 27307 19505
rect 27249 19465 27261 19499
rect 27295 19496 27307 19499
rect 27706 19496 27712 19508
rect 27295 19468 27712 19496
rect 27295 19465 27307 19468
rect 27249 19459 27307 19465
rect 27706 19456 27712 19468
rect 27764 19456 27770 19508
rect 30009 19499 30067 19505
rect 30009 19496 30021 19499
rect 27816 19468 30021 19496
rect 22738 19428 22744 19440
rect 22388 19400 22744 19428
rect 22388 19369 22416 19400
rect 22738 19388 22744 19400
rect 22796 19428 22802 19440
rect 23382 19428 23388 19440
rect 22796 19400 23388 19428
rect 22796 19388 22802 19400
rect 23382 19388 23388 19400
rect 23440 19388 23446 19440
rect 27614 19428 27620 19440
rect 27575 19400 27620 19428
rect 27614 19388 27620 19400
rect 27672 19388 27678 19440
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 22640 19363 22698 19369
rect 22640 19329 22652 19363
rect 22686 19360 22698 19363
rect 22922 19360 22928 19372
rect 22686 19332 22928 19360
rect 22686 19329 22698 19332
rect 22640 19323 22698 19329
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 26142 19360 26148 19372
rect 24351 19332 26148 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 26142 19320 26148 19332
rect 26200 19320 26206 19372
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 27816 19360 27844 19468
rect 30009 19465 30021 19468
rect 30055 19465 30067 19499
rect 33502 19496 33508 19508
rect 33463 19468 33508 19496
rect 30009 19459 30067 19465
rect 33502 19456 33508 19468
rect 33560 19456 33566 19508
rect 35066 19496 35072 19508
rect 35027 19468 35072 19496
rect 35066 19456 35072 19468
rect 35124 19456 35130 19508
rect 35437 19499 35495 19505
rect 35437 19496 35449 19499
rect 35176 19468 35449 19496
rect 34790 19388 34796 19440
rect 34848 19428 34854 19440
rect 35176 19428 35204 19468
rect 35437 19465 35449 19468
rect 35483 19465 35495 19499
rect 38657 19499 38715 19505
rect 38657 19496 38669 19499
rect 35437 19459 35495 19465
rect 35728 19468 38669 19496
rect 34848 19400 35204 19428
rect 34848 19388 34854 19400
rect 27488 19332 27844 19360
rect 28813 19363 28871 19369
rect 27488 19320 27494 19332
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 30190 19360 30196 19372
rect 28859 19332 30196 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 30190 19320 30196 19332
rect 30248 19320 30254 19372
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19360 32367 19363
rect 35728 19360 35756 19468
rect 38657 19465 38669 19468
rect 38703 19465 38715 19499
rect 38657 19459 38715 19465
rect 40497 19499 40555 19505
rect 40497 19465 40509 19499
rect 40543 19496 40555 19499
rect 40862 19496 40868 19508
rect 40543 19468 40868 19496
rect 40543 19465 40555 19468
rect 40497 19459 40555 19465
rect 40862 19456 40868 19468
rect 40920 19456 40926 19508
rect 40972 19468 41184 19496
rect 35802 19388 35808 19440
rect 35860 19428 35866 19440
rect 40972 19428 41000 19468
rect 35860 19400 36492 19428
rect 35860 19388 35866 19400
rect 36464 19369 36492 19400
rect 36556 19400 41000 19428
rect 41156 19428 41184 19468
rect 41230 19456 41236 19508
rect 41288 19496 41294 19508
rect 41690 19496 41696 19508
rect 41288 19468 41696 19496
rect 41288 19456 41294 19468
rect 41690 19456 41696 19468
rect 41748 19496 41754 19508
rect 48222 19496 48228 19508
rect 41748 19468 48228 19496
rect 41748 19456 41754 19468
rect 48222 19456 48228 19468
rect 48280 19456 48286 19508
rect 48958 19456 48964 19508
rect 49016 19496 49022 19508
rect 58253 19499 58311 19505
rect 58253 19496 58265 19499
rect 49016 19468 58265 19496
rect 49016 19456 49022 19468
rect 58253 19465 58265 19468
rect 58299 19465 58311 19499
rect 58253 19459 58311 19465
rect 47762 19428 47768 19440
rect 41156 19400 47768 19428
rect 36449 19363 36507 19369
rect 32355 19332 35756 19360
rect 35820 19332 36400 19360
rect 32355 19329 32367 19332
rect 32309 19323 32367 19329
rect 27709 19295 27767 19301
rect 22204 19264 22416 19292
rect 19484 19252 19490 19264
rect 22388 19236 22416 19264
rect 27709 19261 27721 19295
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 31570 19292 31576 19304
rect 27939 19264 31576 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 18506 19224 18512 19236
rect 18419 19196 18512 19224
rect 18506 19184 18512 19196
rect 18564 19224 18570 19236
rect 19978 19224 19984 19236
rect 18564 19196 19984 19224
rect 18564 19184 18570 19196
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 20070 19184 20076 19236
rect 20128 19224 20134 19236
rect 20128 19196 22094 19224
rect 20128 19184 20134 19196
rect 2409 19159 2467 19165
rect 2409 19125 2421 19159
rect 2455 19156 2467 19159
rect 7558 19156 7564 19168
rect 2455 19128 7564 19156
rect 2455 19125 2467 19128
rect 2409 19119 2467 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 17497 19159 17555 19165
rect 17497 19125 17509 19159
rect 17543 19156 17555 19159
rect 20622 19156 20628 19168
rect 17543 19128 20628 19156
rect 17543 19125 17555 19128
rect 17497 19119 17555 19125
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 22066 19156 22094 19196
rect 22370 19184 22376 19236
rect 22428 19184 22434 19236
rect 24302 19184 24308 19236
rect 24360 19224 24366 19236
rect 27614 19224 27620 19236
rect 24360 19196 27620 19224
rect 24360 19184 24366 19196
rect 27614 19184 27620 19196
rect 27672 19184 27678 19236
rect 27724 19224 27752 19255
rect 31570 19252 31576 19264
rect 31628 19252 31634 19304
rect 35526 19252 35532 19304
rect 35584 19292 35590 19304
rect 35710 19292 35716 19304
rect 35584 19264 35629 19292
rect 35671 19264 35716 19292
rect 35584 19252 35590 19264
rect 35710 19252 35716 19264
rect 35768 19252 35774 19304
rect 27982 19224 27988 19236
rect 27724 19196 27988 19224
rect 27982 19184 27988 19196
rect 28040 19184 28046 19236
rect 28350 19184 28356 19236
rect 28408 19224 28414 19236
rect 35820 19224 35848 19332
rect 36262 19292 36268 19304
rect 36223 19264 36268 19292
rect 36262 19252 36268 19264
rect 36320 19252 36326 19304
rect 36372 19292 36400 19332
rect 36449 19329 36461 19363
rect 36495 19329 36507 19363
rect 36449 19323 36507 19329
rect 36556 19292 36584 19400
rect 47762 19388 47768 19400
rect 47820 19388 47826 19440
rect 48130 19428 48136 19440
rect 48091 19400 48136 19428
rect 48130 19388 48136 19400
rect 48188 19388 48194 19440
rect 48682 19388 48688 19440
rect 48740 19428 48746 19440
rect 58158 19428 58164 19440
rect 48740 19400 58164 19428
rect 48740 19388 48746 19400
rect 58158 19388 58164 19400
rect 58216 19388 58222 19440
rect 37366 19320 37372 19372
rect 37424 19360 37430 19372
rect 37461 19363 37519 19369
rect 37461 19360 37473 19363
rect 37424 19332 37473 19360
rect 37424 19320 37430 19332
rect 37461 19329 37473 19332
rect 37507 19360 37519 19363
rect 40865 19363 40923 19369
rect 40865 19360 40877 19363
rect 37507 19332 40877 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 40865 19329 40877 19332
rect 40911 19329 40923 19363
rect 41414 19360 41420 19372
rect 40865 19323 40923 19329
rect 41156 19332 41420 19360
rect 36372 19264 36584 19292
rect 37090 19252 37096 19304
rect 37148 19292 37154 19304
rect 40678 19292 40684 19304
rect 37148 19264 40684 19292
rect 37148 19252 37154 19264
rect 40678 19252 40684 19264
rect 40736 19252 40742 19304
rect 40586 19224 40592 19236
rect 28408 19196 35848 19224
rect 35912 19196 40592 19224
rect 28408 19184 28414 19196
rect 28074 19156 28080 19168
rect 22066 19128 28080 19156
rect 28074 19116 28080 19128
rect 28132 19116 28138 19168
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 35912 19156 35940 19196
rect 40586 19184 40592 19196
rect 40644 19184 40650 19236
rect 40880 19224 40908 19323
rect 40957 19295 41015 19301
rect 40957 19261 40969 19295
rect 41003 19292 41015 19295
rect 41046 19292 41052 19304
rect 41003 19264 41052 19292
rect 41003 19261 41015 19264
rect 40957 19255 41015 19261
rect 41046 19252 41052 19264
rect 41104 19252 41110 19304
rect 41156 19301 41184 19332
rect 41414 19320 41420 19332
rect 41472 19320 41478 19372
rect 42705 19363 42763 19369
rect 42705 19329 42717 19363
rect 42751 19360 42763 19363
rect 43898 19360 43904 19372
rect 42751 19332 43904 19360
rect 42751 19329 42763 19332
rect 42705 19323 42763 19329
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 47854 19320 47860 19372
rect 47912 19360 47918 19372
rect 47912 19332 47957 19360
rect 47912 19320 47918 19332
rect 48038 19320 48044 19372
rect 48096 19360 48102 19372
rect 48271 19363 48329 19369
rect 48096 19332 48141 19360
rect 48096 19320 48102 19332
rect 48271 19329 48283 19363
rect 48317 19360 48329 19363
rect 48866 19360 48872 19372
rect 48317 19332 48443 19360
rect 48827 19332 48872 19360
rect 48317 19329 48329 19332
rect 48271 19323 48329 19329
rect 41141 19295 41199 19301
rect 41141 19261 41153 19295
rect 41187 19261 41199 19295
rect 41141 19255 41199 19261
rect 41230 19252 41236 19304
rect 41288 19292 41294 19304
rect 46106 19292 46112 19304
rect 41288 19264 46112 19292
rect 41288 19252 41294 19264
rect 46106 19252 46112 19264
rect 46164 19252 46170 19304
rect 48415 19292 48443 19332
rect 48866 19320 48872 19332
rect 48924 19320 48930 19372
rect 49050 19360 49056 19372
rect 49011 19332 49056 19360
rect 49050 19320 49056 19332
rect 49108 19320 49114 19372
rect 58066 19360 58072 19372
rect 58027 19332 58072 19360
rect 58066 19320 58072 19332
rect 58124 19320 58130 19372
rect 49142 19292 49148 19304
rect 48415 19264 49148 19292
rect 49142 19252 49148 19264
rect 49200 19252 49206 19304
rect 41874 19224 41880 19236
rect 40880 19196 41880 19224
rect 41874 19184 41880 19196
rect 41932 19184 41938 19236
rect 48130 19184 48136 19236
rect 48188 19224 48194 19236
rect 58250 19224 58256 19236
rect 48188 19196 58256 19224
rect 48188 19184 48194 19196
rect 58250 19184 58256 19196
rect 58308 19184 58314 19236
rect 36630 19156 36636 19168
rect 33192 19128 35940 19156
rect 36591 19128 36636 19156
rect 33192 19116 33198 19128
rect 36630 19116 36636 19128
rect 36688 19116 36694 19168
rect 40126 19116 40132 19168
rect 40184 19156 40190 19168
rect 40221 19159 40279 19165
rect 40221 19156 40233 19159
rect 40184 19128 40233 19156
rect 40184 19116 40190 19128
rect 40221 19125 40233 19128
rect 40267 19156 40279 19159
rect 41046 19156 41052 19168
rect 40267 19128 41052 19156
rect 40267 19125 40279 19128
rect 40221 19119 40279 19125
rect 41046 19116 41052 19128
rect 41104 19116 41110 19168
rect 41230 19116 41236 19168
rect 41288 19156 41294 19168
rect 42978 19156 42984 19168
rect 41288 19128 42984 19156
rect 41288 19116 41294 19128
rect 42978 19116 42984 19128
rect 43036 19116 43042 19168
rect 48409 19159 48467 19165
rect 48409 19125 48421 19159
rect 48455 19156 48467 19159
rect 48590 19156 48596 19168
rect 48455 19128 48596 19156
rect 48455 19125 48467 19128
rect 48409 19119 48467 19125
rect 48590 19116 48596 19128
rect 48648 19116 48654 19168
rect 49234 19156 49240 19168
rect 49195 19128 49240 19156
rect 49234 19116 49240 19128
rect 49292 19116 49298 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 22002 18952 22008 18964
rect 18708 18924 22008 18952
rect 15930 18776 15936 18828
rect 15988 18816 15994 18828
rect 17586 18816 17592 18828
rect 15988 18788 16988 18816
rect 17547 18788 17592 18816
rect 15988 18776 15994 18788
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 16666 18748 16672 18760
rect 1627 18720 2452 18748
rect 16627 18720 16672 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 2424 18621 2452 18720
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18717 16911 18751
rect 16960 18748 16988 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 17862 18816 17868 18828
rect 17823 18788 17868 18816
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 18506 18816 18512 18828
rect 18467 18788 18512 18816
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 18708 18825 18736 18924
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22462 18912 22468 18964
rect 22520 18952 22526 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22520 18924 22937 18952
rect 22520 18912 22526 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23106 18912 23112 18964
rect 23164 18952 23170 18964
rect 24302 18952 24308 18964
rect 23164 18924 24308 18952
rect 23164 18912 23170 18924
rect 24302 18912 24308 18924
rect 24360 18912 24366 18964
rect 26050 18952 26056 18964
rect 24596 18924 26056 18952
rect 21269 18887 21327 18893
rect 21269 18853 21281 18887
rect 21315 18884 21327 18887
rect 24596 18884 24624 18924
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 27614 18912 27620 18964
rect 27672 18952 27678 18964
rect 30006 18952 30012 18964
rect 27672 18924 30012 18952
rect 27672 18912 27678 18924
rect 30006 18912 30012 18924
rect 30064 18912 30070 18964
rect 30190 18912 30196 18964
rect 30248 18952 30254 18964
rect 32585 18955 32643 18961
rect 32585 18952 32597 18955
rect 30248 18924 32597 18952
rect 30248 18912 30254 18924
rect 32585 18921 32597 18924
rect 32631 18921 32643 18955
rect 32585 18915 32643 18921
rect 34422 18912 34428 18964
rect 34480 18952 34486 18964
rect 35802 18952 35808 18964
rect 34480 18924 35808 18952
rect 34480 18912 34486 18924
rect 35802 18912 35808 18924
rect 35860 18912 35866 18964
rect 48409 18955 48467 18961
rect 36556 18924 45692 18952
rect 21315 18856 24624 18884
rect 21315 18853 21327 18856
rect 21269 18847 21327 18853
rect 26418 18844 26424 18896
rect 26476 18884 26482 18896
rect 28350 18884 28356 18896
rect 26476 18856 28356 18884
rect 26476 18844 26482 18856
rect 28350 18844 28356 18856
rect 28408 18844 28414 18896
rect 30285 18887 30343 18893
rect 30285 18853 30297 18887
rect 30331 18884 30343 18887
rect 36556 18884 36584 18924
rect 30331 18856 36584 18884
rect 30331 18853 30343 18856
rect 30285 18847 30343 18853
rect 39390 18844 39396 18896
rect 39448 18884 39454 18896
rect 39669 18887 39727 18893
rect 39669 18884 39681 18887
rect 39448 18856 39681 18884
rect 39448 18844 39454 18856
rect 39669 18853 39681 18856
rect 39715 18884 39727 18887
rect 40126 18884 40132 18896
rect 39715 18856 40132 18884
rect 39715 18853 39727 18856
rect 39669 18847 39727 18853
rect 40126 18844 40132 18856
rect 40184 18844 40190 18896
rect 41874 18884 41880 18896
rect 41835 18856 41880 18884
rect 41874 18844 41880 18856
rect 41932 18844 41938 18896
rect 42429 18887 42487 18893
rect 42429 18853 42441 18887
rect 42475 18884 42487 18887
rect 44082 18884 44088 18896
rect 42475 18856 44088 18884
rect 42475 18853 42487 18856
rect 42429 18847 42487 18853
rect 44082 18844 44088 18856
rect 44140 18844 44146 18896
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 18831 18788 20024 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 17310 18748 17316 18760
rect 16960 18720 17316 18748
rect 16853 18711 16911 18717
rect 16776 18680 16804 18708
rect 2746 18652 16804 18680
rect 16868 18680 16896 18711
rect 17310 18708 17316 18720
rect 17368 18748 17374 18760
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17368 18720 17509 18748
rect 17368 18708 17374 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 18472 18720 18613 18748
rect 18472 18708 18478 18720
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 19484 18720 19901 18748
rect 19484 18708 19490 18720
rect 19889 18717 19901 18720
rect 19935 18717 19947 18751
rect 19996 18748 20024 18788
rect 20916 18788 23336 18816
rect 19996 18720 20484 18748
rect 19889 18711 19947 18717
rect 19978 18680 19984 18692
rect 16868 18652 19984 18680
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2746 18612 2774 18652
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 20156 18683 20214 18689
rect 20156 18649 20168 18683
rect 20202 18680 20214 18683
rect 20346 18680 20352 18692
rect 20202 18652 20352 18680
rect 20202 18649 20214 18652
rect 20156 18643 20214 18649
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 20456 18680 20484 18720
rect 20530 18708 20536 18760
rect 20588 18748 20594 18760
rect 20916 18748 20944 18788
rect 21726 18748 21732 18760
rect 20588 18720 20944 18748
rect 21687 18720 21732 18748
rect 20588 18708 20594 18720
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 23308 18680 23336 18788
rect 23382 18776 23388 18828
rect 23440 18816 23446 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 23440 18788 24593 18816
rect 23440 18776 23446 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 26050 18776 26056 18828
rect 26108 18816 26114 18828
rect 26108 18788 31432 18816
rect 26108 18776 26114 18788
rect 24854 18757 24860 18760
rect 24848 18748 24860 18757
rect 24815 18720 24860 18748
rect 24848 18711 24860 18720
rect 24854 18708 24860 18711
rect 24912 18708 24918 18760
rect 26878 18748 26884 18760
rect 26839 18720 26884 18748
rect 26878 18708 26884 18720
rect 26936 18748 26942 18760
rect 28442 18748 28448 18760
rect 26936 18720 28448 18748
rect 26936 18708 26942 18720
rect 28442 18708 28448 18720
rect 28500 18748 28506 18760
rect 29822 18748 29828 18760
rect 28500 18720 29828 18748
rect 28500 18708 28506 18720
rect 29822 18708 29828 18720
rect 29880 18748 29886 18760
rect 31404 18757 31432 18788
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 36909 18819 36967 18825
rect 36909 18816 36921 18819
rect 33100 18788 36921 18816
rect 33100 18776 33106 18788
rect 36909 18785 36921 18788
rect 36955 18785 36967 18819
rect 36909 18779 36967 18785
rect 38102 18776 38108 18828
rect 38160 18816 38166 18828
rect 39117 18819 39175 18825
rect 39117 18816 39129 18819
rect 38160 18788 39129 18816
rect 38160 18776 38166 18788
rect 39117 18785 39129 18788
rect 39163 18785 39175 18819
rect 39117 18779 39175 18785
rect 30561 18751 30619 18757
rect 30561 18748 30573 18751
rect 29880 18720 30573 18748
rect 29880 18708 29886 18720
rect 30561 18717 30573 18720
rect 30607 18717 30619 18751
rect 30561 18711 30619 18717
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 34790 18748 34796 18760
rect 31435 18720 34796 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 34790 18708 34796 18720
rect 34848 18708 34854 18760
rect 34882 18708 34888 18760
rect 34940 18748 34946 18760
rect 35069 18751 35127 18757
rect 34940 18720 34985 18748
rect 34940 18708 34946 18720
rect 35069 18717 35081 18751
rect 35115 18717 35127 18751
rect 35802 18748 35808 18760
rect 35763 18720 35808 18748
rect 35069 18711 35127 18717
rect 27614 18680 27620 18692
rect 20456 18652 23244 18680
rect 23308 18652 27620 18680
rect 2455 18584 2774 18612
rect 16761 18615 16819 18621
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 18230 18612 18236 18624
rect 16807 18584 18236 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 18325 18615 18383 18621
rect 18325 18581 18337 18615
rect 18371 18612 18383 18615
rect 21082 18612 21088 18624
rect 18371 18584 21088 18612
rect 18371 18581 18383 18584
rect 18325 18575 18383 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 23106 18612 23112 18624
rect 21324 18584 23112 18612
rect 21324 18572 21330 18584
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 23216 18612 23244 18652
rect 27614 18640 27620 18652
rect 27672 18640 27678 18692
rect 30006 18640 30012 18692
rect 30064 18680 30070 18692
rect 30064 18652 30696 18680
rect 30064 18640 30070 18652
rect 24578 18612 24584 18624
rect 23216 18584 24584 18612
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25961 18615 26019 18621
rect 25961 18581 25973 18615
rect 26007 18612 26019 18615
rect 26050 18612 26056 18624
rect 26007 18584 26056 18612
rect 26007 18581 26019 18584
rect 25961 18575 26019 18581
rect 26050 18572 26056 18584
rect 26108 18572 26114 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 28077 18615 28135 18621
rect 28077 18612 28089 18615
rect 26292 18584 28089 18612
rect 26292 18572 26298 18584
rect 28077 18581 28089 18584
rect 28123 18581 28135 18615
rect 30668 18612 30696 18652
rect 30834 18640 30840 18692
rect 30892 18680 30898 18692
rect 33962 18680 33968 18692
rect 30892 18652 33968 18680
rect 30892 18640 30898 18652
rect 33962 18640 33968 18652
rect 34020 18640 34026 18692
rect 34698 18640 34704 18692
rect 34756 18680 34762 18692
rect 35084 18680 35112 18711
rect 35802 18708 35808 18720
rect 35860 18748 35866 18760
rect 38838 18748 38844 18760
rect 35860 18720 38844 18748
rect 35860 18708 35866 18720
rect 38838 18708 38844 18720
rect 38896 18708 38902 18760
rect 38933 18751 38991 18757
rect 38933 18717 38945 18751
rect 38979 18748 38991 18751
rect 39206 18748 39212 18760
rect 38979 18720 39212 18748
rect 38979 18717 38991 18720
rect 38933 18711 38991 18717
rect 39206 18708 39212 18720
rect 39264 18708 39270 18760
rect 40497 18751 40555 18757
rect 40497 18717 40509 18751
rect 40543 18748 40555 18751
rect 40586 18748 40592 18760
rect 40543 18720 40592 18748
rect 40543 18717 40555 18720
rect 40497 18711 40555 18717
rect 40586 18708 40592 18720
rect 40644 18708 40650 18760
rect 40770 18757 40776 18760
rect 40764 18748 40776 18757
rect 40731 18720 40776 18748
rect 40764 18711 40776 18720
rect 40770 18708 40776 18711
rect 40828 18708 40834 18760
rect 41892 18748 41920 18844
rect 42978 18816 42984 18828
rect 42939 18788 42984 18816
rect 42978 18776 42984 18788
rect 43036 18776 43042 18828
rect 42797 18751 42855 18757
rect 42797 18748 42809 18751
rect 41892 18720 42809 18748
rect 42797 18717 42809 18720
rect 42843 18717 42855 18751
rect 43622 18748 43628 18760
rect 43583 18720 43628 18748
rect 42797 18711 42855 18717
rect 43622 18708 43628 18720
rect 43680 18708 43686 18760
rect 43990 18748 43996 18760
rect 43951 18720 43996 18748
rect 43990 18708 43996 18720
rect 44048 18708 44054 18760
rect 45373 18751 45431 18757
rect 45373 18717 45385 18751
rect 45419 18717 45431 18751
rect 45554 18748 45560 18760
rect 45515 18720 45560 18748
rect 45373 18711 45431 18717
rect 34756 18652 35112 18680
rect 34756 18640 34762 18652
rect 40678 18640 40684 18692
rect 40736 18680 40742 18692
rect 42889 18683 42947 18689
rect 42889 18680 42901 18683
rect 40736 18652 42901 18680
rect 40736 18640 40742 18652
rect 42889 18649 42901 18652
rect 42935 18649 42947 18683
rect 42889 18643 42947 18649
rect 43070 18640 43076 18692
rect 43128 18680 43134 18692
rect 43809 18683 43867 18689
rect 43809 18680 43821 18683
rect 43128 18652 43821 18680
rect 43128 18640 43134 18652
rect 43809 18649 43821 18652
rect 43855 18649 43867 18683
rect 43809 18643 43867 18649
rect 43901 18683 43959 18689
rect 43901 18649 43913 18683
rect 43947 18680 43959 18683
rect 44266 18680 44272 18692
rect 43947 18652 44272 18680
rect 43947 18649 43959 18652
rect 43901 18643 43959 18649
rect 44266 18640 44272 18652
rect 44324 18640 44330 18692
rect 45388 18680 45416 18711
rect 45554 18708 45560 18720
rect 45612 18708 45618 18760
rect 45664 18748 45692 18924
rect 48409 18921 48421 18955
rect 48455 18952 48467 18955
rect 49050 18952 49056 18964
rect 48455 18924 49056 18952
rect 48455 18921 48467 18924
rect 48409 18915 48467 18921
rect 49050 18912 49056 18924
rect 49108 18912 49114 18964
rect 48038 18844 48044 18896
rect 48096 18884 48102 18896
rect 48096 18856 49004 18884
rect 48096 18844 48102 18856
rect 46106 18776 46112 18828
rect 46164 18816 46170 18828
rect 48590 18816 48596 18828
rect 46164 18788 48596 18816
rect 46164 18776 46170 18788
rect 48590 18776 48596 18788
rect 48648 18776 48654 18828
rect 48976 18816 49004 18856
rect 48976 18788 49050 18816
rect 47857 18751 47915 18757
rect 47857 18748 47869 18751
rect 45664 18720 47869 18748
rect 47857 18717 47869 18720
rect 47903 18717 47915 18751
rect 48222 18748 48228 18760
rect 48183 18720 48228 18748
rect 47857 18711 47915 18717
rect 48222 18708 48228 18720
rect 48280 18708 48286 18760
rect 48682 18708 48688 18760
rect 48740 18748 48746 18760
rect 49022 18757 49050 18788
rect 49142 18776 49148 18828
rect 49200 18816 49206 18828
rect 49200 18788 49280 18816
rect 49200 18776 49206 18788
rect 49252 18757 49280 18788
rect 48869 18751 48927 18757
rect 48869 18748 48881 18751
rect 48740 18720 48881 18748
rect 48740 18708 48746 18720
rect 48869 18717 48881 18720
rect 48915 18717 48927 18751
rect 48869 18711 48927 18717
rect 49007 18751 49065 18757
rect 49007 18717 49019 18751
rect 49053 18717 49065 18751
rect 49007 18711 49065 18717
rect 49237 18751 49295 18757
rect 49237 18717 49249 18751
rect 49283 18717 49295 18751
rect 57882 18748 57888 18760
rect 57843 18720 57888 18748
rect 49237 18711 49295 18717
rect 57882 18708 57888 18720
rect 57940 18708 57946 18760
rect 46842 18680 46848 18692
rect 45388 18652 46848 18680
rect 46842 18640 46848 18652
rect 46900 18640 46906 18692
rect 48038 18680 48044 18692
rect 47999 18652 48044 18680
rect 48038 18640 48044 18652
rect 48096 18640 48102 18692
rect 48130 18640 48136 18692
rect 48188 18680 48194 18692
rect 49145 18683 49203 18689
rect 48188 18652 48233 18680
rect 48188 18640 48194 18652
rect 49145 18649 49157 18683
rect 49191 18680 49203 18683
rect 49878 18680 49884 18692
rect 49191 18652 49884 18680
rect 49191 18649 49203 18652
rect 49145 18643 49203 18649
rect 49878 18640 49884 18652
rect 49936 18680 49942 18692
rect 50706 18680 50712 18692
rect 49936 18652 50712 18680
rect 49936 18640 49942 18652
rect 50706 18640 50712 18652
rect 50764 18640 50770 18692
rect 58158 18680 58164 18692
rect 58119 18652 58164 18680
rect 58158 18640 58164 18652
rect 58216 18640 58222 18692
rect 30742 18612 30748 18624
rect 30668 18584 30748 18612
rect 28077 18575 28135 18581
rect 30742 18572 30748 18584
rect 30800 18612 30806 18624
rect 30800 18584 30893 18612
rect 30800 18572 30806 18584
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 35253 18615 35311 18621
rect 35253 18612 35265 18615
rect 34572 18584 35265 18612
rect 34572 18572 34578 18584
rect 35253 18581 35265 18584
rect 35299 18581 35311 18615
rect 38562 18612 38568 18624
rect 38523 18584 38568 18612
rect 35253 18575 35311 18581
rect 38562 18572 38568 18584
rect 38620 18572 38626 18624
rect 39025 18615 39083 18621
rect 39025 18581 39037 18615
rect 39071 18612 39083 18615
rect 39206 18612 39212 18624
rect 39071 18584 39212 18612
rect 39071 18581 39083 18584
rect 39025 18575 39083 18581
rect 39206 18572 39212 18584
rect 39264 18572 39270 18624
rect 42978 18572 42984 18624
rect 43036 18612 43042 18624
rect 44177 18615 44235 18621
rect 44177 18612 44189 18615
rect 43036 18584 44189 18612
rect 43036 18572 43042 18584
rect 44177 18581 44189 18584
rect 44223 18581 44235 18615
rect 45738 18612 45744 18624
rect 45699 18584 45744 18612
rect 44177 18575 44235 18581
rect 45738 18572 45744 18584
rect 45796 18572 45802 18624
rect 45922 18572 45928 18624
rect 45980 18612 45986 18624
rect 48682 18612 48688 18624
rect 45980 18584 48688 18612
rect 45980 18572 45986 18584
rect 48682 18572 48688 18584
rect 48740 18572 48746 18624
rect 49418 18612 49424 18624
rect 49379 18584 49424 18612
rect 49418 18572 49424 18584
rect 49476 18572 49482 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 17126 18408 17132 18420
rect 7616 18380 17132 18408
rect 7616 18368 7622 18380
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 18506 18408 18512 18420
rect 17552 18380 18512 18408
rect 17552 18368 17558 18380
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 18601 18411 18659 18417
rect 18601 18377 18613 18411
rect 18647 18408 18659 18411
rect 24302 18408 24308 18420
rect 18647 18380 24308 18408
rect 18647 18377 18659 18380
rect 18601 18371 18659 18377
rect 24302 18368 24308 18380
rect 24360 18368 24366 18420
rect 24394 18368 24400 18420
rect 24452 18408 24458 18420
rect 24489 18411 24547 18417
rect 24489 18408 24501 18411
rect 24452 18380 24501 18408
rect 24452 18368 24458 18380
rect 24489 18377 24501 18380
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 27062 18368 27068 18420
rect 27120 18408 27126 18420
rect 27157 18411 27215 18417
rect 27157 18408 27169 18411
rect 27120 18380 27169 18408
rect 27120 18368 27126 18380
rect 27157 18377 27169 18380
rect 27203 18377 27215 18411
rect 27157 18371 27215 18377
rect 27890 18368 27896 18420
rect 27948 18408 27954 18420
rect 29457 18411 29515 18417
rect 29457 18408 29469 18411
rect 27948 18380 29469 18408
rect 27948 18368 27954 18380
rect 29457 18377 29469 18380
rect 29503 18377 29515 18411
rect 31386 18408 31392 18420
rect 31347 18380 31392 18408
rect 29457 18371 29515 18377
rect 31386 18368 31392 18380
rect 31444 18368 31450 18420
rect 34790 18368 34796 18420
rect 34848 18408 34854 18420
rect 36449 18411 36507 18417
rect 36449 18408 36461 18411
rect 34848 18380 36461 18408
rect 34848 18368 34854 18380
rect 36449 18377 36461 18380
rect 36495 18408 36507 18411
rect 37182 18408 37188 18420
rect 36495 18380 37188 18408
rect 36495 18377 36507 18380
rect 36449 18371 36507 18377
rect 37182 18368 37188 18380
rect 37240 18368 37246 18420
rect 37458 18408 37464 18420
rect 37419 18380 37464 18408
rect 37458 18368 37464 18380
rect 37516 18368 37522 18420
rect 38838 18368 38844 18420
rect 38896 18408 38902 18420
rect 40129 18411 40187 18417
rect 40129 18408 40141 18411
rect 38896 18380 40141 18408
rect 38896 18368 38902 18380
rect 40129 18377 40141 18380
rect 40175 18377 40187 18411
rect 40129 18371 40187 18377
rect 40681 18411 40739 18417
rect 40681 18377 40693 18411
rect 40727 18408 40739 18411
rect 43622 18408 43628 18420
rect 40727 18380 43628 18408
rect 40727 18377 40739 18380
rect 40681 18371 40739 18377
rect 17862 18300 17868 18352
rect 17920 18340 17926 18352
rect 17920 18312 19196 18340
rect 17920 18300 17926 18312
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 14240 18244 15393 18272
rect 14240 18232 14246 18244
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 15746 18272 15752 18284
rect 15611 18244 15752 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 19168 18281 19196 18312
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 21266 18340 21272 18352
rect 20036 18312 21272 18340
rect 20036 18300 20042 18312
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 22649 18343 22707 18349
rect 22649 18309 22661 18343
rect 22695 18340 22707 18343
rect 24026 18340 24032 18352
rect 22695 18312 24032 18340
rect 22695 18309 22707 18312
rect 22649 18303 22707 18309
rect 24026 18300 24032 18312
rect 24084 18300 24090 18352
rect 25866 18300 25872 18352
rect 25924 18340 25930 18352
rect 26418 18340 26424 18352
rect 25924 18312 26424 18340
rect 25924 18300 25930 18312
rect 26418 18300 26424 18312
rect 26476 18300 26482 18352
rect 27522 18300 27528 18352
rect 27580 18340 27586 18352
rect 35336 18343 35394 18349
rect 27580 18312 31754 18340
rect 27580 18300 27586 18312
rect 17488 18275 17546 18281
rect 17488 18241 17500 18275
rect 17534 18272 17546 18275
rect 19153 18275 19211 18281
rect 17534 18244 18920 18272
rect 17534 18241 17546 18244
rect 17488 18235 17546 18241
rect 17218 18204 17224 18216
rect 17179 18176 17224 18204
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 18892 18204 18920 18244
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 23293 18275 23351 18281
rect 23293 18272 23305 18275
rect 21140 18244 23305 18272
rect 21140 18232 21146 18244
rect 23293 18241 23305 18244
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 26237 18275 26295 18281
rect 26237 18241 26249 18275
rect 26283 18272 26295 18275
rect 26283 18244 27108 18272
rect 26283 18241 26295 18244
rect 26237 18235 26295 18241
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 18892 18176 20269 18204
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 20257 18167 20315 18173
rect 22066 18176 22569 18204
rect 13722 18096 13728 18148
rect 13780 18136 13786 18148
rect 13780 18108 15884 18136
rect 13780 18096 13786 18108
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 10836 18040 15761 18068
rect 10836 18028 10842 18040
rect 15749 18037 15761 18040
rect 15795 18037 15807 18071
rect 15856 18068 15884 18108
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 20530 18136 20536 18148
rect 18564 18108 20536 18136
rect 18564 18096 18570 18108
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 22066 18068 22094 18176
rect 22557 18173 22569 18176
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 22741 18207 22799 18213
rect 22741 18173 22753 18207
rect 22787 18204 22799 18207
rect 26050 18204 26056 18216
rect 22787 18176 26056 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 26050 18164 26056 18176
rect 26108 18164 26114 18216
rect 26329 18207 26387 18213
rect 26329 18173 26341 18207
rect 26375 18204 26387 18207
rect 27080 18204 27108 18244
rect 27154 18232 27160 18284
rect 27212 18278 27218 18284
rect 27334 18281 27392 18287
rect 27334 18278 27346 18281
rect 27212 18250 27346 18278
rect 27212 18232 27218 18250
rect 27334 18247 27346 18250
rect 27380 18247 27392 18281
rect 27614 18272 27620 18284
rect 27334 18241 27392 18247
rect 27575 18244 27620 18272
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 27801 18275 27859 18281
rect 27801 18241 27813 18275
rect 27847 18272 27859 18275
rect 27890 18272 27896 18284
rect 27847 18244 27896 18272
rect 27847 18241 27859 18244
rect 27801 18235 27859 18241
rect 27890 18232 27896 18244
rect 27948 18232 27954 18284
rect 28258 18272 28264 18284
rect 28219 18244 28264 18272
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 29822 18232 29828 18284
rect 29880 18272 29886 18284
rect 30650 18272 30656 18284
rect 29880 18244 30656 18272
rect 29880 18232 29886 18244
rect 30650 18232 30656 18244
rect 30708 18232 30714 18284
rect 31726 18272 31754 18312
rect 35336 18309 35348 18343
rect 35382 18340 35394 18343
rect 36630 18340 36636 18352
rect 35382 18312 36636 18340
rect 35382 18309 35394 18312
rect 35336 18303 35394 18309
rect 36630 18300 36636 18312
rect 36688 18300 36694 18352
rect 40144 18340 40172 18371
rect 43622 18368 43628 18380
rect 43680 18368 43686 18420
rect 44266 18408 44272 18420
rect 44227 18380 44272 18408
rect 44266 18368 44272 18380
rect 44324 18368 44330 18420
rect 45922 18408 45928 18420
rect 44376 18380 45928 18408
rect 41049 18343 41107 18349
rect 41049 18340 41061 18343
rect 38580 18312 39160 18340
rect 40144 18312 41061 18340
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 31726 18244 32321 18272
rect 32309 18241 32321 18244
rect 32355 18272 32367 18275
rect 37274 18272 37280 18284
rect 32355 18244 37280 18272
rect 32355 18241 32367 18244
rect 32309 18235 32367 18241
rect 37274 18232 37280 18244
rect 37332 18272 37338 18284
rect 37829 18275 37887 18281
rect 37829 18272 37841 18275
rect 37332 18244 37841 18272
rect 37332 18232 37338 18244
rect 37829 18241 37841 18244
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 26375 18176 27016 18204
rect 27080 18176 27200 18204
rect 26375 18173 26387 18176
rect 26329 18167 26387 18173
rect 22186 18096 22192 18148
rect 22244 18136 22250 18148
rect 22244 18108 22289 18136
rect 22244 18096 22250 18108
rect 24026 18096 24032 18148
rect 24084 18136 24090 18148
rect 24670 18136 24676 18148
rect 24084 18108 24676 18136
rect 24084 18096 24090 18108
rect 24670 18096 24676 18108
rect 24728 18096 24734 18148
rect 26142 18096 26148 18148
rect 26200 18136 26206 18148
rect 26605 18139 26663 18145
rect 26605 18136 26617 18139
rect 26200 18108 26617 18136
rect 26200 18096 26206 18108
rect 26605 18105 26617 18108
rect 26651 18105 26663 18139
rect 26605 18099 26663 18105
rect 15856 18040 22094 18068
rect 15749 18031 15807 18037
rect 23750 18028 23756 18080
rect 23808 18068 23814 18080
rect 26878 18068 26884 18080
rect 23808 18040 26884 18068
rect 23808 18028 23814 18040
rect 26878 18028 26884 18040
rect 26936 18028 26942 18080
rect 26988 18068 27016 18176
rect 27172 18136 27200 18176
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 30466 18204 30472 18216
rect 27488 18176 30472 18204
rect 27488 18164 27494 18176
rect 30466 18164 30472 18176
rect 30524 18164 30530 18216
rect 31110 18164 31116 18216
rect 31168 18204 31174 18216
rect 31481 18207 31539 18213
rect 31481 18204 31493 18207
rect 31168 18176 31493 18204
rect 31168 18164 31174 18176
rect 31481 18173 31493 18176
rect 31527 18173 31539 18207
rect 31481 18167 31539 18173
rect 31570 18164 31576 18216
rect 31628 18204 31634 18216
rect 31628 18176 31673 18204
rect 31628 18164 31634 18176
rect 34238 18164 34244 18216
rect 34296 18204 34302 18216
rect 35069 18207 35127 18213
rect 35069 18204 35081 18207
rect 34296 18176 35081 18204
rect 34296 18164 34302 18176
rect 35069 18173 35081 18176
rect 35115 18173 35127 18207
rect 37918 18204 37924 18216
rect 37879 18176 37924 18204
rect 35069 18167 35127 18173
rect 37918 18164 37924 18176
rect 37976 18164 37982 18216
rect 38105 18207 38163 18213
rect 38105 18173 38117 18207
rect 38151 18204 38163 18207
rect 38580 18204 38608 18312
rect 39022 18281 39028 18284
rect 39016 18272 39028 18281
rect 38983 18244 39028 18272
rect 39016 18235 39028 18244
rect 39022 18232 39028 18235
rect 39080 18232 39086 18284
rect 39132 18272 39160 18312
rect 41049 18309 41061 18312
rect 41095 18309 41107 18343
rect 44376 18340 44404 18380
rect 45922 18368 45928 18380
rect 45980 18368 45986 18420
rect 46750 18368 46756 18420
rect 46808 18408 46814 18420
rect 46845 18411 46903 18417
rect 46845 18408 46857 18411
rect 46808 18380 46857 18408
rect 46808 18368 46814 18380
rect 46845 18377 46857 18380
rect 46891 18377 46903 18411
rect 46845 18371 46903 18377
rect 48130 18368 48136 18420
rect 48188 18408 48194 18420
rect 49513 18411 49571 18417
rect 49513 18408 49525 18411
rect 48188 18380 49525 18408
rect 48188 18368 48194 18380
rect 49513 18377 49525 18380
rect 49559 18408 49571 18411
rect 57698 18408 57704 18420
rect 49559 18380 57704 18408
rect 49559 18377 49571 18380
rect 49513 18371 49571 18377
rect 57698 18368 57704 18380
rect 57756 18368 57762 18420
rect 58250 18408 58256 18420
rect 58211 18380 58256 18408
rect 58250 18368 58256 18380
rect 58308 18368 58314 18420
rect 45738 18349 45744 18352
rect 45732 18340 45744 18349
rect 41049 18303 41107 18309
rect 41386 18312 44404 18340
rect 45699 18312 45744 18340
rect 40310 18272 40316 18284
rect 39132 18244 40316 18272
rect 40310 18232 40316 18244
rect 40368 18232 40374 18284
rect 38151 18176 38608 18204
rect 38151 18173 38163 18176
rect 38105 18167 38163 18173
rect 31754 18136 31760 18148
rect 27172 18108 31760 18136
rect 31754 18096 31760 18108
rect 31812 18096 31818 18148
rect 37550 18096 37556 18148
rect 37608 18136 37614 18148
rect 38120 18136 38148 18167
rect 38654 18164 38660 18216
rect 38712 18204 38718 18216
rect 38749 18207 38807 18213
rect 38749 18204 38761 18207
rect 38712 18176 38761 18204
rect 38712 18164 38718 18176
rect 38749 18173 38761 18176
rect 38795 18173 38807 18207
rect 38749 18167 38807 18173
rect 40126 18164 40132 18216
rect 40184 18204 40190 18216
rect 40497 18207 40555 18213
rect 40497 18204 40509 18207
rect 40184 18176 40509 18204
rect 40184 18164 40190 18176
rect 40497 18173 40509 18176
rect 40543 18173 40555 18207
rect 40497 18167 40555 18173
rect 40862 18164 40868 18216
rect 40920 18204 40926 18216
rect 41141 18207 41199 18213
rect 41141 18204 41153 18207
rect 40920 18176 41153 18204
rect 40920 18164 40926 18176
rect 41141 18173 41153 18176
rect 41187 18173 41199 18207
rect 41141 18167 41199 18173
rect 41230 18164 41236 18216
rect 41288 18204 41294 18216
rect 41288 18176 41333 18204
rect 41288 18164 41294 18176
rect 41386 18136 41414 18312
rect 45732 18303 45744 18312
rect 45738 18300 45744 18303
rect 45796 18300 45802 18352
rect 47486 18300 47492 18352
rect 47544 18340 47550 18352
rect 48222 18340 48228 18352
rect 47544 18312 48228 18340
rect 47544 18300 47550 18312
rect 48222 18300 48228 18312
rect 48280 18300 48286 18352
rect 48400 18343 48458 18349
rect 48400 18309 48412 18343
rect 48446 18340 48458 18343
rect 49234 18340 49240 18352
rect 48446 18312 49240 18340
rect 48446 18309 48458 18312
rect 48400 18303 48458 18309
rect 49234 18300 49240 18312
rect 49292 18300 49298 18352
rect 41690 18272 41696 18284
rect 41651 18244 41696 18272
rect 41690 18232 41696 18244
rect 41748 18232 41754 18284
rect 42794 18232 42800 18284
rect 42852 18272 42858 18284
rect 43145 18275 43203 18281
rect 43145 18272 43157 18275
rect 42852 18244 43157 18272
rect 42852 18232 42858 18244
rect 43145 18241 43157 18244
rect 43191 18241 43203 18275
rect 43145 18235 43203 18241
rect 45480 18244 46704 18272
rect 42886 18204 42892 18216
rect 42847 18176 42892 18204
rect 42886 18164 42892 18176
rect 42944 18164 42950 18216
rect 44174 18164 44180 18216
rect 44232 18204 44238 18216
rect 45480 18213 45508 18244
rect 45465 18207 45523 18213
rect 45465 18204 45477 18207
rect 44232 18176 45477 18204
rect 44232 18164 44238 18176
rect 45465 18173 45477 18176
rect 45511 18173 45523 18207
rect 46676 18204 46704 18244
rect 46842 18232 46848 18284
rect 46900 18272 46906 18284
rect 46900 18244 49188 18272
rect 46900 18232 46906 18244
rect 48130 18204 48136 18216
rect 46676 18176 48136 18204
rect 45465 18167 45523 18173
rect 48130 18164 48136 18176
rect 48188 18164 48194 18216
rect 49160 18204 49188 18244
rect 49418 18232 49424 18284
rect 49476 18272 49482 18284
rect 50249 18275 50307 18281
rect 50249 18272 50261 18275
rect 49476 18244 50261 18272
rect 49476 18232 49482 18244
rect 50249 18241 50261 18244
rect 50295 18241 50307 18275
rect 58066 18272 58072 18284
rect 58027 18244 58072 18272
rect 50249 18235 50307 18241
rect 58066 18232 58072 18244
rect 58124 18232 58130 18284
rect 50065 18207 50123 18213
rect 50065 18204 50077 18207
rect 49160 18176 50077 18204
rect 50065 18173 50077 18176
rect 50111 18173 50123 18207
rect 50065 18167 50123 18173
rect 37608 18108 38148 18136
rect 39684 18108 41414 18136
rect 37608 18096 37614 18108
rect 27798 18068 27804 18080
rect 26988 18040 27804 18068
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 27890 18028 27896 18080
rect 27948 18068 27954 18080
rect 28350 18068 28356 18080
rect 27948 18040 28356 18068
rect 27948 18028 27954 18040
rect 28350 18028 28356 18040
rect 28408 18028 28414 18080
rect 28994 18028 29000 18080
rect 29052 18068 29058 18080
rect 30834 18068 30840 18080
rect 29052 18040 30840 18068
rect 29052 18028 29058 18040
rect 30834 18028 30840 18040
rect 30892 18028 30898 18080
rect 31018 18068 31024 18080
rect 30979 18040 31024 18068
rect 31018 18028 31024 18040
rect 31076 18028 31082 18080
rect 31386 18028 31392 18080
rect 31444 18068 31450 18080
rect 33134 18068 33140 18080
rect 31444 18040 33140 18068
rect 31444 18028 31450 18040
rect 33134 18028 33140 18040
rect 33192 18028 33198 18080
rect 33502 18068 33508 18080
rect 33463 18040 33508 18068
rect 33502 18028 33508 18040
rect 33560 18028 33566 18080
rect 33870 18028 33876 18080
rect 33928 18068 33934 18080
rect 39684 18068 39712 18108
rect 33928 18040 39712 18068
rect 33928 18028 33934 18040
rect 46198 18028 46204 18080
rect 46256 18068 46262 18080
rect 47026 18068 47032 18080
rect 46256 18040 47032 18068
rect 46256 18028 46262 18040
rect 47026 18028 47032 18040
rect 47084 18028 47090 18080
rect 49694 18028 49700 18080
rect 49752 18068 49758 18080
rect 50433 18071 50491 18077
rect 50433 18068 50445 18071
rect 49752 18040 50445 18068
rect 49752 18028 49758 18040
rect 50433 18037 50445 18040
rect 50479 18037 50491 18071
rect 50433 18031 50491 18037
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 16666 17864 16672 17876
rect 15028 17836 16672 17864
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 11054 17660 11060 17672
rect 1627 17632 11060 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 15028 17669 15056 17836
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 26786 17864 26792 17876
rect 20128 17836 24716 17864
rect 26747 17836 26792 17864
rect 20128 17824 20134 17836
rect 16022 17796 16028 17808
rect 15983 17768 16028 17796
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 20809 17799 20867 17805
rect 20809 17765 20821 17799
rect 20855 17765 20867 17799
rect 20809 17759 20867 17765
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15151 17700 19564 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14240 17632 14289 17660
rect 14240 17620 14246 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 15194 17660 15200 17672
rect 15155 17632 15200 17660
rect 15013 17623 15071 17629
rect 1854 17592 1860 17604
rect 1815 17564 1860 17592
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 11606 17484 11612 17536
rect 11664 17524 11670 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 11664 17496 14381 17524
rect 11664 17484 11670 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14476 17524 14504 17623
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 16574 17660 16580 17672
rect 16535 17632 16580 17660
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 19426 17660 19432 17672
rect 17276 17632 19432 17660
rect 17276 17620 17282 17632
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19536 17660 19564 17700
rect 20714 17660 20720 17672
rect 19536 17632 20720 17660
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 14826 17552 14832 17604
rect 14884 17592 14890 17604
rect 15657 17595 15715 17601
rect 15657 17592 15669 17595
rect 14884 17564 15669 17592
rect 14884 17552 14890 17564
rect 15657 17561 15669 17564
rect 15703 17561 15715 17595
rect 15657 17555 15715 17561
rect 18877 17595 18935 17601
rect 18877 17561 18889 17595
rect 18923 17592 18935 17595
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 18923 17564 19686 17592
rect 18923 17561 18935 17564
rect 18877 17555 18935 17561
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 20824 17592 20852 17759
rect 20898 17756 20904 17808
rect 20956 17796 20962 17808
rect 24394 17796 24400 17808
rect 20956 17768 24400 17796
rect 20956 17756 20962 17768
rect 24394 17756 24400 17768
rect 24452 17756 24458 17808
rect 24578 17796 24584 17808
rect 24539 17768 24584 17796
rect 24578 17756 24584 17768
rect 24636 17756 24642 17808
rect 21450 17688 21456 17740
rect 21508 17728 21514 17740
rect 24486 17728 24492 17740
rect 21508 17700 24492 17728
rect 21508 17688 21514 17700
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 24688 17728 24716 17836
rect 26786 17824 26792 17836
rect 26844 17824 26850 17876
rect 26878 17824 26884 17876
rect 26936 17864 26942 17876
rect 27890 17864 27896 17876
rect 26936 17836 27896 17864
rect 26936 17824 26942 17836
rect 27890 17824 27896 17836
rect 27948 17824 27954 17876
rect 28445 17867 28503 17873
rect 28445 17833 28457 17867
rect 28491 17864 28503 17867
rect 29178 17864 29184 17876
rect 28491 17836 29184 17864
rect 28491 17833 28503 17836
rect 28445 17827 28503 17833
rect 29178 17824 29184 17836
rect 29236 17824 29242 17876
rect 32490 17824 32496 17876
rect 32548 17864 32554 17876
rect 33045 17867 33103 17873
rect 33045 17864 33057 17867
rect 32548 17836 33057 17864
rect 32548 17824 32554 17836
rect 33045 17833 33057 17836
rect 33091 17833 33103 17867
rect 41138 17864 41144 17876
rect 33045 17827 33103 17833
rect 33152 17836 41144 17864
rect 33152 17796 33180 17836
rect 41138 17824 41144 17836
rect 41196 17824 41202 17876
rect 42429 17867 42487 17873
rect 42429 17833 42441 17867
rect 42475 17864 42487 17867
rect 42794 17864 42800 17876
rect 42475 17836 42800 17864
rect 42475 17833 42487 17836
rect 42429 17827 42487 17833
rect 42794 17824 42800 17836
rect 42852 17824 42858 17876
rect 44269 17867 44327 17873
rect 42904 17836 43852 17864
rect 28276 17768 33180 17796
rect 24949 17731 25007 17737
rect 24949 17728 24961 17731
rect 24688 17700 24961 17728
rect 24949 17697 24961 17700
rect 24995 17728 25007 17731
rect 27890 17728 27896 17740
rect 24995 17700 27896 17728
rect 24995 17697 25007 17700
rect 24949 17691 25007 17697
rect 27890 17688 27896 17700
rect 27948 17688 27954 17740
rect 21729 17663 21787 17669
rect 21729 17629 21741 17663
rect 21775 17660 21787 17663
rect 24578 17660 24584 17672
rect 21775 17632 24584 17660
rect 21775 17629 21787 17632
rect 21729 17623 21787 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 24854 17620 24860 17672
rect 24912 17660 24918 17672
rect 25041 17663 25099 17669
rect 24912 17632 24957 17660
rect 24912 17620 24918 17632
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 25593 17663 25651 17669
rect 25593 17629 25605 17663
rect 25639 17660 25651 17663
rect 26234 17660 26240 17672
rect 25639 17632 26240 17660
rect 25639 17629 25651 17632
rect 25593 17623 25651 17629
rect 24026 17592 24032 17604
rect 20824 17564 23888 17592
rect 23987 17564 24032 17592
rect 19674 17555 19732 17561
rect 15746 17524 15752 17536
rect 14476 17496 15752 17524
rect 14369 17487 14427 17493
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 16117 17527 16175 17533
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 16574 17524 16580 17536
rect 16163 17496 16580 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 16758 17484 16764 17536
rect 16816 17524 16822 17536
rect 23750 17524 23756 17536
rect 16816 17496 23756 17524
rect 16816 17484 16822 17496
rect 23750 17484 23756 17496
rect 23808 17484 23814 17536
rect 23860 17524 23888 17564
rect 24026 17552 24032 17564
rect 24084 17552 24090 17604
rect 25056 17592 25084 17623
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 26418 17620 26424 17672
rect 26476 17660 26482 17672
rect 28276 17660 28304 17768
rect 41046 17756 41052 17808
rect 41104 17796 41110 17808
rect 42904 17796 42932 17836
rect 41104 17768 42932 17796
rect 43824 17796 43852 17836
rect 44269 17833 44281 17867
rect 44315 17864 44327 17867
rect 44358 17864 44364 17876
rect 44315 17836 44364 17864
rect 44315 17833 44327 17836
rect 44269 17827 44327 17833
rect 44358 17824 44364 17836
rect 44416 17824 44422 17876
rect 45554 17824 45560 17876
rect 45612 17864 45618 17876
rect 45741 17867 45799 17873
rect 45741 17864 45753 17867
rect 45612 17836 45753 17864
rect 45612 17824 45618 17836
rect 45741 17833 45753 17836
rect 45787 17833 45799 17867
rect 51718 17864 51724 17876
rect 45741 17827 45799 17833
rect 47412 17836 51724 17864
rect 43824 17768 47164 17796
rect 41104 17756 41110 17768
rect 29089 17731 29147 17737
rect 29089 17697 29101 17731
rect 29135 17697 29147 17731
rect 29089 17691 29147 17697
rect 26476 17632 28304 17660
rect 26476 17620 26482 17632
rect 28442 17620 28448 17672
rect 28500 17660 28506 17672
rect 28813 17663 28871 17669
rect 28813 17660 28825 17663
rect 28500 17632 28825 17660
rect 28500 17620 28506 17632
rect 28813 17629 28825 17632
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 28902 17620 28908 17672
rect 28960 17660 28966 17672
rect 29104 17660 29132 17691
rect 31754 17688 31760 17740
rect 31812 17728 31818 17740
rect 33689 17731 33747 17737
rect 31812 17700 31857 17728
rect 31812 17688 31818 17700
rect 33689 17697 33701 17731
rect 33735 17728 33747 17731
rect 33735 17700 33824 17728
rect 33735 17697 33747 17700
rect 33689 17691 33747 17697
rect 30282 17660 30288 17672
rect 28960 17632 29132 17660
rect 30243 17632 30288 17660
rect 28960 17620 28966 17632
rect 30282 17620 30288 17632
rect 30340 17620 30346 17672
rect 31294 17620 31300 17672
rect 31352 17660 31358 17672
rect 33318 17660 33324 17672
rect 31352 17632 33324 17660
rect 31352 17620 31358 17632
rect 33318 17620 33324 17632
rect 33376 17660 33382 17672
rect 33505 17663 33563 17669
rect 33505 17660 33517 17663
rect 33376 17632 33517 17660
rect 33376 17620 33382 17632
rect 33505 17629 33517 17632
rect 33551 17629 33563 17663
rect 33505 17623 33563 17629
rect 28994 17592 29000 17604
rect 25056 17564 29000 17592
rect 28994 17552 29000 17564
rect 29052 17552 29058 17604
rect 33796 17592 33824 17700
rect 41064 17700 42932 17728
rect 34882 17660 34888 17672
rect 34843 17632 34888 17660
rect 34882 17620 34888 17632
rect 34940 17620 34946 17672
rect 35897 17663 35955 17669
rect 35897 17629 35909 17663
rect 35943 17660 35955 17663
rect 35986 17660 35992 17672
rect 35943 17632 35992 17660
rect 35943 17629 35955 17632
rect 35897 17623 35955 17629
rect 35986 17620 35992 17632
rect 36044 17660 36050 17672
rect 37458 17660 37464 17672
rect 36044 17632 37464 17660
rect 36044 17620 36050 17632
rect 37458 17620 37464 17632
rect 37516 17660 37522 17672
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37516 17632 37841 17660
rect 37516 17620 37522 17632
rect 37829 17629 37841 17632
rect 37875 17660 37887 17663
rect 38654 17660 38660 17672
rect 37875 17632 38660 17660
rect 37875 17629 37887 17632
rect 37829 17623 37887 17629
rect 38654 17620 38660 17632
rect 38712 17660 38718 17672
rect 40037 17663 40095 17669
rect 40037 17660 40049 17663
rect 38712 17632 40049 17660
rect 38712 17620 38718 17632
rect 40037 17629 40049 17632
rect 40083 17660 40095 17663
rect 40586 17660 40592 17672
rect 40083 17632 40592 17660
rect 40083 17629 40095 17632
rect 40037 17623 40095 17629
rect 40586 17620 40592 17632
rect 40644 17660 40650 17672
rect 41064 17660 41092 17700
rect 42904 17672 42932 17700
rect 45388 17700 47072 17728
rect 40644 17632 41092 17660
rect 42153 17663 42211 17669
rect 40644 17620 40650 17632
rect 42153 17629 42165 17663
rect 42199 17629 42211 17663
rect 42153 17623 42211 17629
rect 42245 17663 42303 17669
rect 42245 17629 42257 17663
rect 42291 17662 42303 17663
rect 42291 17660 42380 17662
rect 42886 17660 42892 17672
rect 42291 17634 42748 17660
rect 42291 17629 42303 17634
rect 42352 17632 42748 17634
rect 42847 17632 42892 17660
rect 42245 17623 42303 17629
rect 33152 17564 33824 17592
rect 26878 17524 26884 17536
rect 23860 17496 26884 17524
rect 26878 17484 26884 17496
rect 26936 17484 26942 17536
rect 27614 17484 27620 17536
rect 27672 17524 27678 17536
rect 28166 17524 28172 17536
rect 27672 17496 28172 17524
rect 27672 17484 27678 17496
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 28905 17527 28963 17533
rect 28905 17524 28917 17527
rect 28868 17496 28917 17524
rect 28868 17484 28874 17496
rect 28905 17493 28917 17496
rect 28951 17493 28963 17527
rect 28905 17487 28963 17493
rect 29362 17484 29368 17536
rect 29420 17524 29426 17536
rect 33152 17524 33180 17564
rect 33410 17524 33416 17536
rect 29420 17496 33180 17524
rect 33323 17496 33416 17524
rect 29420 17484 29426 17496
rect 33410 17484 33416 17496
rect 33468 17524 33474 17536
rect 33686 17524 33692 17536
rect 33468 17496 33692 17524
rect 33468 17484 33474 17496
rect 33686 17484 33692 17496
rect 33744 17484 33750 17536
rect 33796 17524 33824 17564
rect 34422 17552 34428 17604
rect 34480 17592 34486 17604
rect 35161 17595 35219 17601
rect 35161 17592 35173 17595
rect 34480 17564 35173 17592
rect 34480 17552 34486 17564
rect 35161 17561 35173 17564
rect 35207 17561 35219 17595
rect 35161 17555 35219 17561
rect 36164 17595 36222 17601
rect 36164 17561 36176 17595
rect 36210 17592 36222 17595
rect 36814 17592 36820 17604
rect 36210 17564 36820 17592
rect 36210 17561 36222 17564
rect 36164 17555 36222 17561
rect 36814 17552 36820 17564
rect 36872 17552 36878 17604
rect 37366 17592 37372 17604
rect 36924 17564 37372 17592
rect 36924 17524 36952 17564
rect 37366 17552 37372 17564
rect 37424 17552 37430 17604
rect 38096 17595 38154 17601
rect 38096 17561 38108 17595
rect 38142 17592 38154 17595
rect 38562 17592 38568 17604
rect 38142 17564 38568 17592
rect 38142 17561 38154 17564
rect 38096 17555 38154 17561
rect 38562 17552 38568 17564
rect 38620 17552 38626 17604
rect 40304 17595 40362 17601
rect 40304 17561 40316 17595
rect 40350 17592 40362 17595
rect 41782 17592 41788 17604
rect 40350 17564 41788 17592
rect 40350 17561 40362 17564
rect 40304 17555 40362 17561
rect 41782 17552 41788 17564
rect 41840 17552 41846 17604
rect 42168 17592 42196 17623
rect 42610 17592 42616 17604
rect 42168 17564 42616 17592
rect 42610 17552 42616 17564
rect 42668 17552 42674 17604
rect 42720 17592 42748 17632
rect 42886 17620 42892 17632
rect 42944 17620 42950 17672
rect 44082 17620 44088 17672
rect 44140 17660 44146 17672
rect 45189 17663 45247 17669
rect 45189 17660 45201 17663
rect 44140 17632 45201 17660
rect 44140 17620 44146 17632
rect 45189 17629 45201 17632
rect 45235 17629 45247 17663
rect 45189 17623 45247 17629
rect 42978 17592 42984 17604
rect 42720 17564 42984 17592
rect 42978 17552 42984 17564
rect 43036 17552 43042 17604
rect 43162 17601 43168 17604
rect 43156 17555 43168 17601
rect 43220 17592 43226 17604
rect 43220 17564 43256 17592
rect 43162 17552 43168 17555
rect 43220 17552 43226 17564
rect 44450 17552 44456 17604
rect 44508 17592 44514 17604
rect 45388 17601 45416 17700
rect 45554 17660 45560 17672
rect 45515 17632 45560 17660
rect 45554 17620 45560 17632
rect 45612 17620 45618 17672
rect 45373 17595 45431 17601
rect 45373 17592 45385 17595
rect 44508 17564 45385 17592
rect 44508 17552 44514 17564
rect 45373 17561 45385 17564
rect 45419 17561 45431 17595
rect 45373 17555 45431 17561
rect 45465 17595 45523 17601
rect 45465 17561 45477 17595
rect 45511 17592 45523 17595
rect 46750 17592 46756 17604
rect 45511 17564 46756 17592
rect 45511 17561 45523 17564
rect 45465 17555 45523 17561
rect 46750 17552 46756 17564
rect 46808 17552 46814 17604
rect 47044 17592 47072 17700
rect 47136 17669 47164 17768
rect 47412 17669 47440 17836
rect 51718 17824 51724 17836
rect 51776 17824 51782 17876
rect 48130 17728 48136 17740
rect 48091 17700 48136 17728
rect 48130 17688 48136 17700
rect 48188 17688 48194 17740
rect 47121 17663 47179 17669
rect 47121 17629 47133 17663
rect 47167 17629 47179 17663
rect 47121 17623 47179 17629
rect 47397 17663 47455 17669
rect 47397 17629 47409 17663
rect 47443 17629 47455 17663
rect 47397 17623 47455 17629
rect 47486 17620 47492 17672
rect 47544 17660 47550 17672
rect 48148 17660 48176 17688
rect 50341 17663 50399 17669
rect 50341 17660 50353 17663
rect 47544 17632 47589 17660
rect 48148 17632 50353 17660
rect 47544 17620 47550 17632
rect 50341 17629 50353 17632
rect 50387 17629 50399 17663
rect 50341 17623 50399 17629
rect 47305 17595 47363 17601
rect 47305 17592 47317 17595
rect 47044 17564 47317 17592
rect 47305 17561 47317 17564
rect 47351 17592 47363 17595
rect 48038 17592 48044 17604
rect 47351 17564 48044 17592
rect 47351 17561 47363 17564
rect 47305 17555 47363 17561
rect 48038 17552 48044 17564
rect 48096 17552 48102 17604
rect 48400 17595 48458 17601
rect 48400 17561 48412 17595
rect 48446 17592 48458 17595
rect 48498 17592 48504 17604
rect 48446 17564 48504 17592
rect 48446 17561 48458 17564
rect 48400 17555 48458 17561
rect 48498 17552 48504 17564
rect 48556 17552 48562 17604
rect 48590 17552 48596 17604
rect 48648 17592 48654 17604
rect 48648 17564 49556 17592
rect 48648 17552 48654 17564
rect 37274 17524 37280 17536
rect 33796 17496 36952 17524
rect 37235 17496 37280 17524
rect 37274 17484 37280 17496
rect 37332 17484 37338 17536
rect 37642 17484 37648 17536
rect 37700 17524 37706 17536
rect 39022 17524 39028 17536
rect 37700 17496 39028 17524
rect 37700 17484 37706 17496
rect 39022 17484 39028 17496
rect 39080 17484 39086 17536
rect 39206 17524 39212 17536
rect 39167 17496 39212 17524
rect 39206 17484 39212 17496
rect 39264 17484 39270 17536
rect 40586 17484 40592 17536
rect 40644 17524 40650 17536
rect 41417 17527 41475 17533
rect 41417 17524 41429 17527
rect 40644 17496 41429 17524
rect 40644 17484 40650 17496
rect 41417 17493 41429 17496
rect 41463 17493 41475 17527
rect 41417 17487 41475 17493
rect 41690 17484 41696 17536
rect 41748 17524 41754 17536
rect 46290 17524 46296 17536
rect 41748 17496 46296 17524
rect 41748 17484 41754 17496
rect 46290 17484 46296 17496
rect 46348 17484 46354 17536
rect 47673 17527 47731 17533
rect 47673 17493 47685 17527
rect 47719 17524 47731 17527
rect 49234 17524 49240 17536
rect 47719 17496 49240 17524
rect 47719 17493 47731 17496
rect 47673 17487 47731 17493
rect 49234 17484 49240 17496
rect 49292 17484 49298 17536
rect 49528 17533 49556 17564
rect 49970 17552 49976 17604
rect 50028 17592 50034 17604
rect 50586 17595 50644 17601
rect 50586 17592 50598 17595
rect 50028 17564 50598 17592
rect 50028 17552 50034 17564
rect 50586 17561 50598 17564
rect 50632 17561 50644 17595
rect 50586 17555 50644 17561
rect 49513 17527 49571 17533
rect 49513 17493 49525 17527
rect 49559 17493 49571 17527
rect 49513 17487 49571 17493
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 15252 17292 20361 17320
rect 15252 17280 15258 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 21174 17280 21180 17332
rect 21232 17320 21238 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 21232 17292 22385 17320
rect 21232 17280 21238 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 24118 17320 24124 17332
rect 24079 17292 24124 17320
rect 22373 17283 22431 17289
rect 24118 17280 24124 17292
rect 24176 17280 24182 17332
rect 25774 17280 25780 17332
rect 25832 17320 25838 17332
rect 25869 17323 25927 17329
rect 25869 17320 25881 17323
rect 25832 17292 25881 17320
rect 25832 17280 25838 17292
rect 25869 17289 25881 17292
rect 25915 17289 25927 17323
rect 26237 17323 26295 17329
rect 26237 17320 26249 17323
rect 25869 17283 25927 17289
rect 25976 17292 26249 17320
rect 3694 17212 3700 17264
rect 3752 17252 3758 17264
rect 13722 17252 13728 17264
rect 3752 17224 13728 17252
rect 3752 17212 3758 17224
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 17580 17255 17638 17261
rect 17580 17221 17592 17255
rect 17626 17252 17638 17255
rect 17626 17224 19564 17252
rect 17626 17221 17638 17224
rect 17580 17215 17638 17221
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 1627 17156 2452 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2424 16989 2452 17156
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13872 17156 14013 17184
rect 13872 17144 13878 17156
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 19153 17187 19211 17193
rect 19153 17184 19165 17187
rect 18656 17156 19165 17184
rect 18656 17144 18662 17156
rect 19153 17153 19165 17156
rect 19199 17153 19211 17187
rect 19536 17184 19564 17224
rect 19610 17212 19616 17264
rect 19668 17252 19674 17264
rect 19668 17224 22968 17252
rect 19668 17212 19674 17224
rect 20530 17184 20536 17196
rect 19536 17156 20536 17184
rect 19153 17147 19211 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20640 17156 22140 17184
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 17218 17116 17224 17128
rect 16908 17088 17224 17116
rect 16908 17076 16914 17088
rect 17218 17076 17224 17088
rect 17276 17116 17282 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 17276 17088 17325 17116
rect 17276 17076 17282 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 18414 17076 18420 17128
rect 18472 17116 18478 17128
rect 18874 17116 18880 17128
rect 18472 17088 18880 17116
rect 18472 17076 18478 17088
rect 18874 17076 18880 17088
rect 18932 17076 18938 17128
rect 19610 17116 19616 17128
rect 19168 17088 19616 17116
rect 18598 17008 18604 17060
rect 18656 17048 18662 17060
rect 18693 17051 18751 17057
rect 18693 17048 18705 17051
rect 18656 17020 18705 17048
rect 18656 17008 18662 17020
rect 18693 17017 18705 17020
rect 18739 17048 18751 17051
rect 19168 17048 19196 17088
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 20162 17076 20168 17128
rect 20220 17116 20226 17128
rect 20640 17116 20668 17156
rect 20220 17088 20668 17116
rect 20220 17076 20226 17088
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21358 17116 21364 17128
rect 20772 17088 21364 17116
rect 20772 17076 20778 17088
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 21910 17076 21916 17128
rect 21968 17116 21974 17128
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21968 17088 22017 17116
rect 21968 17076 21974 17088
rect 22005 17085 22017 17088
rect 22051 17085 22063 17119
rect 22112 17116 22140 17156
rect 22186 17144 22192 17196
rect 22244 17184 22250 17196
rect 22940 17193 22968 17224
rect 24486 17212 24492 17264
rect 24544 17252 24550 17264
rect 25682 17252 25688 17264
rect 24544 17224 25688 17252
rect 24544 17212 24550 17224
rect 25682 17212 25688 17224
rect 25740 17212 25746 17264
rect 22925 17187 22983 17193
rect 22244 17156 22289 17184
rect 22244 17144 22250 17156
rect 22925 17153 22937 17187
rect 22971 17184 22983 17187
rect 25976 17184 26004 17292
rect 26237 17289 26249 17292
rect 26283 17320 26295 17323
rect 27430 17320 27436 17332
rect 26283 17292 27436 17320
rect 26283 17289 26295 17292
rect 26237 17283 26295 17289
rect 27430 17280 27436 17292
rect 27488 17280 27494 17332
rect 27525 17323 27583 17329
rect 27525 17289 27537 17323
rect 27571 17320 27583 17323
rect 29822 17320 29828 17332
rect 27571 17292 29828 17320
rect 27571 17289 27583 17292
rect 27525 17283 27583 17289
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 30282 17280 30288 17332
rect 30340 17320 30346 17332
rect 33781 17323 33839 17329
rect 33781 17320 33793 17323
rect 30340 17292 33793 17320
rect 30340 17280 30346 17292
rect 33781 17289 33793 17292
rect 33827 17289 33839 17323
rect 33781 17283 33839 17289
rect 34790 17280 34796 17332
rect 34848 17320 34854 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 34848 17292 37841 17320
rect 34848 17280 34854 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 38654 17320 38660 17332
rect 37829 17283 37887 17289
rect 38396 17292 38660 17320
rect 33502 17252 33508 17264
rect 22971 17156 26004 17184
rect 26059 17224 27936 17252
rect 22971 17153 22983 17156
rect 22925 17147 22983 17153
rect 26059 17116 26087 17224
rect 26326 17144 26332 17196
rect 26384 17184 26390 17196
rect 27062 17184 27068 17196
rect 26384 17156 27068 17184
rect 26384 17144 26390 17156
rect 27062 17144 27068 17156
rect 27120 17144 27126 17196
rect 27338 17184 27344 17196
rect 27299 17156 27344 17184
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 22112 17088 26087 17116
rect 26513 17119 26571 17125
rect 22005 17079 22063 17085
rect 26513 17085 26525 17119
rect 26559 17116 26571 17119
rect 26694 17116 26700 17128
rect 26559 17088 26700 17116
rect 26559 17085 26571 17088
rect 26513 17079 26571 17085
rect 20898 17048 20904 17060
rect 18739 17020 19196 17048
rect 19306 17020 20904 17048
rect 18739 17017 18751 17020
rect 18693 17011 18751 17017
rect 2409 16983 2467 16989
rect 2409 16949 2421 16983
rect 2455 16980 2467 16983
rect 14918 16980 14924 16992
rect 2455 16952 14924 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 15378 16980 15384 16992
rect 15339 16952 15384 16980
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 19306 16980 19334 17020
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 22020 17048 22048 17079
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27614 17116 27620 17128
rect 27203 17088 27620 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 27908 17116 27936 17224
rect 28966 17224 33508 17252
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 28966 17184 28994 17224
rect 33502 17212 33508 17224
rect 33560 17212 33566 17264
rect 33686 17212 33692 17264
rect 33744 17252 33750 17264
rect 35713 17255 35771 17261
rect 35713 17252 35725 17255
rect 33744 17224 35725 17252
rect 33744 17212 33750 17224
rect 35713 17221 35725 17224
rect 35759 17221 35771 17255
rect 35713 17215 35771 17221
rect 35897 17255 35955 17261
rect 35897 17221 35909 17255
rect 35943 17221 35955 17255
rect 35897 17215 35955 17221
rect 28031 17156 28994 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 31294 17144 31300 17196
rect 31352 17187 31358 17196
rect 31389 17187 31447 17193
rect 31352 17159 31401 17187
rect 31352 17144 31358 17159
rect 31389 17153 31401 17159
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 31481 17187 31539 17193
rect 31481 17153 31493 17187
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 32585 17187 32643 17193
rect 32585 17153 32597 17187
rect 32631 17184 32643 17187
rect 32674 17184 32680 17196
rect 32631 17156 32680 17184
rect 32631 17153 32643 17156
rect 32585 17147 32643 17153
rect 31202 17116 31208 17128
rect 27908 17088 31208 17116
rect 31202 17076 31208 17088
rect 31260 17116 31266 17128
rect 31496 17116 31524 17147
rect 32674 17144 32680 17156
rect 32732 17144 32738 17196
rect 35912 17184 35940 17215
rect 33796 17156 35940 17184
rect 31260 17088 31524 17116
rect 31260 17076 31266 17088
rect 31570 17076 31576 17128
rect 31628 17116 31634 17128
rect 31628 17088 31673 17116
rect 31628 17076 31634 17088
rect 23106 17048 23112 17060
rect 22020 17020 23112 17048
rect 23106 17008 23112 17020
rect 23164 17008 23170 17060
rect 23750 17008 23756 17060
rect 23808 17048 23814 17060
rect 33796 17048 33824 17156
rect 36078 17144 36084 17196
rect 36136 17184 36142 17196
rect 36725 17187 36783 17193
rect 36725 17184 36737 17187
rect 36136 17156 36737 17184
rect 36136 17144 36142 17156
rect 36725 17153 36737 17156
rect 36771 17153 36783 17187
rect 36725 17147 36783 17153
rect 37182 17144 37188 17196
rect 37240 17184 37246 17196
rect 37461 17187 37519 17193
rect 37461 17184 37473 17187
rect 37240 17156 37473 17184
rect 37240 17144 37246 17156
rect 37461 17153 37473 17156
rect 37507 17153 37519 17187
rect 37642 17184 37648 17196
rect 37603 17156 37648 17184
rect 37461 17147 37519 17153
rect 37642 17144 37648 17156
rect 37700 17144 37706 17196
rect 38396 17193 38424 17292
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 39761 17323 39819 17329
rect 39761 17289 39773 17323
rect 39807 17320 39819 17323
rect 39850 17320 39856 17332
rect 39807 17292 39856 17320
rect 39807 17289 39819 17292
rect 39761 17283 39819 17289
rect 39850 17280 39856 17292
rect 39908 17280 39914 17332
rect 40586 17280 40592 17332
rect 40644 17320 40650 17332
rect 40681 17323 40739 17329
rect 40681 17320 40693 17323
rect 40644 17292 40693 17320
rect 40644 17280 40650 17292
rect 40681 17289 40693 17292
rect 40727 17289 40739 17323
rect 40681 17283 40739 17289
rect 41138 17280 41144 17332
rect 41196 17320 41202 17332
rect 42150 17320 42156 17332
rect 41196 17292 42156 17320
rect 41196 17280 41202 17292
rect 42150 17280 42156 17292
rect 42208 17280 42214 17332
rect 43622 17280 43628 17332
rect 43680 17320 43686 17332
rect 45557 17323 45615 17329
rect 45557 17320 45569 17323
rect 43680 17292 45569 17320
rect 43680 17280 43686 17292
rect 45557 17289 45569 17292
rect 45603 17320 45615 17323
rect 45646 17320 45652 17332
rect 45603 17292 45652 17320
rect 45603 17289 45615 17292
rect 45557 17283 45615 17289
rect 45646 17280 45652 17292
rect 45704 17280 45710 17332
rect 49878 17320 49884 17332
rect 49839 17292 49884 17320
rect 49878 17280 49884 17292
rect 49936 17280 49942 17332
rect 41877 17255 41935 17261
rect 41877 17252 41889 17255
rect 40052 17224 41889 17252
rect 38381 17187 38439 17193
rect 38381 17153 38393 17187
rect 38427 17153 38439 17187
rect 38381 17147 38439 17153
rect 38648 17187 38706 17193
rect 38648 17153 38660 17187
rect 38694 17184 38706 17187
rect 40052 17184 40080 17224
rect 41877 17221 41889 17224
rect 41923 17221 41935 17255
rect 41877 17215 41935 17221
rect 42981 17255 43039 17261
rect 42981 17221 42993 17255
rect 43027 17252 43039 17255
rect 44358 17252 44364 17264
rect 43027 17224 44364 17252
rect 43027 17221 43039 17224
rect 42981 17215 43039 17221
rect 44358 17212 44364 17224
rect 44416 17212 44422 17264
rect 48768 17255 48826 17261
rect 48768 17221 48780 17255
rect 48814 17252 48826 17255
rect 49694 17252 49700 17264
rect 48814 17224 49700 17252
rect 48814 17221 48826 17224
rect 48768 17215 48826 17221
rect 49694 17212 49700 17224
rect 49752 17212 49758 17264
rect 38694 17156 40080 17184
rect 38694 17153 38706 17156
rect 38648 17147 38706 17153
rect 40218 17144 40224 17196
rect 40276 17184 40282 17196
rect 40773 17187 40831 17193
rect 40773 17184 40785 17187
rect 40276 17156 40785 17184
rect 40276 17144 40282 17156
rect 40773 17153 40785 17156
rect 40819 17153 40831 17187
rect 41693 17187 41751 17193
rect 41693 17184 41705 17187
rect 40773 17147 40831 17153
rect 40871 17156 41705 17184
rect 33962 17076 33968 17128
rect 34020 17116 34026 17128
rect 35989 17119 36047 17125
rect 35989 17116 36001 17119
rect 34020 17088 36001 17116
rect 34020 17076 34026 17088
rect 35989 17085 36001 17088
rect 36035 17116 36047 17119
rect 36354 17116 36360 17128
rect 36035 17088 36360 17116
rect 36035 17085 36047 17088
rect 35989 17079 36047 17085
rect 36354 17076 36360 17088
rect 36412 17076 36418 17128
rect 36538 17116 36544 17128
rect 36499 17088 36544 17116
rect 36538 17076 36544 17088
rect 36596 17076 36602 17128
rect 39942 17076 39948 17128
rect 40000 17116 40006 17128
rect 40871 17116 40899 17156
rect 41693 17153 41705 17156
rect 41739 17153 41751 17187
rect 41693 17147 41751 17153
rect 42705 17187 42763 17193
rect 42705 17153 42717 17187
rect 42751 17153 42763 17187
rect 42705 17147 42763 17153
rect 42889 17187 42947 17193
rect 42889 17153 42901 17187
rect 42935 17153 42947 17187
rect 42889 17147 42947 17153
rect 43073 17187 43131 17193
rect 43073 17153 43085 17187
rect 43119 17184 43131 17187
rect 43806 17184 43812 17196
rect 43119 17156 43812 17184
rect 43119 17153 43131 17156
rect 43073 17147 43131 17153
rect 40000 17088 40899 17116
rect 40957 17119 41015 17125
rect 40000 17076 40006 17088
rect 40957 17085 40969 17119
rect 41003 17116 41015 17119
rect 41003 17088 41184 17116
rect 41003 17085 41015 17088
rect 40957 17079 41015 17085
rect 41046 17048 41052 17060
rect 23808 17020 33824 17048
rect 36832 17020 38424 17048
rect 23808 17008 23814 17020
rect 16724 16952 19334 16980
rect 16724 16940 16730 16952
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20806 16980 20812 16992
rect 19852 16952 20812 16980
rect 19852 16940 19858 16952
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 24118 16940 24124 16992
rect 24176 16980 24182 16992
rect 24762 16980 24768 16992
rect 24176 16952 24768 16980
rect 24176 16940 24182 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 25682 16940 25688 16992
rect 25740 16980 25746 16992
rect 29181 16983 29239 16989
rect 29181 16980 29193 16983
rect 25740 16952 29193 16980
rect 25740 16940 25746 16952
rect 29181 16949 29193 16952
rect 29227 16949 29239 16983
rect 29181 16943 29239 16949
rect 30282 16940 30288 16992
rect 30340 16980 30346 16992
rect 30742 16980 30748 16992
rect 30340 16952 30748 16980
rect 30340 16940 30346 16952
rect 30742 16940 30748 16952
rect 30800 16940 30806 16992
rect 31021 16983 31079 16989
rect 31021 16949 31033 16983
rect 31067 16980 31079 16983
rect 32398 16980 32404 16992
rect 31067 16952 32404 16980
rect 31067 16949 31079 16952
rect 31021 16943 31079 16949
rect 32398 16940 32404 16952
rect 32456 16940 32462 16992
rect 35437 16983 35495 16989
rect 35437 16949 35449 16983
rect 35483 16980 35495 16983
rect 36832 16980 36860 17020
rect 35483 16952 36860 16980
rect 35483 16949 35495 16952
rect 35437 16943 35495 16949
rect 36906 16940 36912 16992
rect 36964 16980 36970 16992
rect 36964 16952 37009 16980
rect 36964 16940 36970 16952
rect 37826 16940 37832 16992
rect 37884 16980 37890 16992
rect 38286 16980 38292 16992
rect 37884 16952 38292 16980
rect 37884 16940 37890 16952
rect 38286 16940 38292 16952
rect 38344 16940 38350 16992
rect 38396 16980 38424 17020
rect 40144 17020 41052 17048
rect 40144 16980 40172 17020
rect 41046 17008 41052 17020
rect 41104 17008 41110 17060
rect 40310 16980 40316 16992
rect 38396 16952 40172 16980
rect 40271 16952 40316 16980
rect 40310 16940 40316 16952
rect 40368 16940 40374 16992
rect 40402 16940 40408 16992
rect 40460 16980 40466 16992
rect 41156 16980 41184 17088
rect 41414 17076 41420 17128
rect 41472 17116 41478 17128
rect 41509 17119 41567 17125
rect 41509 17116 41521 17119
rect 41472 17088 41521 17116
rect 41472 17076 41478 17088
rect 41509 17085 41521 17088
rect 41555 17085 41567 17119
rect 41509 17079 41567 17085
rect 40460 16952 41184 16980
rect 40460 16940 40466 16952
rect 41506 16940 41512 16992
rect 41564 16980 41570 16992
rect 42720 16980 42748 17147
rect 42904 17116 42932 17147
rect 43806 17144 43812 17156
rect 43864 17184 43870 17196
rect 43990 17184 43996 17196
rect 43864 17156 43996 17184
rect 43864 17144 43870 17156
rect 43990 17144 43996 17156
rect 44048 17144 44054 17196
rect 44444 17187 44502 17193
rect 44444 17153 44456 17187
rect 44490 17184 44502 17187
rect 45554 17184 45560 17196
rect 44490 17156 45560 17184
rect 44490 17153 44502 17156
rect 44444 17147 44502 17153
rect 45554 17144 45560 17156
rect 45612 17144 45618 17196
rect 42978 17116 42984 17128
rect 42904 17088 42984 17116
rect 42978 17076 42984 17088
rect 43036 17076 43042 17128
rect 44174 17116 44180 17128
rect 44135 17088 44180 17116
rect 44174 17076 44180 17088
rect 44232 17076 44238 17128
rect 48130 17076 48136 17128
rect 48188 17116 48194 17128
rect 48501 17119 48559 17125
rect 48501 17116 48513 17119
rect 48188 17088 48513 17116
rect 48188 17076 48194 17088
rect 48501 17085 48513 17088
rect 48547 17085 48559 17119
rect 48501 17079 48559 17085
rect 43254 16980 43260 16992
rect 41564 16952 42748 16980
rect 43215 16952 43260 16980
rect 41564 16940 41570 16952
rect 43254 16940 43260 16952
rect 43312 16940 43318 16992
rect 43990 16940 43996 16992
rect 44048 16980 44054 16992
rect 45462 16980 45468 16992
rect 44048 16952 45468 16980
rect 44048 16940 44054 16952
rect 45462 16940 45468 16952
rect 45520 16940 45526 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 30374 16776 30380 16788
rect 13464 16748 30380 16776
rect 13464 16649 13492 16748
rect 30374 16736 30380 16748
rect 30432 16736 30438 16788
rect 30834 16736 30840 16788
rect 30892 16776 30898 16788
rect 36078 16776 36084 16788
rect 30892 16748 36084 16776
rect 30892 16736 30898 16748
rect 36078 16736 36084 16748
rect 36136 16736 36142 16788
rect 57149 16779 57207 16785
rect 57149 16776 57161 16779
rect 37568 16748 57161 16776
rect 15565 16711 15623 16717
rect 15565 16677 15577 16711
rect 15611 16708 15623 16711
rect 16758 16708 16764 16720
rect 15611 16680 16764 16708
rect 15611 16677 15623 16680
rect 15565 16671 15623 16677
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 25961 16711 26019 16717
rect 25961 16677 25973 16711
rect 26007 16677 26019 16711
rect 25961 16671 26019 16677
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 14826 16640 14832 16652
rect 14787 16612 14832 16640
rect 13449 16603 13507 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 16206 16640 16212 16652
rect 15151 16612 16212 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 19794 16640 19800 16652
rect 16500 16612 19800 16640
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13357 16575 13415 16581
rect 13357 16572 13369 16575
rect 13228 16544 13369 16572
rect 13228 16532 13234 16544
rect 13357 16541 13369 16544
rect 13403 16541 13415 16575
rect 13538 16572 13544 16584
rect 13499 16544 13544 16572
rect 13357 16535 13415 16541
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 14737 16575 14795 16581
rect 13688 16544 13733 16572
rect 13688 16532 13694 16544
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 15930 16572 15936 16584
rect 15891 16544 15936 16572
rect 14737 16535 14795 16541
rect 1854 16504 1860 16516
rect 1815 16476 1860 16504
rect 1854 16464 1860 16476
rect 1912 16464 1918 16516
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 14752 16504 14780 16535
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16500 16572 16528 16612
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 23032 16612 23336 16640
rect 16163 16544 16528 16572
rect 16577 16575 16635 16581
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16577 16541 16589 16575
rect 16623 16569 16635 16575
rect 18046 16572 18052 16584
rect 16684 16569 18052 16572
rect 16623 16544 18052 16569
rect 16623 16541 16712 16544
rect 16577 16535 16635 16541
rect 18046 16532 18052 16544
rect 18104 16532 18110 16584
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18840 16544 18889 16572
rect 18840 16532 18846 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 19484 16544 19901 16572
rect 19484 16532 19490 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 21729 16575 21787 16581
rect 21729 16572 21741 16575
rect 20680 16544 21741 16572
rect 20680 16532 20686 16544
rect 21729 16541 21741 16544
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 12400 16476 14780 16504
rect 15841 16507 15899 16513
rect 12400 16464 12406 16476
rect 15841 16473 15853 16507
rect 15887 16504 15899 16507
rect 18598 16504 18604 16516
rect 15887 16476 18604 16504
rect 15887 16473 15899 16476
rect 15841 16467 15899 16473
rect 18598 16464 18604 16476
rect 18656 16464 18662 16516
rect 20156 16507 20214 16513
rect 20156 16473 20168 16507
rect 20202 16504 20214 16507
rect 23032 16504 23060 16612
rect 23106 16532 23112 16584
rect 23164 16572 23170 16584
rect 23308 16572 23336 16612
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 24581 16643 24639 16649
rect 24581 16640 24593 16643
rect 23440 16612 24593 16640
rect 23440 16600 23446 16612
rect 24581 16609 24593 16612
rect 24627 16609 24639 16643
rect 24581 16603 24639 16609
rect 23164 16544 23244 16572
rect 23308 16544 23428 16572
rect 23164 16532 23170 16544
rect 20202 16476 23060 16504
rect 20202 16473 20214 16476
rect 20156 16467 20214 16473
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 11112 16408 13185 16436
rect 11112 16396 11118 16408
rect 13173 16405 13185 16408
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 18322 16436 18328 16448
rect 15795 16408 18328 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16436 21327 16439
rect 22922 16436 22928 16448
rect 21315 16408 22928 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 23106 16436 23112 16448
rect 23067 16408 23112 16436
rect 23106 16396 23112 16408
rect 23164 16396 23170 16448
rect 23216 16436 23244 16544
rect 23400 16504 23428 16544
rect 24026 16532 24032 16584
rect 24084 16572 24090 16584
rect 24837 16575 24895 16581
rect 24837 16572 24849 16575
rect 24084 16544 24849 16572
rect 24084 16532 24090 16544
rect 24837 16541 24849 16544
rect 24883 16541 24895 16575
rect 25976 16572 26004 16671
rect 26050 16668 26056 16720
rect 26108 16708 26114 16720
rect 26694 16708 26700 16720
rect 26108 16680 26700 16708
rect 26108 16668 26114 16680
rect 26694 16668 26700 16680
rect 26752 16708 26758 16720
rect 29362 16708 29368 16720
rect 26752 16680 29368 16708
rect 26752 16668 26758 16680
rect 29362 16668 29368 16680
rect 29420 16668 29426 16720
rect 32674 16668 32680 16720
rect 32732 16708 32738 16720
rect 34974 16708 34980 16720
rect 32732 16680 34980 16708
rect 32732 16668 32738 16680
rect 34974 16668 34980 16680
rect 35032 16668 35038 16720
rect 37568 16708 37596 16748
rect 57149 16745 57161 16748
rect 57195 16745 57207 16779
rect 57149 16739 57207 16745
rect 35360 16680 36124 16708
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 28718 16640 28724 16652
rect 27672 16612 28724 16640
rect 27672 16600 27678 16612
rect 28718 16600 28724 16612
rect 28776 16600 28782 16652
rect 29730 16640 29736 16652
rect 29691 16612 29736 16640
rect 29730 16600 29736 16612
rect 29788 16600 29794 16652
rect 30742 16600 30748 16652
rect 30800 16640 30806 16652
rect 35360 16640 35388 16680
rect 30800 16612 35388 16640
rect 35529 16643 35587 16649
rect 30800 16600 30806 16612
rect 35529 16609 35541 16643
rect 35575 16640 35587 16643
rect 35710 16640 35716 16652
rect 35575 16612 35716 16640
rect 35575 16609 35587 16612
rect 35529 16603 35587 16609
rect 35710 16600 35716 16612
rect 35768 16600 35774 16652
rect 26878 16572 26884 16584
rect 25976 16544 26740 16572
rect 26839 16544 26884 16572
rect 24837 16535 24895 16541
rect 25038 16504 25044 16516
rect 23400 16476 25044 16504
rect 25038 16464 25044 16476
rect 25096 16464 25102 16516
rect 26712 16504 26740 16544
rect 26878 16532 26884 16544
rect 26936 16572 26942 16584
rect 29822 16572 29828 16584
rect 26936 16544 29828 16572
rect 26936 16532 26942 16544
rect 29822 16532 29828 16544
rect 29880 16532 29886 16584
rect 30000 16575 30058 16581
rect 30000 16541 30012 16575
rect 30046 16572 30058 16575
rect 31018 16572 31024 16584
rect 30046 16544 31024 16572
rect 30046 16541 30058 16544
rect 30000 16535 30058 16541
rect 31018 16532 31024 16544
rect 31076 16532 31082 16584
rect 31849 16575 31907 16581
rect 31849 16572 31861 16575
rect 31726 16544 31861 16572
rect 31726 16504 31754 16544
rect 31849 16541 31861 16544
rect 31895 16572 31907 16575
rect 35158 16572 35164 16584
rect 31895 16544 35164 16572
rect 31895 16541 31907 16544
rect 31849 16535 31907 16541
rect 35158 16532 35164 16544
rect 35216 16532 35222 16584
rect 35342 16572 35348 16584
rect 35303 16544 35348 16572
rect 35342 16532 35348 16544
rect 35400 16532 35406 16584
rect 36096 16572 36124 16680
rect 37200 16680 37596 16708
rect 38105 16711 38163 16717
rect 36170 16600 36176 16652
rect 36228 16640 36234 16652
rect 36228 16612 36273 16640
rect 36228 16600 36234 16612
rect 37200 16572 37228 16680
rect 38105 16677 38117 16711
rect 38151 16677 38163 16711
rect 38105 16671 38163 16677
rect 38120 16640 38148 16671
rect 38286 16668 38292 16720
rect 38344 16708 38350 16720
rect 38344 16680 38700 16708
rect 38344 16668 38350 16680
rect 38194 16640 38200 16652
rect 38120 16612 38200 16640
rect 38194 16600 38200 16612
rect 38252 16600 38258 16652
rect 38470 16600 38476 16652
rect 38528 16640 38534 16652
rect 38672 16649 38700 16680
rect 38746 16668 38752 16720
rect 38804 16708 38810 16720
rect 40218 16708 40224 16720
rect 38804 16680 40224 16708
rect 38804 16668 38810 16680
rect 40218 16668 40224 16680
rect 40276 16668 40282 16720
rect 40310 16668 40316 16720
rect 40368 16708 40374 16720
rect 41782 16708 41788 16720
rect 40368 16680 41644 16708
rect 41743 16680 41788 16708
rect 40368 16668 40374 16680
rect 38565 16643 38623 16649
rect 38565 16640 38577 16643
rect 38528 16612 38577 16640
rect 38528 16600 38534 16612
rect 38565 16609 38577 16612
rect 38611 16609 38623 16643
rect 38565 16603 38623 16609
rect 38657 16643 38715 16649
rect 38657 16609 38669 16643
rect 38703 16609 38715 16643
rect 38657 16603 38715 16609
rect 39114 16600 39120 16652
rect 39172 16640 39178 16652
rect 40865 16643 40923 16649
rect 39172 16612 40816 16640
rect 39172 16600 39178 16612
rect 36096 16544 37228 16572
rect 37274 16532 37280 16584
rect 37332 16572 37338 16584
rect 40402 16572 40408 16584
rect 37332 16544 40408 16572
rect 37332 16532 37338 16544
rect 40402 16532 40408 16544
rect 40460 16532 40466 16584
rect 40788 16572 40816 16612
rect 40865 16609 40877 16643
rect 40911 16640 40923 16643
rect 41046 16640 41052 16652
rect 40911 16612 41052 16640
rect 40911 16609 40923 16612
rect 40865 16603 40923 16609
rect 41046 16600 41052 16612
rect 41104 16600 41110 16652
rect 41414 16640 41420 16652
rect 41156 16612 41420 16640
rect 41156 16572 41184 16612
rect 41414 16600 41420 16612
rect 41472 16640 41478 16652
rect 41472 16612 41517 16640
rect 41472 16600 41478 16612
rect 41616 16581 41644 16680
rect 41782 16668 41788 16680
rect 41840 16668 41846 16720
rect 45554 16708 45560 16720
rect 42904 16680 45232 16708
rect 45515 16680 45560 16708
rect 40788 16544 41184 16572
rect 41601 16575 41659 16581
rect 41601 16541 41613 16575
rect 41647 16541 41659 16575
rect 41601 16535 41659 16541
rect 42610 16532 42616 16584
rect 42668 16572 42674 16584
rect 42904 16581 42932 16680
rect 43254 16640 43260 16652
rect 43088 16612 43260 16640
rect 43088 16581 43116 16612
rect 43254 16600 43260 16612
rect 43312 16600 43318 16652
rect 43622 16600 43628 16652
rect 43680 16640 43686 16652
rect 44358 16640 44364 16652
rect 43680 16612 43852 16640
rect 43680 16600 43686 16612
rect 42889 16575 42947 16581
rect 42889 16572 42901 16575
rect 42668 16544 42901 16572
rect 42668 16532 42674 16544
rect 42889 16541 42901 16544
rect 42935 16541 42947 16575
rect 42889 16535 42947 16541
rect 43073 16575 43131 16581
rect 43073 16541 43085 16575
rect 43119 16541 43131 16575
rect 43073 16535 43131 16541
rect 43717 16575 43775 16581
rect 43717 16541 43729 16575
rect 43763 16541 43775 16575
rect 43717 16535 43775 16541
rect 26712 16476 31754 16504
rect 32214 16464 32220 16516
rect 32272 16504 32278 16516
rect 36440 16507 36498 16513
rect 32272 16476 36400 16504
rect 32272 16464 32278 16476
rect 28077 16439 28135 16445
rect 28077 16436 28089 16439
rect 23216 16408 28089 16436
rect 28077 16405 28089 16408
rect 28123 16405 28135 16439
rect 28077 16399 28135 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 29638 16436 29644 16448
rect 28316 16408 29644 16436
rect 28316 16396 28322 16408
rect 29638 16396 29644 16408
rect 29696 16396 29702 16448
rect 31110 16436 31116 16448
rect 31071 16408 31116 16436
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 33042 16436 33048 16448
rect 33003 16408 33048 16436
rect 33042 16396 33048 16408
rect 33100 16396 33106 16448
rect 34698 16396 34704 16448
rect 34756 16436 34762 16448
rect 34885 16439 34943 16445
rect 34885 16436 34897 16439
rect 34756 16408 34897 16436
rect 34756 16396 34762 16408
rect 34885 16405 34897 16408
rect 34931 16405 34943 16439
rect 34885 16399 34943 16405
rect 34974 16396 34980 16448
rect 35032 16436 35038 16448
rect 35253 16439 35311 16445
rect 35253 16436 35265 16439
rect 35032 16408 35265 16436
rect 35032 16396 35038 16408
rect 35253 16405 35265 16408
rect 35299 16436 35311 16439
rect 35618 16436 35624 16448
rect 35299 16408 35624 16436
rect 35299 16405 35311 16408
rect 35253 16399 35311 16405
rect 35618 16396 35624 16408
rect 35676 16396 35682 16448
rect 36372 16436 36400 16476
rect 36440 16473 36452 16507
rect 36486 16504 36498 16507
rect 39758 16504 39764 16516
rect 36486 16476 39764 16504
rect 36486 16473 36498 16476
rect 36440 16467 36498 16473
rect 39758 16464 39764 16476
rect 39816 16464 39822 16516
rect 41506 16504 41512 16516
rect 40236 16476 41512 16504
rect 37553 16439 37611 16445
rect 37553 16436 37565 16439
rect 36372 16408 37565 16436
rect 37553 16405 37565 16408
rect 37599 16436 37611 16439
rect 38473 16439 38531 16445
rect 38473 16436 38485 16439
rect 37599 16408 38485 16436
rect 37599 16405 37611 16408
rect 37553 16399 37611 16405
rect 38473 16405 38485 16408
rect 38519 16436 38531 16439
rect 40126 16436 40132 16448
rect 38519 16408 40132 16436
rect 38519 16405 38531 16408
rect 38473 16399 38531 16405
rect 40126 16396 40132 16408
rect 40184 16396 40190 16448
rect 40236 16445 40264 16476
rect 41506 16464 41512 16476
rect 41564 16464 41570 16516
rect 41708 16476 41920 16504
rect 40221 16439 40279 16445
rect 40221 16405 40233 16439
rect 40267 16405 40279 16439
rect 40586 16436 40592 16448
rect 40547 16408 40592 16436
rect 40221 16399 40279 16405
rect 40586 16396 40592 16408
rect 40644 16396 40650 16448
rect 40681 16439 40739 16445
rect 40681 16405 40693 16439
rect 40727 16436 40739 16439
rect 41138 16436 41144 16448
rect 40727 16408 41144 16436
rect 40727 16405 40739 16408
rect 40681 16399 40739 16405
rect 41138 16396 41144 16408
rect 41196 16396 41202 16448
rect 41322 16396 41328 16448
rect 41380 16436 41386 16448
rect 41708 16436 41736 16476
rect 41380 16408 41736 16436
rect 41892 16436 41920 16476
rect 43162 16464 43168 16516
rect 43220 16504 43226 16516
rect 43257 16507 43315 16513
rect 43257 16504 43269 16507
rect 43220 16476 43269 16504
rect 43220 16464 43226 16476
rect 43257 16473 43269 16476
rect 43303 16473 43315 16507
rect 43257 16467 43315 16473
rect 43732 16436 43760 16535
rect 43824 16504 43852 16612
rect 44008 16612 44364 16640
rect 43901 16575 43959 16581
rect 43901 16541 43913 16575
rect 43947 16572 43959 16575
rect 44008 16572 44036 16612
rect 44358 16600 44364 16612
rect 44416 16600 44422 16652
rect 45204 16649 45232 16680
rect 45554 16668 45560 16680
rect 45612 16668 45618 16720
rect 45189 16643 45247 16649
rect 45189 16609 45201 16643
rect 45235 16609 45247 16643
rect 45189 16603 45247 16609
rect 46842 16600 46848 16652
rect 46900 16640 46906 16652
rect 47489 16643 47547 16649
rect 47489 16640 47501 16643
rect 46900 16612 47501 16640
rect 46900 16600 46906 16612
rect 47489 16609 47501 16612
rect 47535 16609 47547 16643
rect 47489 16603 47547 16609
rect 47857 16643 47915 16649
rect 47857 16609 47869 16643
rect 47903 16640 47915 16643
rect 47903 16612 48084 16640
rect 47903 16609 47915 16612
rect 47857 16603 47915 16609
rect 43947 16544 44036 16572
rect 44085 16575 44143 16581
rect 43947 16541 43959 16544
rect 43901 16535 43959 16541
rect 44085 16541 44097 16575
rect 44131 16572 44143 16575
rect 45373 16575 45431 16581
rect 44131 16544 44211 16572
rect 44131 16541 44143 16544
rect 44085 16535 44143 16541
rect 43993 16507 44051 16513
rect 43993 16504 44005 16507
rect 43824 16476 44005 16504
rect 43993 16473 44005 16476
rect 44039 16473 44051 16507
rect 43993 16467 44051 16473
rect 41892 16408 43760 16436
rect 41380 16396 41386 16408
rect 44082 16396 44088 16448
rect 44140 16436 44146 16448
rect 44183 16436 44211 16544
rect 45373 16541 45385 16575
rect 45419 16541 45431 16575
rect 45373 16535 45431 16541
rect 47673 16575 47731 16581
rect 47673 16541 47685 16575
rect 47719 16541 47731 16575
rect 48056 16572 48084 16612
rect 48130 16600 48136 16652
rect 48188 16640 48194 16652
rect 48317 16643 48375 16649
rect 48317 16640 48329 16643
rect 48188 16612 48329 16640
rect 48188 16600 48194 16612
rect 48317 16609 48329 16612
rect 48363 16609 48375 16643
rect 48317 16603 48375 16609
rect 48573 16575 48631 16581
rect 48573 16572 48585 16575
rect 48056 16544 48585 16572
rect 47673 16535 47731 16541
rect 48573 16541 48585 16544
rect 48619 16541 48631 16575
rect 57885 16575 57943 16581
rect 57885 16572 57897 16575
rect 48573 16535 48631 16541
rect 55186 16544 57897 16572
rect 45388 16504 45416 16535
rect 44284 16476 45416 16504
rect 47688 16504 47716 16535
rect 48682 16504 48688 16516
rect 47688 16476 48688 16504
rect 44284 16445 44312 16476
rect 48682 16464 48688 16476
rect 48740 16464 48746 16516
rect 55186 16504 55214 16544
rect 57885 16541 57897 16544
rect 57931 16541 57943 16575
rect 58158 16572 58164 16584
rect 58119 16544 58164 16572
rect 57885 16535 57943 16541
rect 58158 16532 58164 16544
rect 58216 16532 58222 16584
rect 57054 16504 57060 16516
rect 48792 16476 55214 16504
rect 57015 16476 57060 16504
rect 44140 16408 44211 16436
rect 44269 16439 44327 16445
rect 44140 16396 44146 16408
rect 44269 16405 44281 16439
rect 44315 16405 44327 16439
rect 44269 16399 44327 16405
rect 46750 16396 46756 16448
rect 46808 16436 46814 16448
rect 48792 16436 48820 16476
rect 57054 16464 57060 16476
rect 57112 16464 57118 16516
rect 49694 16436 49700 16448
rect 46808 16408 48820 16436
rect 49607 16408 49700 16436
rect 46808 16396 46814 16408
rect 49694 16396 49700 16408
rect 49752 16436 49758 16448
rect 50798 16436 50804 16448
rect 49752 16408 50804 16436
rect 49752 16396 49758 16408
rect 50798 16396 50804 16408
rect 50856 16396 50862 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 12989 16235 13047 16241
rect 12989 16232 13001 16235
rect 1636 16204 13001 16232
rect 1636 16192 1642 16204
rect 12989 16201 13001 16204
rect 13035 16201 13047 16235
rect 12989 16195 13047 16201
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 24486 16232 24492 16244
rect 13228 16204 24492 16232
rect 13228 16192 13234 16204
rect 24486 16192 24492 16204
rect 24544 16192 24550 16244
rect 25038 16232 25044 16244
rect 24999 16204 25044 16232
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 26878 16192 26884 16244
rect 26936 16232 26942 16244
rect 27982 16232 27988 16244
rect 26936 16204 27988 16232
rect 26936 16192 26942 16204
rect 27982 16192 27988 16204
rect 28040 16232 28046 16244
rect 28997 16235 29055 16241
rect 28997 16232 29009 16235
rect 28040 16204 29009 16232
rect 28040 16192 28046 16204
rect 28997 16201 29009 16204
rect 29043 16201 29055 16235
rect 28997 16195 29055 16201
rect 29270 16192 29276 16244
rect 29328 16232 29334 16244
rect 33042 16232 33048 16244
rect 29328 16204 33048 16232
rect 29328 16192 29334 16204
rect 33042 16192 33048 16204
rect 33100 16192 33106 16244
rect 33686 16232 33692 16244
rect 33647 16204 33692 16232
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 35618 16232 35624 16244
rect 35579 16204 35624 16232
rect 35618 16192 35624 16204
rect 35676 16232 35682 16244
rect 36170 16232 36176 16244
rect 35676 16204 36176 16232
rect 35676 16192 35682 16204
rect 36170 16192 36176 16204
rect 36228 16192 36234 16244
rect 36446 16232 36452 16244
rect 36407 16204 36452 16232
rect 36446 16192 36452 16204
rect 36504 16192 36510 16244
rect 38102 16192 38108 16244
rect 38160 16232 38166 16244
rect 40034 16232 40040 16244
rect 38160 16204 40040 16232
rect 38160 16192 38166 16204
rect 40034 16192 40040 16204
rect 40092 16192 40098 16244
rect 40310 16192 40316 16244
rect 40368 16232 40374 16244
rect 41046 16232 41052 16244
rect 40368 16204 41052 16232
rect 40368 16192 40374 16204
rect 41046 16192 41052 16204
rect 41104 16192 41110 16244
rect 41690 16232 41696 16244
rect 41651 16204 41696 16232
rect 41690 16192 41696 16204
rect 41748 16192 41754 16244
rect 42978 16192 42984 16244
rect 43036 16232 43042 16244
rect 44542 16232 44548 16244
rect 43036 16204 44548 16232
rect 43036 16192 43042 16204
rect 11146 16124 11152 16176
rect 11204 16164 11210 16176
rect 22094 16164 22100 16176
rect 11204 16136 13492 16164
rect 11204 16124 11210 16136
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 12161 16099 12219 16105
rect 1627 16068 2452 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2424 15904 2452 16068
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 13170 16096 13176 16108
rect 12207 16068 13176 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13464 16105 13492 16136
rect 22020 16136 22100 16164
rect 13449 16099 13507 16105
rect 13320 16068 13365 16096
rect 13320 16056 13326 16068
rect 13449 16065 13461 16099
rect 13495 16065 13507 16099
rect 13449 16059 13507 16065
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16096 14059 16099
rect 15102 16096 15108 16108
rect 14047 16068 15108 16096
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 17488 16099 17546 16105
rect 17488 16065 17500 16099
rect 17534 16096 17546 16099
rect 17770 16096 17776 16108
rect 17534 16068 17776 16096
rect 17534 16065 17546 16068
rect 17488 16059 17546 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 22020 16105 22048 16136
rect 22094 16124 22100 16136
rect 22152 16124 22158 16176
rect 22278 16173 22284 16176
rect 22272 16164 22284 16173
rect 22239 16136 22284 16164
rect 22272 16127 22284 16136
rect 22278 16124 22284 16127
rect 22336 16124 22342 16176
rect 22922 16124 22928 16176
rect 22980 16164 22986 16176
rect 27522 16164 27528 16176
rect 22980 16136 27528 16164
rect 22980 16124 22986 16136
rect 27522 16124 27528 16136
rect 27580 16124 27586 16176
rect 27706 16124 27712 16176
rect 27764 16164 27770 16176
rect 27873 16167 27931 16173
rect 27873 16164 27885 16167
rect 27764 16136 27885 16164
rect 27764 16124 27770 16136
rect 27873 16133 27885 16136
rect 27919 16133 27931 16167
rect 27873 16127 27931 16133
rect 29822 16124 29828 16176
rect 29880 16164 29886 16176
rect 32214 16164 32220 16176
rect 29880 16136 32220 16164
rect 29880 16124 29886 16136
rect 32214 16124 32220 16136
rect 32272 16124 32278 16176
rect 32324 16136 33732 16164
rect 32324 16108 32352 16136
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 18288 16068 19165 16096
rect 18288 16056 18294 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 23845 16099 23903 16105
rect 22005 16059 22063 16065
rect 22112 16068 23796 16096
rect 4062 15988 4068 16040
rect 4120 16028 4126 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 4120 16000 11989 16028
rect 4120 15988 4126 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 11977 15991 12035 15997
rect 12084 16000 12265 16028
rect 2406 15892 2412 15904
rect 2367 15864 2412 15892
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 12084 15892 12112 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 12345 16031 12403 16037
rect 12345 15997 12357 16031
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 12158 15920 12164 15972
rect 12216 15960 12222 15972
rect 12360 15960 12388 15991
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 12492 16000 12537 16028
rect 12636 16000 13369 16028
rect 12492 15988 12498 16000
rect 12636 15960 12664 16000
rect 13357 15997 13369 16000
rect 13403 16028 13415 16031
rect 13538 16028 13544 16040
rect 13403 16000 13544 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 16908 16000 17233 16028
rect 16908 15988 16914 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 22112 16028 22140 16068
rect 21232 16000 22140 16028
rect 23768 16028 23796 16068
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 27154 16096 27160 16108
rect 23891 16068 27160 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27617 16099 27675 16105
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 27663 16068 29408 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 29380 16028 29408 16068
rect 29454 16056 29460 16108
rect 29512 16096 29518 16108
rect 29512 16068 29557 16096
rect 29512 16056 29518 16068
rect 29638 16056 29644 16108
rect 29696 16096 29702 16108
rect 32306 16096 32312 16108
rect 29696 16068 31754 16096
rect 32219 16068 32312 16096
rect 29696 16056 29702 16068
rect 29822 16028 29828 16040
rect 23768 16000 27614 16028
rect 29380 16000 29828 16028
rect 21232 15988 21238 16000
rect 27586 15972 27614 16000
rect 29822 15988 29828 16000
rect 29880 15988 29886 16040
rect 31726 16028 31754 16068
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 32565 16099 32623 16105
rect 32565 16096 32577 16099
rect 32456 16068 32577 16096
rect 32456 16056 32462 16068
rect 32565 16065 32577 16068
rect 32611 16065 32623 16099
rect 32565 16059 32623 16065
rect 33704 16040 33732 16136
rect 34422 16124 34428 16176
rect 34480 16164 34486 16176
rect 34480 16136 35112 16164
rect 34480 16124 34486 16136
rect 34514 16105 34520 16108
rect 34508 16096 34520 16105
rect 34475 16068 34520 16096
rect 34508 16059 34520 16068
rect 34514 16056 34520 16059
rect 34572 16056 34578 16108
rect 35084 16096 35112 16136
rect 35158 16124 35164 16176
rect 35216 16164 35222 16176
rect 40586 16164 40592 16176
rect 35216 16136 40592 16164
rect 35216 16124 35222 16136
rect 40586 16124 40592 16136
rect 40644 16124 40650 16176
rect 41506 16124 41512 16176
rect 41564 16164 41570 16176
rect 43088 16173 43116 16204
rect 44542 16192 44548 16204
rect 44600 16232 44606 16244
rect 48682 16232 48688 16244
rect 44600 16204 48360 16232
rect 48643 16204 48688 16232
rect 44600 16192 44606 16204
rect 43073 16167 43131 16173
rect 43073 16164 43085 16167
rect 41564 16136 43085 16164
rect 41564 16124 41570 16136
rect 43073 16133 43085 16136
rect 43119 16133 43131 16167
rect 43073 16127 43131 16133
rect 43165 16167 43223 16173
rect 43165 16133 43177 16167
rect 43211 16164 43223 16167
rect 44168 16167 44226 16173
rect 43211 16136 44128 16164
rect 43211 16133 43223 16136
rect 43165 16127 43223 16133
rect 37458 16096 37464 16108
rect 35084 16068 36676 16096
rect 37419 16068 37464 16096
rect 31726 16000 32352 16028
rect 12216 15932 12664 15960
rect 12216 15920 12222 15932
rect 13262 15920 13268 15972
rect 13320 15960 13326 15972
rect 18601 15963 18659 15969
rect 13320 15932 17264 15960
rect 13320 15920 13326 15932
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12084 15864 12909 15892
rect 12897 15861 12909 15864
rect 12943 15892 12955 15895
rect 14550 15892 14556 15904
rect 12943 15864 14556 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 14550 15852 14556 15864
rect 14608 15852 14614 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 17236 15892 17264 15932
rect 18601 15929 18613 15963
rect 18647 15960 18659 15963
rect 24210 15960 24216 15972
rect 18647 15932 20484 15960
rect 18647 15929 18659 15932
rect 18601 15923 18659 15929
rect 17862 15892 17868 15904
rect 17236 15864 17868 15892
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 18230 15852 18236 15904
rect 18288 15892 18294 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 18288 15864 20361 15892
rect 18288 15852 18294 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20456 15892 20484 15932
rect 23216 15932 24216 15960
rect 23216 15892 23244 15932
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 27586 15932 27620 15972
rect 27614 15920 27620 15932
rect 27672 15920 27678 15972
rect 20456 15864 23244 15892
rect 23385 15895 23443 15901
rect 20349 15855 20407 15861
rect 23385 15861 23397 15895
rect 23431 15892 23443 15895
rect 24026 15892 24032 15904
rect 23431 15864 24032 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 24486 15852 24492 15904
rect 24544 15892 24550 15904
rect 30098 15892 30104 15904
rect 24544 15864 30104 15892
rect 24544 15852 24550 15864
rect 30098 15852 30104 15864
rect 30156 15852 30162 15904
rect 30650 15892 30656 15904
rect 30611 15864 30656 15892
rect 30650 15852 30656 15864
rect 30708 15852 30714 15904
rect 32324 15892 32352 16000
rect 33686 15988 33692 16040
rect 33744 16028 33750 16040
rect 34238 16028 34244 16040
rect 33744 16000 34244 16028
rect 33744 15988 33750 16000
rect 34238 15988 34244 16000
rect 34296 15988 34302 16040
rect 35618 15988 35624 16040
rect 35676 16028 35682 16040
rect 36648 16037 36676 16068
rect 37458 16056 37464 16068
rect 37516 16056 37522 16108
rect 37550 16056 37556 16108
rect 37608 16096 37614 16108
rect 37717 16099 37775 16105
rect 37717 16096 37729 16099
rect 37608 16068 37729 16096
rect 37608 16056 37614 16068
rect 37717 16065 37729 16068
rect 37763 16065 37775 16099
rect 37717 16059 37775 16065
rect 38194 16056 38200 16108
rect 38252 16096 38258 16108
rect 39577 16099 39635 16105
rect 39577 16096 39589 16099
rect 38252 16094 39436 16096
rect 39500 16094 39589 16096
rect 38252 16068 39589 16094
rect 38252 16056 38258 16068
rect 39408 16066 39528 16068
rect 39577 16065 39589 16068
rect 39623 16065 39635 16099
rect 39577 16059 39635 16065
rect 39758 16056 39764 16108
rect 39816 16096 39822 16108
rect 40218 16096 40224 16108
rect 39816 16068 39861 16096
rect 40179 16068 40224 16096
rect 39816 16056 39822 16068
rect 40218 16056 40224 16068
rect 40276 16056 40282 16108
rect 40402 16096 40408 16108
rect 40363 16068 40408 16096
rect 40402 16056 40408 16068
rect 40460 16056 40466 16108
rect 40512 16068 42012 16096
rect 36541 16031 36599 16037
rect 36541 16028 36553 16031
rect 35676 16000 36553 16028
rect 35676 15988 35682 16000
rect 36541 15997 36553 16000
rect 36587 15997 36599 16031
rect 36541 15991 36599 15997
rect 36633 16031 36691 16037
rect 36633 15997 36645 16031
rect 36679 15997 36691 16031
rect 36633 15991 36691 15997
rect 38654 15988 38660 16040
rect 38712 16028 38718 16040
rect 39114 16028 39120 16040
rect 38712 16000 39120 16028
rect 38712 15988 38718 16000
rect 39114 15988 39120 16000
rect 39172 16028 39178 16040
rect 39393 16031 39451 16037
rect 39393 16028 39405 16031
rect 39172 16000 39405 16028
rect 39172 15988 39178 16000
rect 39393 15997 39405 16000
rect 39439 15997 39451 16031
rect 40512 16028 40540 16068
rect 41782 16028 41788 16040
rect 39393 15991 39451 15997
rect 39500 16000 40540 16028
rect 41743 16000 41788 16028
rect 36081 15963 36139 15969
rect 36081 15960 36093 15963
rect 35176 15932 36093 15960
rect 33410 15892 33416 15904
rect 32324 15864 33416 15892
rect 33410 15852 33416 15864
rect 33468 15852 33474 15904
rect 33962 15852 33968 15904
rect 34020 15892 34026 15904
rect 35176 15892 35204 15932
rect 36081 15929 36093 15932
rect 36127 15929 36139 15963
rect 36081 15923 36139 15929
rect 36170 15920 36176 15972
rect 36228 15960 36234 15972
rect 37182 15960 37188 15972
rect 36228 15932 37188 15960
rect 36228 15920 36234 15932
rect 37182 15920 37188 15932
rect 37240 15920 37246 15972
rect 39206 15920 39212 15972
rect 39264 15960 39270 15972
rect 39500 15960 39528 16000
rect 41782 15988 41788 16000
rect 41840 15988 41846 16040
rect 41877 16031 41935 16037
rect 41877 15997 41889 16031
rect 41923 15997 41935 16031
rect 41984 16028 42012 16068
rect 42150 16056 42156 16108
rect 42208 16096 42214 16108
rect 42889 16099 42947 16105
rect 42889 16096 42901 16099
rect 42208 16068 42901 16096
rect 42208 16056 42214 16068
rect 42889 16065 42901 16068
rect 42935 16065 42947 16099
rect 42889 16059 42947 16065
rect 43257 16099 43315 16105
rect 43257 16065 43269 16099
rect 43303 16096 43315 16099
rect 43990 16096 43996 16108
rect 43303 16068 43996 16096
rect 43303 16065 43315 16068
rect 43257 16059 43315 16065
rect 43272 16028 43300 16059
rect 43990 16056 43996 16068
rect 44048 16056 44054 16108
rect 44100 16096 44128 16136
rect 44168 16133 44180 16167
rect 44214 16164 44226 16167
rect 44266 16164 44272 16176
rect 44214 16136 44272 16164
rect 44214 16133 44226 16136
rect 44168 16127 44226 16133
rect 44266 16124 44272 16136
rect 44324 16124 44330 16176
rect 45462 16124 45468 16176
rect 45520 16164 45526 16176
rect 48332 16173 48360 16204
rect 48682 16192 48688 16204
rect 48740 16192 48746 16244
rect 49513 16235 49571 16241
rect 49513 16201 49525 16235
rect 49559 16232 49571 16235
rect 49970 16232 49976 16244
rect 49559 16204 49976 16232
rect 49559 16201 49571 16204
rect 49513 16195 49571 16201
rect 49970 16192 49976 16204
rect 50028 16192 50034 16244
rect 48317 16167 48375 16173
rect 45520 16136 48268 16164
rect 45520 16124 45526 16136
rect 44100 16068 45324 16096
rect 41984 16000 43300 16028
rect 43901 16031 43959 16037
rect 41877 15991 41935 15997
rect 43901 15997 43913 16031
rect 43947 15997 43959 16031
rect 43901 15991 43959 15997
rect 39264 15932 39528 15960
rect 39264 15920 39270 15932
rect 40034 15920 40040 15972
rect 40092 15960 40098 15972
rect 41892 15960 41920 15991
rect 43162 15960 43168 15972
rect 40092 15932 43168 15960
rect 40092 15920 40098 15932
rect 43162 15920 43168 15932
rect 43220 15920 43226 15972
rect 34020 15864 35204 15892
rect 34020 15852 34026 15864
rect 37734 15852 37740 15904
rect 37792 15892 37798 15904
rect 38841 15895 38899 15901
rect 38841 15892 38853 15895
rect 37792 15864 38853 15892
rect 37792 15852 37798 15864
rect 38841 15861 38853 15864
rect 38887 15861 38899 15895
rect 40586 15892 40592 15904
rect 40547 15864 40592 15892
rect 38841 15855 38899 15861
rect 40586 15852 40592 15864
rect 40644 15852 40650 15904
rect 41322 15892 41328 15904
rect 41283 15864 41328 15892
rect 41322 15852 41328 15864
rect 41380 15852 41386 15904
rect 43438 15892 43444 15904
rect 43399 15864 43444 15892
rect 43438 15852 43444 15864
rect 43496 15852 43502 15904
rect 43916 15892 43944 15991
rect 45296 15969 45324 16068
rect 45738 16056 45744 16108
rect 45796 16096 45802 16108
rect 46385 16099 46443 16105
rect 46385 16096 46397 16099
rect 45796 16068 46397 16096
rect 45796 16056 45802 16068
rect 46385 16065 46397 16068
rect 46431 16065 46443 16099
rect 46385 16059 46443 16065
rect 46474 16056 46480 16108
rect 46532 16096 46538 16108
rect 48133 16099 48191 16105
rect 48133 16096 48145 16099
rect 46532 16068 48145 16096
rect 46532 16056 46538 16068
rect 48133 16065 48145 16068
rect 48179 16065 48191 16099
rect 48240 16096 48268 16136
rect 48317 16133 48329 16167
rect 48363 16133 48375 16167
rect 48317 16127 48375 16133
rect 48409 16167 48467 16173
rect 48409 16133 48421 16167
rect 48455 16164 48467 16167
rect 49694 16164 49700 16176
rect 48455 16136 49700 16164
rect 48455 16133 48467 16136
rect 48409 16127 48467 16133
rect 49694 16124 49700 16136
rect 49752 16124 49758 16176
rect 48501 16099 48559 16105
rect 48501 16096 48513 16099
rect 48240 16068 48513 16096
rect 48133 16059 48191 16065
rect 48501 16065 48513 16068
rect 48547 16065 48559 16099
rect 48501 16059 48559 16065
rect 46198 16028 46204 16040
rect 46111 16000 46204 16028
rect 46198 15988 46204 16000
rect 46256 16028 46262 16040
rect 46842 16028 46848 16040
rect 46256 16000 46848 16028
rect 46256 15988 46262 16000
rect 46842 15988 46848 16000
rect 46900 15988 46906 16040
rect 48516 16028 48544 16059
rect 48866 16056 48872 16108
rect 48924 16096 48930 16108
rect 49145 16099 49203 16105
rect 49145 16096 49157 16099
rect 48924 16068 49157 16096
rect 48924 16056 48930 16068
rect 49145 16065 49157 16068
rect 49191 16065 49203 16099
rect 49145 16059 49203 16065
rect 49234 16056 49240 16108
rect 49292 16096 49298 16108
rect 49329 16099 49387 16105
rect 49329 16096 49341 16099
rect 49292 16068 49341 16096
rect 49292 16056 49298 16068
rect 49329 16065 49341 16068
rect 49375 16065 49387 16099
rect 49329 16059 49387 16065
rect 49418 16028 49424 16040
rect 48516 16000 49424 16028
rect 49418 15988 49424 16000
rect 49476 15988 49482 16040
rect 45281 15963 45339 15969
rect 45281 15929 45293 15963
rect 45327 15960 45339 15963
rect 57790 15960 57796 15972
rect 45327 15932 57796 15960
rect 45327 15929 45339 15932
rect 45281 15923 45339 15929
rect 57790 15920 57796 15932
rect 57848 15920 57854 15972
rect 44174 15892 44180 15904
rect 43916 15864 44180 15892
rect 44174 15852 44180 15864
rect 44232 15852 44238 15904
rect 46566 15892 46572 15904
rect 46527 15864 46572 15892
rect 46566 15852 46572 15864
rect 46624 15852 46630 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 17770 15688 17776 15700
rect 17731 15660 17776 15688
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 17862 15648 17868 15700
rect 17920 15688 17926 15700
rect 17920 15660 26832 15688
rect 17920 15648 17926 15660
rect 17310 15580 17316 15632
rect 17368 15620 17374 15632
rect 18230 15620 18236 15632
rect 17368 15592 18236 15620
rect 17368 15580 17374 15592
rect 18230 15580 18236 15592
rect 18288 15580 18294 15632
rect 20530 15580 20536 15632
rect 20588 15620 20594 15632
rect 22557 15623 22615 15629
rect 22557 15620 22569 15623
rect 20588 15592 22569 15620
rect 20588 15580 20594 15592
rect 22557 15589 22569 15592
rect 22603 15589 22615 15623
rect 22557 15583 22615 15589
rect 23474 15580 23480 15632
rect 23532 15620 23538 15632
rect 24762 15620 24768 15632
rect 23532 15592 24768 15620
rect 23532 15580 23538 15592
rect 24762 15580 24768 15592
rect 24820 15580 24826 15632
rect 25222 15580 25228 15632
rect 25280 15620 25286 15632
rect 26510 15620 26516 15632
rect 25280 15592 26516 15620
rect 25280 15580 25286 15592
rect 26510 15580 26516 15592
rect 26568 15580 26574 15632
rect 26804 15620 26832 15660
rect 27154 15648 27160 15700
rect 27212 15688 27218 15700
rect 41782 15688 41788 15700
rect 27212 15660 41788 15688
rect 27212 15648 27218 15660
rect 41782 15648 41788 15660
rect 41840 15648 41846 15700
rect 42886 15688 42892 15700
rect 42847 15660 42892 15688
rect 42886 15648 42892 15660
rect 42944 15648 42950 15700
rect 45738 15688 45744 15700
rect 45699 15660 45744 15688
rect 45738 15648 45744 15660
rect 45796 15648 45802 15700
rect 48130 15688 48136 15700
rect 48091 15660 48136 15688
rect 48130 15648 48136 15660
rect 48188 15648 48194 15700
rect 30285 15623 30343 15629
rect 26804 15592 29132 15620
rect 2406 15512 2412 15564
rect 2464 15552 2470 15564
rect 13725 15555 13783 15561
rect 2464 15524 2774 15552
rect 2464 15512 2470 15524
rect 2746 15348 2774 15524
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 13771 15524 14749 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 16390 15512 16396 15564
rect 16448 15552 16454 15564
rect 17770 15552 17776 15564
rect 16448 15524 17776 15552
rect 16448 15512 16454 15524
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 25130 15552 25136 15564
rect 20916 15524 25136 15552
rect 11422 15484 11428 15496
rect 11383 15456 11428 15484
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13964 15456 14473 15484
rect 13964 15444 13970 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 16574 15484 16580 15496
rect 14608 15456 16436 15484
rect 16535 15456 16580 15484
rect 14608 15444 14614 15456
rect 16117 15419 16175 15425
rect 16117 15385 16129 15419
rect 16163 15416 16175 15419
rect 16298 15416 16304 15428
rect 16163 15388 16304 15416
rect 16163 15385 16175 15388
rect 16117 15379 16175 15385
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 16408 15416 16436 15456
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19484 15456 19533 15484
rect 19484 15444 19490 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19788 15487 19846 15493
rect 19788 15453 19800 15487
rect 19834 15484 19846 15487
rect 20916 15484 20944 15524
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 25777 15555 25835 15561
rect 25777 15521 25789 15555
rect 25823 15552 25835 15555
rect 26050 15552 26056 15564
rect 25823 15524 26056 15552
rect 25823 15521 25835 15524
rect 25777 15515 25835 15521
rect 26050 15512 26056 15524
rect 26108 15512 26114 15564
rect 28074 15552 28080 15564
rect 28035 15524 28080 15552
rect 28074 15512 28080 15524
rect 28132 15512 28138 15564
rect 21358 15484 21364 15496
rect 19834 15456 20944 15484
rect 21319 15456 21364 15484
rect 19834 15453 19846 15456
rect 19788 15447 19846 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 22020 15456 22140 15484
rect 22020 15416 22048 15456
rect 16408 15388 22048 15416
rect 22112 15416 22140 15456
rect 25038 15444 25044 15496
rect 25096 15484 25102 15496
rect 26329 15487 26387 15493
rect 26329 15484 26341 15487
rect 25096 15456 26341 15484
rect 25096 15444 25102 15456
rect 26329 15453 26341 15456
rect 26375 15484 26387 15487
rect 28994 15484 29000 15496
rect 26375 15456 29000 15484
rect 26375 15453 26387 15456
rect 26329 15447 26387 15453
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 27154 15416 27160 15428
rect 22112 15388 27160 15416
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 28442 15416 28448 15428
rect 27448 15388 28448 15416
rect 19978 15348 19984 15360
rect 2746 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20898 15348 20904 15360
rect 20859 15320 20904 15348
rect 20898 15308 20904 15320
rect 20956 15348 20962 15360
rect 25038 15348 25044 15360
rect 20956 15320 25044 15348
rect 20956 15308 20962 15320
rect 25038 15308 25044 15320
rect 25096 15308 25102 15360
rect 25133 15351 25191 15357
rect 25133 15317 25145 15351
rect 25179 15348 25191 15351
rect 25222 15348 25228 15360
rect 25179 15320 25228 15348
rect 25179 15317 25191 15320
rect 25133 15311 25191 15317
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 25498 15348 25504 15360
rect 25459 15320 25504 15348
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 25866 15348 25872 15360
rect 25639 15320 25872 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 25866 15308 25872 15320
rect 25924 15348 25930 15360
rect 27448 15348 27476 15388
rect 28442 15376 28448 15388
rect 28500 15376 28506 15428
rect 29104 15416 29132 15592
rect 30285 15589 30297 15623
rect 30331 15620 30343 15623
rect 31294 15620 31300 15632
rect 30331 15592 31300 15620
rect 30331 15589 30343 15592
rect 30285 15583 30343 15589
rect 31294 15580 31300 15592
rect 31352 15580 31358 15632
rect 31478 15580 31484 15632
rect 31536 15580 31542 15632
rect 32861 15623 32919 15629
rect 32861 15589 32873 15623
rect 32907 15620 32919 15623
rect 33410 15620 33416 15632
rect 32907 15592 33416 15620
rect 32907 15589 32919 15592
rect 32861 15583 32919 15589
rect 33410 15580 33416 15592
rect 33468 15580 33474 15632
rect 34054 15580 34060 15632
rect 34112 15620 34118 15632
rect 37461 15623 37519 15629
rect 34112 15592 35379 15620
rect 34112 15580 34118 15592
rect 29914 15512 29920 15564
rect 29972 15552 29978 15564
rect 30837 15555 30895 15561
rect 30837 15552 30849 15555
rect 29972 15524 30849 15552
rect 29972 15512 29978 15524
rect 30837 15521 30849 15524
rect 30883 15552 30895 15555
rect 31496 15552 31524 15580
rect 34149 15555 34207 15561
rect 34149 15552 34161 15555
rect 30883 15524 31524 15552
rect 32488 15524 34161 15552
rect 30883 15521 30895 15524
rect 30837 15515 30895 15521
rect 30653 15487 30711 15493
rect 30653 15453 30665 15487
rect 30699 15484 30711 15487
rect 30926 15484 30932 15496
rect 30699 15456 30932 15484
rect 30699 15453 30711 15456
rect 30653 15447 30711 15453
rect 30926 15444 30932 15456
rect 30984 15444 30990 15496
rect 31481 15487 31539 15493
rect 31481 15453 31493 15487
rect 31527 15484 31539 15487
rect 32306 15484 32312 15496
rect 31527 15456 32312 15484
rect 31527 15453 31539 15456
rect 31481 15447 31539 15453
rect 32306 15444 32312 15456
rect 32364 15444 32370 15496
rect 31570 15416 31576 15428
rect 29104 15388 31576 15416
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 31748 15419 31806 15425
rect 31748 15385 31760 15419
rect 31794 15416 31806 15419
rect 31846 15416 31852 15428
rect 31794 15388 31852 15416
rect 31794 15385 31806 15388
rect 31748 15379 31806 15385
rect 31846 15376 31852 15388
rect 31904 15376 31910 15428
rect 25924 15320 27476 15348
rect 25924 15308 25930 15320
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 29454 15348 29460 15360
rect 27580 15320 29460 15348
rect 27580 15308 27586 15320
rect 29454 15308 29460 15320
rect 29512 15348 29518 15360
rect 30558 15348 30564 15360
rect 29512 15320 30564 15348
rect 29512 15308 29518 15320
rect 30558 15308 30564 15320
rect 30616 15308 30622 15360
rect 30742 15348 30748 15360
rect 30703 15320 30748 15348
rect 30742 15308 30748 15320
rect 30800 15308 30806 15360
rect 31478 15308 31484 15360
rect 31536 15348 31542 15360
rect 32488 15348 32516 15524
rect 34149 15521 34161 15524
rect 34195 15552 34207 15555
rect 34422 15552 34428 15564
rect 34195 15524 34428 15552
rect 34195 15521 34207 15524
rect 34149 15515 34207 15521
rect 34422 15512 34428 15524
rect 34480 15512 34486 15564
rect 34054 15484 34060 15496
rect 34015 15456 34060 15484
rect 34054 15444 34060 15456
rect 34112 15444 34118 15496
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34756 15456 34897 15484
rect 34756 15444 34762 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 35066 15484 35072 15496
rect 35027 15456 35072 15484
rect 34885 15447 34943 15453
rect 35066 15444 35072 15456
rect 35124 15444 35130 15496
rect 35351 15484 35379 15592
rect 37461 15589 37473 15623
rect 37507 15620 37519 15623
rect 37550 15620 37556 15632
rect 37507 15592 37556 15620
rect 37507 15589 37519 15592
rect 37461 15583 37519 15589
rect 37550 15580 37556 15592
rect 37608 15580 37614 15632
rect 38657 15623 38715 15629
rect 38657 15589 38669 15623
rect 38703 15620 38715 15623
rect 39942 15620 39948 15632
rect 38703 15592 39948 15620
rect 38703 15589 38715 15592
rect 38657 15583 38715 15589
rect 39942 15580 39948 15592
rect 40000 15580 40006 15632
rect 35434 15512 35440 15564
rect 35492 15552 35498 15564
rect 35529 15555 35587 15561
rect 35529 15552 35541 15555
rect 35492 15524 35541 15552
rect 35492 15512 35498 15524
rect 35529 15521 35541 15524
rect 35575 15521 35587 15555
rect 35529 15515 35587 15521
rect 36906 15512 36912 15564
rect 36964 15552 36970 15564
rect 38102 15552 38108 15564
rect 36964 15524 37274 15552
rect 38063 15524 38108 15552
rect 36964 15512 36970 15524
rect 35351 15456 36952 15484
rect 35774 15419 35832 15425
rect 35774 15416 35786 15419
rect 33612 15388 35786 15416
rect 33612 15357 33640 15388
rect 35774 15385 35786 15388
rect 35820 15385 35832 15419
rect 35774 15379 35832 15385
rect 31536 15320 32516 15348
rect 33597 15351 33655 15357
rect 31536 15308 31542 15320
rect 33597 15317 33609 15351
rect 33643 15317 33655 15351
rect 33597 15311 33655 15317
rect 33965 15351 34023 15357
rect 33965 15317 33977 15351
rect 34011 15348 34023 15351
rect 34882 15348 34888 15360
rect 34011 15320 34888 15348
rect 34011 15317 34023 15320
rect 33965 15311 34023 15317
rect 34882 15308 34888 15320
rect 34940 15308 34946 15360
rect 34977 15351 35035 15357
rect 34977 15317 34989 15351
rect 35023 15348 35035 15351
rect 35342 15348 35348 15360
rect 35023 15320 35348 15348
rect 35023 15317 35035 15320
rect 34977 15311 35035 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 36078 15308 36084 15360
rect 36136 15348 36142 15360
rect 36630 15348 36636 15360
rect 36136 15320 36636 15348
rect 36136 15308 36142 15320
rect 36630 15308 36636 15320
rect 36688 15308 36694 15360
rect 36924 15357 36952 15456
rect 37246 15416 37274 15524
rect 38102 15512 38108 15524
rect 38160 15512 38166 15564
rect 38672 15524 38976 15552
rect 37734 15444 37740 15496
rect 37792 15484 37798 15496
rect 37921 15487 37979 15493
rect 37921 15484 37933 15487
rect 37792 15456 37933 15484
rect 37792 15444 37798 15456
rect 37921 15453 37933 15456
rect 37967 15453 37979 15487
rect 37921 15447 37979 15453
rect 38672 15416 38700 15524
rect 38948 15493 38976 15524
rect 41046 15512 41052 15564
rect 41104 15552 41110 15564
rect 41104 15524 46888 15552
rect 41104 15512 41110 15524
rect 39206 15493 39212 15496
rect 38934 15487 38992 15493
rect 38842 15465 38900 15471
rect 38842 15431 38854 15465
rect 38888 15431 38900 15465
rect 38934 15453 38946 15487
rect 38980 15453 38992 15487
rect 38934 15447 38992 15453
rect 39163 15487 39212 15493
rect 39163 15453 39175 15487
rect 39209 15453 39212 15487
rect 39163 15447 39212 15453
rect 39206 15444 39212 15447
rect 39264 15444 39270 15496
rect 39301 15487 39359 15493
rect 39301 15453 39313 15487
rect 39347 15484 39359 15487
rect 39850 15484 39856 15496
rect 39347 15456 39856 15484
rect 39347 15453 39359 15456
rect 39301 15447 39359 15453
rect 39850 15444 39856 15456
rect 39908 15444 39914 15496
rect 41506 15484 41512 15496
rect 39960 15456 41512 15484
rect 38842 15428 38900 15431
rect 37246 15388 38700 15416
rect 38838 15376 38844 15428
rect 38896 15376 38902 15428
rect 39050 15419 39108 15425
rect 39050 15385 39062 15419
rect 39096 15416 39108 15419
rect 39960 15416 39988 15456
rect 41506 15444 41512 15456
rect 41564 15444 41570 15496
rect 41616 15493 41644 15524
rect 41601 15487 41659 15493
rect 41601 15453 41613 15487
rect 41647 15453 41659 15487
rect 41601 15447 41659 15453
rect 44082 15444 44088 15496
rect 44140 15484 44146 15496
rect 44177 15487 44235 15493
rect 44177 15484 44189 15487
rect 44140 15456 44189 15484
rect 44140 15444 44146 15456
rect 44177 15453 44189 15456
rect 44223 15484 44235 15487
rect 44542 15484 44548 15496
rect 44223 15456 44548 15484
rect 44223 15453 44235 15456
rect 44177 15447 44235 15453
rect 44542 15444 44548 15456
rect 44600 15444 44606 15496
rect 45186 15484 45192 15496
rect 45147 15456 45192 15484
rect 45186 15444 45192 15456
rect 45244 15444 45250 15496
rect 45557 15487 45615 15493
rect 45557 15453 45569 15487
rect 45603 15484 45615 15487
rect 46658 15484 46664 15496
rect 45603 15456 46664 15484
rect 45603 15453 45615 15456
rect 45557 15447 45615 15453
rect 46658 15444 46664 15456
rect 46716 15444 46722 15496
rect 39096 15388 39988 15416
rect 40037 15419 40095 15425
rect 39096 15385 39108 15388
rect 39050 15379 39108 15385
rect 40037 15385 40049 15419
rect 40083 15385 40095 15419
rect 40037 15379 40095 15385
rect 36909 15351 36967 15357
rect 36909 15317 36921 15351
rect 36955 15317 36967 15351
rect 36909 15311 36967 15317
rect 37829 15351 37887 15357
rect 37829 15317 37841 15351
rect 37875 15348 37887 15351
rect 38746 15348 38752 15360
rect 37875 15320 38752 15348
rect 37875 15317 37887 15320
rect 37829 15311 37887 15317
rect 38746 15308 38752 15320
rect 38804 15308 38810 15360
rect 40052 15348 40080 15379
rect 40126 15376 40132 15428
rect 40184 15416 40190 15428
rect 40221 15419 40279 15425
rect 40221 15416 40233 15419
rect 40184 15388 40233 15416
rect 40184 15376 40190 15388
rect 40221 15385 40233 15388
rect 40267 15385 40279 15419
rect 40221 15379 40279 15385
rect 44358 15376 44364 15428
rect 44416 15416 44422 15428
rect 44453 15419 44511 15425
rect 44453 15416 44465 15419
rect 44416 15388 44465 15416
rect 44416 15376 44422 15388
rect 44453 15385 44465 15388
rect 44499 15416 44511 15419
rect 45373 15419 45431 15425
rect 45373 15416 45385 15419
rect 44499 15388 45385 15416
rect 44499 15385 44511 15388
rect 44453 15379 44511 15385
rect 45373 15385 45385 15388
rect 45419 15385 45431 15419
rect 45373 15379 45431 15385
rect 45465 15419 45523 15425
rect 45465 15385 45477 15419
rect 45511 15416 45523 15419
rect 46750 15416 46756 15428
rect 45511 15388 46756 15416
rect 45511 15385 45523 15388
rect 45465 15379 45523 15385
rect 46750 15376 46756 15388
rect 46808 15376 46814 15428
rect 46860 15425 46888 15524
rect 48866 15512 48872 15564
rect 48924 15552 48930 15564
rect 50341 15555 50399 15561
rect 50341 15552 50353 15555
rect 48924 15524 50353 15552
rect 48924 15512 48930 15524
rect 50341 15521 50353 15524
rect 50387 15521 50399 15555
rect 50341 15515 50399 15521
rect 47118 15444 47124 15496
rect 47176 15484 47182 15496
rect 49053 15487 49111 15493
rect 49053 15484 49065 15487
rect 47176 15456 49065 15484
rect 47176 15444 47182 15456
rect 49053 15453 49065 15456
rect 49099 15453 49111 15487
rect 49418 15484 49424 15496
rect 49379 15456 49424 15484
rect 49053 15447 49111 15453
rect 49418 15444 49424 15456
rect 49476 15444 49482 15496
rect 49786 15484 49792 15496
rect 49528 15456 49792 15484
rect 46845 15419 46903 15425
rect 46845 15385 46857 15419
rect 46891 15416 46903 15419
rect 47210 15416 47216 15428
rect 46891 15388 47216 15416
rect 46891 15385 46903 15388
rect 46845 15379 46903 15385
rect 47210 15376 47216 15388
rect 47268 15376 47274 15428
rect 48038 15376 48044 15428
rect 48096 15416 48102 15428
rect 49237 15419 49295 15425
rect 49237 15416 49249 15419
rect 48096 15388 49249 15416
rect 48096 15376 48102 15388
rect 49237 15385 49249 15388
rect 49283 15385 49295 15419
rect 49237 15379 49295 15385
rect 49329 15419 49387 15425
rect 49329 15385 49341 15419
rect 49375 15416 49387 15419
rect 49528 15416 49556 15456
rect 49786 15444 49792 15456
rect 49844 15444 49850 15496
rect 50525 15487 50583 15493
rect 50525 15453 50537 15487
rect 50571 15453 50583 15487
rect 50525 15447 50583 15453
rect 50540 15416 50568 15447
rect 56502 15444 56508 15496
rect 56560 15484 56566 15496
rect 57885 15487 57943 15493
rect 57885 15484 57897 15487
rect 56560 15456 57897 15484
rect 56560 15444 56566 15456
rect 57885 15453 57897 15456
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 58158 15416 58164 15428
rect 49375 15388 49556 15416
rect 49620 15388 50568 15416
rect 58119 15388 58164 15416
rect 49375 15385 49387 15388
rect 49329 15379 49387 15385
rect 40310 15348 40316 15360
rect 40052 15320 40316 15348
rect 40310 15308 40316 15320
rect 40368 15308 40374 15360
rect 40405 15351 40463 15357
rect 40405 15317 40417 15351
rect 40451 15348 40463 15351
rect 40586 15348 40592 15360
rect 40451 15320 40592 15348
rect 40451 15317 40463 15320
rect 40405 15311 40463 15317
rect 40586 15308 40592 15320
rect 40644 15308 40650 15360
rect 43254 15308 43260 15360
rect 43312 15348 43318 15360
rect 46198 15348 46204 15360
rect 43312 15320 46204 15348
rect 43312 15308 43318 15320
rect 46198 15308 46204 15320
rect 46256 15308 46262 15360
rect 49620 15357 49648 15388
rect 58158 15376 58164 15388
rect 58216 15376 58222 15428
rect 49605 15351 49663 15357
rect 49605 15317 49617 15351
rect 49651 15317 49663 15351
rect 50706 15348 50712 15360
rect 50667 15320 50712 15348
rect 49605 15311 49663 15317
rect 50706 15308 50712 15320
rect 50764 15308 50770 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 10980 15116 15148 15144
rect 10980 15017 11008 15116
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 10965 15011 11023 15017
rect 1627 14980 2452 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 2424 14952 2452 14980
rect 10965 14977 10977 15011
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11238 15008 11244 15020
rect 11195 14980 11244 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 13906 15008 13912 15020
rect 11900 14980 13912 15008
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2406 14940 2412 14952
rect 2367 14912 2412 14940
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 11900 14949 11928 14980
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 15120 15008 15148 15116
rect 16022 15104 16028 15156
rect 16080 15144 16086 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 16080 15116 16221 15144
rect 16080 15104 16086 15116
rect 16209 15113 16221 15116
rect 16255 15113 16267 15147
rect 16209 15107 16267 15113
rect 17034 15104 17040 15156
rect 17092 15144 17098 15156
rect 25130 15144 25136 15156
rect 17092 15116 23980 15144
rect 25091 15116 25136 15144
rect 17092 15104 17098 15116
rect 18322 15036 18328 15088
rect 18380 15076 18386 15088
rect 20898 15076 20904 15088
rect 18380 15048 20904 15076
rect 18380 15036 18386 15048
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 22462 15076 22468 15088
rect 22296 15048 22468 15076
rect 17954 15008 17960 15020
rect 14056 14980 14101 15008
rect 15120 14980 17960 15008
rect 14056 14968 14062 14980
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 8260 14912 11897 14940
rect 8260 14900 8266 14912
rect 11885 14909 11897 14912
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 13924 14940 13952 14968
rect 16850 14940 16856 14952
rect 12207 14912 13860 14940
rect 13924 14912 16856 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 10410 14832 10416 14884
rect 10468 14872 10474 14884
rect 13832 14872 13860 14912
rect 16850 14900 16856 14912
rect 16908 14940 16914 14952
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 16908 14912 17049 14940
rect 16908 14900 16914 14912
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 17276 14912 17325 14940
rect 17276 14900 17282 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 15378 14872 15384 14884
rect 10468 14844 11928 14872
rect 13832 14844 15384 14872
rect 10468 14832 10474 14844
rect 10962 14804 10968 14816
rect 10923 14776 10968 14804
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11900 14804 11928 14844
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 19168 14872 19196 14971
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22296 15008 22324 15048
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 23952 15017 23980 15116
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 28350 15104 28356 15156
rect 28408 15144 28414 15156
rect 29273 15147 29331 15153
rect 29273 15144 29285 15147
rect 28408 15116 29285 15144
rect 28408 15104 28414 15116
rect 29273 15113 29285 15116
rect 29319 15113 29331 15147
rect 30834 15144 30840 15156
rect 30795 15116 30840 15144
rect 29273 15107 29331 15113
rect 30834 15104 30840 15116
rect 30892 15104 30898 15156
rect 30926 15104 30932 15156
rect 30984 15144 30990 15156
rect 31297 15147 31355 15153
rect 31297 15144 31309 15147
rect 30984 15116 31309 15144
rect 30984 15104 30990 15116
rect 31297 15113 31309 15116
rect 31343 15113 31355 15147
rect 31297 15107 31355 15113
rect 32309 15147 32367 15153
rect 32309 15113 32321 15147
rect 32355 15144 32367 15147
rect 36170 15144 36176 15156
rect 32355 15116 36176 15144
rect 32355 15113 32367 15116
rect 32309 15107 32367 15113
rect 36170 15104 36176 15116
rect 36228 15104 36234 15156
rect 36630 15104 36636 15156
rect 36688 15144 36694 15156
rect 38838 15144 38844 15156
rect 36688 15116 38844 15144
rect 36688 15104 36694 15116
rect 38838 15104 38844 15116
rect 38896 15104 38902 15156
rect 39114 15104 39120 15156
rect 39172 15104 39178 15156
rect 41782 15104 41788 15156
rect 41840 15144 41846 15156
rect 41969 15147 42027 15153
rect 41969 15144 41981 15147
rect 41840 15116 41981 15144
rect 41840 15104 41846 15116
rect 41969 15113 41981 15116
rect 42015 15113 42027 15147
rect 41969 15107 42027 15113
rect 43073 15147 43131 15153
rect 43073 15113 43085 15147
rect 43119 15144 43131 15147
rect 44266 15144 44272 15156
rect 43119 15116 44272 15144
rect 43119 15113 43131 15116
rect 43073 15107 43131 15113
rect 44266 15104 44272 15116
rect 44324 15104 44330 15156
rect 44450 15104 44456 15156
rect 44508 15144 44514 15156
rect 45833 15147 45891 15153
rect 45833 15144 45845 15147
rect 44508 15116 45845 15144
rect 44508 15104 44514 15116
rect 45833 15113 45845 15116
rect 45879 15144 45891 15147
rect 45879 15116 51074 15144
rect 45879 15113 45891 15116
rect 45833 15107 45891 15113
rect 28994 15036 29000 15088
rect 29052 15076 29058 15088
rect 31018 15076 31024 15088
rect 29052 15048 31024 15076
rect 29052 15036 29058 15048
rect 31018 15036 31024 15048
rect 31076 15076 31082 15088
rect 32677 15079 32735 15085
rect 32677 15076 32689 15079
rect 31076 15048 32689 15076
rect 31076 15036 31082 15048
rect 32677 15045 32689 15048
rect 32723 15045 32735 15079
rect 32677 15039 32735 15045
rect 32766 15036 32772 15088
rect 32824 15076 32830 15088
rect 33962 15085 33968 15088
rect 33956 15076 33968 15085
rect 32824 15048 32869 15076
rect 33923 15048 33968 15076
rect 32824 15036 32830 15048
rect 33956 15039 33968 15048
rect 33962 15036 33968 15039
rect 34020 15036 34026 15088
rect 34330 15036 34336 15088
rect 34388 15076 34394 15088
rect 36078 15076 36084 15088
rect 34388 15048 36084 15076
rect 34388 15036 34394 15048
rect 22152 14980 22324 15008
rect 22364 15011 22422 15017
rect 22152 14968 22158 14980
rect 22364 14977 22376 15011
rect 22410 15008 22422 15011
rect 23937 15011 23995 15017
rect 22410 14980 23888 15008
rect 22410 14977 22422 14980
rect 22364 14971 22422 14977
rect 23860 14940 23888 14980
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 27246 15008 27252 15020
rect 27207 14980 27252 15008
rect 23937 14971 23995 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 30650 15008 30656 15020
rect 28123 14980 30656 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 30650 14968 30656 14980
rect 30708 14968 30714 15020
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 25590 14940 25596 14952
rect 23860 14912 25596 14940
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 30558 14900 30564 14952
rect 30616 14940 30622 14952
rect 31110 14940 31116 14952
rect 30616 14912 31116 14940
rect 30616 14900 30622 14912
rect 31110 14900 31116 14912
rect 31168 14940 31174 14952
rect 31220 14940 31248 14971
rect 32030 14968 32036 15020
rect 32088 15008 32094 15020
rect 35912 15017 35940 15048
rect 36078 15036 36084 15048
rect 36136 15036 36142 15088
rect 37458 15036 37464 15088
rect 37516 15076 37522 15088
rect 38010 15076 38016 15088
rect 37516 15048 38016 15076
rect 37516 15036 37522 15048
rect 38010 15036 38016 15048
rect 38068 15076 38074 15088
rect 39132 15076 39160 15104
rect 38068 15048 39160 15076
rect 38068 15036 38074 15048
rect 39390 15036 39396 15088
rect 39448 15036 39454 15088
rect 39574 15036 39580 15088
rect 39632 15076 39638 15088
rect 39850 15076 39856 15088
rect 39632 15048 39856 15076
rect 39632 15036 39638 15048
rect 39850 15036 39856 15048
rect 39908 15036 39914 15088
rect 40856 15079 40914 15085
rect 40856 15045 40868 15079
rect 40902 15076 40914 15079
rect 41322 15076 41328 15088
rect 40902 15048 41328 15076
rect 40902 15045 40914 15048
rect 40856 15039 40914 15045
rect 41322 15036 41328 15048
rect 41380 15036 41386 15088
rect 46569 15079 46627 15085
rect 42260 15048 46428 15076
rect 35713 15011 35771 15017
rect 35713 15008 35725 15011
rect 32088 14980 35725 15008
rect 32088 14968 32094 14980
rect 35713 14977 35725 14980
rect 35759 14977 35771 15011
rect 35713 14971 35771 14977
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 14977 35955 15011
rect 35897 14971 35955 14977
rect 35989 15011 36047 15017
rect 35989 14977 36001 15011
rect 36035 14977 36047 15011
rect 36725 15011 36783 15017
rect 36725 15008 36737 15011
rect 35989 14971 36047 14977
rect 36372 14980 36737 15008
rect 31168 14912 31248 14940
rect 31389 14943 31447 14949
rect 31168 14900 31174 14912
rect 31389 14909 31401 14943
rect 31435 14909 31447 14943
rect 31389 14903 31447 14909
rect 32861 14943 32919 14949
rect 32861 14909 32873 14943
rect 32907 14909 32919 14943
rect 32861 14903 32919 14909
rect 17972 14844 19196 14872
rect 23477 14875 23535 14881
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 11900 14776 13277 14804
rect 13265 14773 13277 14776
rect 13311 14804 13323 14807
rect 13446 14804 13452 14816
rect 13311 14776 13452 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 17972 14804 18000 14844
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 25498 14872 25504 14884
rect 23523 14844 25504 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 15620 14776 18000 14804
rect 18601 14807 18659 14813
rect 15620 14764 15626 14776
rect 18601 14773 18613 14807
rect 18647 14804 18659 14807
rect 20898 14804 20904 14816
rect 18647 14776 20904 14804
rect 18647 14773 18659 14776
rect 18601 14767 18659 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21361 14807 21419 14813
rect 21361 14773 21373 14807
rect 21407 14804 21419 14807
rect 22278 14804 22284 14816
rect 21407 14776 22284 14804
rect 21407 14773 21419 14776
rect 21361 14767 21419 14773
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 22830 14764 22836 14816
rect 22888 14804 22894 14816
rect 23382 14804 23388 14816
rect 22888 14776 23388 14804
rect 22888 14764 22894 14776
rect 23382 14764 23388 14776
rect 23440 14804 23446 14816
rect 23492 14804 23520 14835
rect 25498 14832 25504 14844
rect 25556 14832 25562 14884
rect 31202 14872 31208 14884
rect 25608 14844 31208 14872
rect 23440 14776 23520 14804
rect 23440 14764 23446 14776
rect 23566 14764 23572 14816
rect 23624 14804 23630 14816
rect 25608 14804 25636 14844
rect 31202 14832 31208 14844
rect 31260 14832 31266 14884
rect 31404 14872 31432 14903
rect 31478 14872 31484 14884
rect 31391 14844 31484 14872
rect 23624 14776 25636 14804
rect 23624 14764 23630 14776
rect 27338 14764 27344 14816
rect 27396 14804 27402 14816
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 27396 14776 27537 14804
rect 27396 14764 27402 14776
rect 27525 14773 27537 14776
rect 27571 14804 27583 14807
rect 27798 14804 27804 14816
rect 27571 14776 27804 14804
rect 27571 14773 27583 14776
rect 27525 14767 27583 14773
rect 27798 14764 27804 14776
rect 27856 14764 27862 14816
rect 28074 14764 28080 14816
rect 28132 14804 28138 14816
rect 28902 14804 28908 14816
rect 28132 14776 28908 14804
rect 28132 14764 28138 14776
rect 28902 14764 28908 14776
rect 28960 14804 28966 14816
rect 31404 14804 31432 14844
rect 31478 14832 31484 14844
rect 31536 14872 31542 14884
rect 32876 14872 32904 14903
rect 32950 14900 32956 14952
rect 33008 14940 33014 14952
rect 33686 14940 33692 14952
rect 33008 14912 33692 14940
rect 33008 14900 33014 14912
rect 33686 14900 33692 14912
rect 33744 14900 33750 14952
rect 35526 14900 35532 14952
rect 35584 14940 35590 14952
rect 35805 14943 35863 14949
rect 35805 14940 35817 14943
rect 35584 14912 35817 14940
rect 35584 14900 35590 14912
rect 35805 14909 35817 14912
rect 35851 14909 35863 14943
rect 35805 14903 35863 14909
rect 35618 14872 35624 14884
rect 31536 14844 32904 14872
rect 35084 14844 35624 14872
rect 31536 14832 31542 14844
rect 28960 14776 31432 14804
rect 28960 14764 28966 14776
rect 31570 14764 31576 14816
rect 31628 14804 31634 14816
rect 35084 14813 35112 14844
rect 35618 14832 35624 14844
rect 35676 14832 35682 14884
rect 36004 14872 36032 14971
rect 36170 14900 36176 14952
rect 36228 14940 36234 14952
rect 36372 14940 36400 14980
rect 36725 14977 36737 14980
rect 36771 14977 36783 15011
rect 36725 14971 36783 14977
rect 36814 14968 36820 15020
rect 36872 15008 36878 15020
rect 36872 14980 37596 15008
rect 36872 14968 36878 14980
rect 36228 14912 36400 14940
rect 36228 14900 36234 14912
rect 36446 14900 36452 14952
rect 36504 14940 36510 14952
rect 36541 14943 36599 14949
rect 36541 14940 36553 14943
rect 36504 14912 36553 14940
rect 36504 14900 36510 14912
rect 36541 14909 36553 14912
rect 36587 14909 36599 14943
rect 36541 14903 36599 14909
rect 36630 14900 36636 14952
rect 36688 14940 36694 14952
rect 36909 14943 36967 14949
rect 36909 14940 36921 14943
rect 36688 14912 36921 14940
rect 36688 14900 36694 14912
rect 36909 14909 36921 14912
rect 36955 14909 36967 14943
rect 36909 14903 36967 14909
rect 37182 14900 37188 14952
rect 37240 14940 37246 14952
rect 37461 14943 37519 14949
rect 37461 14940 37473 14943
rect 37240 14912 37473 14940
rect 37240 14900 37246 14912
rect 37461 14909 37473 14912
rect 37507 14909 37519 14943
rect 37568 14940 37596 14980
rect 37642 14968 37648 15020
rect 37700 15008 37706 15020
rect 39114 15008 39120 15020
rect 37700 14980 37745 15008
rect 37844 14980 39120 15008
rect 37700 14968 37706 14980
rect 37844 14940 37872 14980
rect 39114 14968 39120 14980
rect 39172 14968 39178 15020
rect 39209 15011 39267 15017
rect 39209 14977 39221 15011
rect 39255 15008 39267 15011
rect 39408 15008 39436 15036
rect 39255 14980 39436 15008
rect 40589 15011 40647 15017
rect 39255 14977 39267 14980
rect 39209 14971 39267 14977
rect 40589 14977 40601 15011
rect 40635 14977 40647 15011
rect 40589 14971 40647 14977
rect 37568 14912 37872 14940
rect 37461 14903 37519 14909
rect 38102 14900 38108 14952
rect 38160 14940 38166 14952
rect 38160 14912 39059 14940
rect 38160 14900 38166 14912
rect 37829 14875 37887 14881
rect 37829 14872 37841 14875
rect 36004 14844 37841 14872
rect 37829 14841 37841 14844
rect 37875 14841 37887 14875
rect 38746 14872 38752 14884
rect 37829 14835 37887 14841
rect 38626 14844 38752 14872
rect 35069 14807 35127 14813
rect 35069 14804 35081 14807
rect 31628 14776 35081 14804
rect 31628 14764 31634 14776
rect 35069 14773 35081 14776
rect 35115 14773 35127 14807
rect 35069 14767 35127 14773
rect 35529 14807 35587 14813
rect 35529 14773 35541 14807
rect 35575 14804 35587 14807
rect 38626 14804 38654 14844
rect 38746 14832 38752 14844
rect 38804 14832 38810 14884
rect 39031 14872 39059 14912
rect 39298 14900 39304 14952
rect 39356 14940 39362 14952
rect 39485 14943 39543 14949
rect 39356 14912 39401 14940
rect 39356 14900 39362 14912
rect 39485 14909 39497 14943
rect 39531 14940 39543 14943
rect 39531 14912 39620 14940
rect 39531 14909 39543 14912
rect 39485 14903 39543 14909
rect 39592 14872 39620 14912
rect 40604 14872 40632 14971
rect 39031 14844 39620 14872
rect 39684 14844 40632 14872
rect 38838 14804 38844 14816
rect 35575 14776 38654 14804
rect 38799 14776 38844 14804
rect 35575 14773 35587 14776
rect 35529 14767 35587 14773
rect 38838 14764 38844 14776
rect 38896 14764 38902 14816
rect 39206 14764 39212 14816
rect 39264 14804 39270 14816
rect 39684 14804 39712 14844
rect 39264 14776 39712 14804
rect 39264 14764 39270 14776
rect 40310 14764 40316 14816
rect 40368 14804 40374 14816
rect 40586 14804 40592 14816
rect 40368 14776 40592 14804
rect 40368 14764 40374 14776
rect 40586 14764 40592 14776
rect 40644 14764 40650 14816
rect 40770 14764 40776 14816
rect 40828 14804 40834 14816
rect 42260 14804 42288 15048
rect 42334 14968 42340 15020
rect 42392 15008 42398 15020
rect 42889 15011 42947 15017
rect 42392 14980 42840 15008
rect 42392 14968 42398 14980
rect 42610 14900 42616 14952
rect 42668 14940 42674 14952
rect 42705 14943 42763 14949
rect 42705 14940 42717 14943
rect 42668 14912 42717 14940
rect 42668 14900 42674 14912
rect 42705 14909 42717 14912
rect 42751 14909 42763 14943
rect 42812 14940 42840 14980
rect 42889 14977 42901 15011
rect 42935 15008 42947 15011
rect 43438 15008 43444 15020
rect 42935 14980 43444 15008
rect 42935 14977 42947 14980
rect 42889 14971 42947 14977
rect 43438 14968 43444 14980
rect 43496 14968 43502 15020
rect 43622 15008 43628 15020
rect 43583 14980 43628 15008
rect 43622 14968 43628 14980
rect 43680 14968 43686 15020
rect 43993 15011 44051 15017
rect 43993 14977 44005 15011
rect 44039 15008 44051 15011
rect 44082 15008 44088 15020
rect 44039 14980 44088 15008
rect 44039 14977 44051 14980
rect 43993 14971 44051 14977
rect 44082 14968 44088 14980
rect 44140 14968 44146 15020
rect 44174 14968 44180 15020
rect 44232 15008 44238 15020
rect 44726 15017 44732 15020
rect 44453 15011 44511 15017
rect 44453 15008 44465 15011
rect 44232 14980 44465 15008
rect 44232 14968 44238 14980
rect 44453 14977 44465 14980
rect 44499 14977 44511 15011
rect 44453 14971 44511 14977
rect 44720 14971 44732 15017
rect 44784 15008 44790 15020
rect 44784 14980 44820 15008
rect 44726 14968 44732 14971
rect 44784 14968 44790 14980
rect 45462 14968 45468 15020
rect 45520 15008 45526 15020
rect 46293 15011 46351 15017
rect 46293 15008 46305 15011
rect 45520 14980 46305 15008
rect 45520 14968 45526 14980
rect 46293 14977 46305 14980
rect 46339 14977 46351 15011
rect 46400 15008 46428 15048
rect 46569 15045 46581 15079
rect 46615 15076 46627 15079
rect 46658 15076 46664 15088
rect 46615 15048 46664 15076
rect 46615 15045 46627 15048
rect 46569 15039 46627 15045
rect 46658 15036 46664 15048
rect 46716 15076 46722 15088
rect 47486 15076 47492 15088
rect 46716 15048 47492 15076
rect 46716 15036 46722 15048
rect 47486 15036 47492 15048
rect 47544 15076 47550 15088
rect 48222 15076 48228 15088
rect 47544 15048 48228 15076
rect 47544 15036 47550 15048
rect 48222 15036 48228 15048
rect 48280 15036 48286 15088
rect 48676 15079 48734 15085
rect 48676 15045 48688 15079
rect 48722 15076 48734 15079
rect 50706 15076 50712 15088
rect 48722 15048 50712 15076
rect 48722 15045 48734 15048
rect 48676 15039 48734 15045
rect 50706 15036 50712 15048
rect 50764 15036 50770 15088
rect 51046 15008 51074 15116
rect 55858 15008 55864 15020
rect 46400 14980 49464 15008
rect 51046 14980 55864 15008
rect 46293 14971 46351 14977
rect 48409 14943 48467 14949
rect 42812 14912 43852 14940
rect 42705 14903 42763 14909
rect 42720 14872 42748 14903
rect 43714 14872 43720 14884
rect 42720 14844 43720 14872
rect 43714 14832 43720 14844
rect 43772 14832 43778 14884
rect 40828 14776 42288 14804
rect 43824 14804 43852 14912
rect 48409 14909 48421 14943
rect 48455 14909 48467 14943
rect 49436 14940 49464 14980
rect 55858 14968 55864 14980
rect 55916 14968 55922 15020
rect 57606 14940 57612 14952
rect 49436 14912 57612 14940
rect 48409 14903 48467 14909
rect 47118 14804 47124 14816
rect 43824 14776 47124 14804
rect 40828 14764 40834 14776
rect 47118 14764 47124 14776
rect 47176 14764 47182 14816
rect 48424 14804 48452 14903
rect 57606 14900 57612 14912
rect 57664 14900 57670 14952
rect 49786 14872 49792 14884
rect 49699 14844 49792 14872
rect 49786 14832 49792 14844
rect 49844 14872 49850 14884
rect 50982 14872 50988 14884
rect 49844 14844 50988 14872
rect 49844 14832 49850 14844
rect 50982 14832 50988 14844
rect 51040 14832 51046 14884
rect 49694 14804 49700 14816
rect 48424 14776 49700 14804
rect 49694 14764 49700 14776
rect 49752 14764 49758 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 10965 14603 11023 14609
rect 10965 14569 10977 14603
rect 11011 14600 11023 14603
rect 11422 14600 11428 14612
rect 11011 14572 11428 14600
rect 11011 14569 11023 14572
rect 10965 14563 11023 14569
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 24578 14600 24584 14612
rect 13504 14572 24440 14600
rect 24539 14572 24584 14600
rect 13504 14560 13510 14572
rect 20809 14535 20867 14541
rect 20809 14501 20821 14535
rect 20855 14501 20867 14535
rect 20809 14495 20867 14501
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 10643 14436 12541 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14461 14467 14519 14473
rect 14461 14464 14473 14467
rect 13964 14436 14473 14464
rect 13964 14424 13970 14436
rect 14461 14433 14473 14436
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14464 14795 14467
rect 15194 14464 15200 14476
rect 14783 14436 15200 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 15988 14436 16712 14464
rect 15988 14424 15994 14436
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 8938 14396 8944 14408
rect 1627 14368 8944 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 10778 14396 10784 14408
rect 10739 14368 10784 14396
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14396 11483 14399
rect 11606 14396 11612 14408
rect 11471 14368 11612 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 13780 14368 16589 14396
rect 13780 14356 13786 14368
rect 16577 14365 16589 14368
rect 16623 14365 16635 14399
rect 16684 14396 16712 14436
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 19426 14464 19432 14476
rect 16908 14436 19432 14464
rect 16908 14424 16914 14436
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 20824 14464 20852 14495
rect 20898 14492 20904 14544
rect 20956 14532 20962 14544
rect 22094 14532 22100 14544
rect 20956 14504 22100 14532
rect 20956 14492 20962 14504
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 24302 14532 24308 14544
rect 22572 14504 24308 14532
rect 22572 14464 22600 14504
rect 24302 14492 24308 14504
rect 24360 14492 24366 14544
rect 24412 14532 24440 14572
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 25590 14560 25596 14612
rect 25648 14600 25654 14612
rect 25648 14572 30696 14600
rect 25648 14560 25654 14572
rect 24412 14504 25360 14532
rect 20824 14436 22600 14464
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 25332 14464 25360 14504
rect 26602 14492 26608 14544
rect 26660 14532 26666 14544
rect 28077 14535 28135 14541
rect 28077 14532 28089 14535
rect 26660 14504 28089 14532
rect 26660 14492 26666 14504
rect 28077 14501 28089 14504
rect 28123 14501 28135 14535
rect 30668 14532 30696 14572
rect 30742 14560 30748 14612
rect 30800 14600 30806 14612
rect 32953 14603 33011 14609
rect 32953 14600 32965 14603
rect 30800 14572 32965 14600
rect 30800 14560 30806 14572
rect 32953 14569 32965 14572
rect 32999 14569 33011 14603
rect 32953 14563 33011 14569
rect 34698 14560 34704 14612
rect 34756 14600 34762 14612
rect 34977 14603 35035 14609
rect 34977 14600 34989 14603
rect 34756 14572 34989 14600
rect 34756 14560 34762 14572
rect 34977 14569 34989 14572
rect 35023 14569 35035 14603
rect 34977 14563 35035 14569
rect 36170 14560 36176 14612
rect 36228 14600 36234 14612
rect 37090 14600 37096 14612
rect 36228 14572 37096 14600
rect 36228 14560 36234 14572
rect 37090 14560 37096 14572
rect 37148 14560 37154 14612
rect 37550 14560 37556 14612
rect 37608 14600 37614 14612
rect 42334 14600 42340 14612
rect 37608 14572 42340 14600
rect 37608 14560 37614 14572
rect 42334 14560 42340 14572
rect 42392 14560 42398 14612
rect 42702 14600 42708 14612
rect 42663 14572 42708 14600
rect 42702 14560 42708 14572
rect 42760 14560 42766 14612
rect 46750 14600 46756 14612
rect 46711 14572 46756 14600
rect 46750 14560 46756 14572
rect 46808 14560 46814 14612
rect 48593 14603 48651 14609
rect 48593 14600 48605 14603
rect 46952 14572 48605 14600
rect 30926 14532 30932 14544
rect 30668 14504 30932 14532
rect 28077 14495 28135 14501
rect 30926 14492 30932 14504
rect 30984 14492 30990 14544
rect 31110 14532 31116 14544
rect 31071 14504 31116 14532
rect 31110 14492 31116 14504
rect 31168 14492 31174 14544
rect 33781 14535 33839 14541
rect 33781 14501 33793 14535
rect 33827 14532 33839 14535
rect 33870 14532 33876 14544
rect 33827 14504 33876 14532
rect 33827 14501 33839 14504
rect 33781 14495 33839 14501
rect 33870 14492 33876 14504
rect 33928 14492 33934 14544
rect 34238 14492 34244 14544
rect 34296 14532 34302 14544
rect 36081 14535 36139 14541
rect 34296 14504 36032 14532
rect 34296 14492 34302 14504
rect 28350 14464 28356 14476
rect 22704 14436 24891 14464
rect 25332 14436 28356 14464
rect 22704 14424 22710 14436
rect 21729 14399 21787 14405
rect 16684 14368 21680 14396
rect 16577 14359 16635 14365
rect 1854 14328 1860 14340
rect 1815 14300 1860 14328
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 18877 14331 18935 14337
rect 18877 14297 18889 14331
rect 18923 14328 18935 14331
rect 19674 14331 19732 14337
rect 19674 14328 19686 14331
rect 18923 14300 19686 14328
rect 18923 14297 18935 14300
rect 18877 14291 18935 14297
rect 19674 14297 19686 14300
rect 19720 14297 19732 14331
rect 21652 14328 21680 14368
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 22830 14396 22836 14408
rect 21775 14368 22836 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 23106 14356 23112 14408
rect 23164 14396 23170 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 23164 14368 24593 14396
rect 23164 14356 23170 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24581 14359 24639 14365
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 24863 14396 24891 14436
rect 28350 14424 28356 14436
rect 28408 14424 28414 14476
rect 28534 14464 28540 14476
rect 28495 14436 28540 14464
rect 28534 14424 28540 14436
rect 28592 14424 28598 14476
rect 28721 14467 28779 14473
rect 28721 14433 28733 14467
rect 28767 14464 28779 14467
rect 29362 14464 29368 14476
rect 28767 14436 29368 14464
rect 28767 14433 28779 14436
rect 28721 14427 28779 14433
rect 29362 14424 29368 14436
rect 29420 14424 29426 14476
rect 33965 14467 34023 14473
rect 33965 14464 33977 14467
rect 33888 14436 33977 14464
rect 33888 14408 33916 14436
rect 33965 14433 33977 14436
rect 34011 14433 34023 14467
rect 33965 14427 34023 14433
rect 34149 14467 34207 14473
rect 34149 14433 34161 14467
rect 34195 14464 34207 14467
rect 34330 14464 34336 14476
rect 34195 14436 34336 14464
rect 34195 14433 34207 14436
rect 34149 14427 34207 14433
rect 34330 14424 34336 14436
rect 34388 14424 34394 14476
rect 34698 14424 34704 14476
rect 34756 14464 34762 14476
rect 35529 14467 35587 14473
rect 35529 14464 35541 14467
rect 34756 14436 35541 14464
rect 34756 14424 34762 14436
rect 25317 14399 25375 14405
rect 25317 14396 25329 14399
rect 24863 14368 25329 14396
rect 25317 14365 25329 14368
rect 25363 14396 25375 14399
rect 25363 14368 25452 14396
rect 25363 14365 25375 14368
rect 25317 14359 25375 14365
rect 25424 14328 25452 14368
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 28445 14399 28503 14405
rect 28445 14396 28457 14399
rect 25556 14368 28457 14396
rect 25556 14356 25562 14368
rect 28445 14365 28457 14368
rect 28491 14365 28503 14399
rect 28445 14359 28503 14365
rect 29733 14399 29791 14405
rect 29733 14365 29745 14399
rect 29779 14396 29791 14399
rect 29822 14396 29828 14408
rect 29779 14368 29828 14396
rect 29779 14365 29791 14368
rect 29733 14359 29791 14365
rect 29822 14356 29828 14368
rect 29880 14396 29886 14408
rect 31573 14399 31631 14405
rect 31573 14396 31585 14399
rect 29880 14368 31585 14396
rect 29880 14356 29886 14368
rect 31573 14365 31585 14368
rect 31619 14365 31631 14399
rect 31573 14359 31631 14365
rect 33870 14356 33876 14408
rect 33928 14356 33934 14408
rect 34057 14399 34115 14405
rect 34057 14365 34069 14399
rect 34103 14365 34115 14399
rect 34057 14359 34115 14365
rect 34241 14399 34299 14405
rect 34241 14365 34253 14399
rect 34287 14396 34299 14399
rect 34790 14396 34796 14408
rect 34287 14368 34796 14396
rect 34287 14365 34299 14368
rect 34241 14359 34299 14365
rect 25590 14328 25596 14340
rect 21652 14300 23060 14328
rect 25424 14300 25596 14328
rect 19674 14291 19732 14297
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 13078 14260 13084 14272
rect 11020 14232 13084 14260
rect 11020 14220 11026 14232
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 15838 14260 15844 14272
rect 15799 14232 15844 14260
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16022 14220 16028 14272
rect 16080 14260 16086 14272
rect 17126 14260 17132 14272
rect 16080 14232 17132 14260
rect 16080 14220 16086 14232
rect 17126 14220 17132 14232
rect 17184 14260 17190 14272
rect 22925 14263 22983 14269
rect 22925 14260 22937 14263
rect 17184 14232 22937 14260
rect 17184 14220 17190 14232
rect 22925 14229 22937 14232
rect 22971 14229 22983 14263
rect 23032 14260 23060 14300
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 30006 14337 30012 14340
rect 30000 14328 30012 14337
rect 29967 14300 30012 14328
rect 30000 14291 30012 14300
rect 30006 14288 30012 14291
rect 30064 14288 30070 14340
rect 31294 14288 31300 14340
rect 31352 14328 31358 14340
rect 31818 14331 31876 14337
rect 31818 14328 31830 14331
rect 31352 14300 31830 14328
rect 31352 14288 31358 14300
rect 31818 14297 31830 14300
rect 31864 14297 31876 14331
rect 31818 14291 31876 14297
rect 33962 14288 33968 14340
rect 34020 14328 34026 14340
rect 34072 14328 34100 14359
rect 34790 14356 34796 14368
rect 34848 14356 34854 14408
rect 35158 14399 35216 14405
rect 35158 14365 35170 14399
rect 35204 14365 35216 14399
rect 35158 14359 35216 14365
rect 35452 14390 35480 14436
rect 35529 14433 35541 14436
rect 35575 14433 35587 14467
rect 35529 14427 35587 14433
rect 35621 14467 35679 14473
rect 35621 14433 35633 14467
rect 35667 14464 35679 14467
rect 35710 14464 35716 14476
rect 35667 14436 35716 14464
rect 35667 14433 35679 14436
rect 35621 14427 35679 14433
rect 35710 14424 35716 14436
rect 35768 14424 35774 14476
rect 35897 14467 35955 14473
rect 35897 14433 35909 14467
rect 35943 14433 35955 14467
rect 36004 14464 36032 14504
rect 36081 14501 36093 14535
rect 36127 14532 36139 14535
rect 36630 14532 36636 14544
rect 36127 14504 36636 14532
rect 36127 14501 36139 14504
rect 36081 14495 36139 14501
rect 36630 14492 36636 14504
rect 36688 14492 36694 14544
rect 37182 14492 37188 14544
rect 37240 14532 37246 14544
rect 37461 14535 37519 14541
rect 37461 14532 37473 14535
rect 37240 14504 37473 14532
rect 37240 14492 37246 14504
rect 37461 14501 37473 14504
rect 37507 14501 37519 14535
rect 37461 14495 37519 14501
rect 40037 14535 40095 14541
rect 40037 14501 40049 14535
rect 40083 14532 40095 14535
rect 41322 14532 41328 14544
rect 40083 14504 41328 14532
rect 40083 14501 40095 14504
rect 40037 14495 40095 14501
rect 41322 14492 41328 14504
rect 41380 14492 41386 14544
rect 41414 14492 41420 14544
rect 41472 14532 41478 14544
rect 41472 14504 44036 14532
rect 41472 14492 41478 14504
rect 38010 14464 38016 14476
rect 36004 14436 36207 14464
rect 37971 14436 38016 14464
rect 35897 14427 35955 14433
rect 35912 14396 35940 14427
rect 35636 14390 35940 14396
rect 35452 14368 35940 14390
rect 36179 14398 36207 14436
rect 38010 14424 38016 14436
rect 38068 14424 38074 14476
rect 39206 14424 39212 14476
rect 39264 14464 39270 14476
rect 40681 14467 40739 14473
rect 39264 14436 40356 14464
rect 39264 14424 39270 14436
rect 36268 14399 36326 14405
rect 36268 14398 36280 14399
rect 36179 14370 36280 14398
rect 35452 14362 35664 14368
rect 36268 14365 36280 14370
rect 36314 14365 36326 14399
rect 36268 14359 36326 14365
rect 34020 14300 34100 14328
rect 35173 14328 35201 14359
rect 36354 14356 36360 14408
rect 36412 14356 36418 14408
rect 37185 14399 37243 14405
rect 37185 14365 37197 14399
rect 37231 14365 37243 14399
rect 37185 14359 37243 14365
rect 37297 14399 37355 14405
rect 37297 14365 37309 14399
rect 37343 14396 37355 14399
rect 37734 14396 37740 14408
rect 37343 14368 37740 14396
rect 37343 14365 37355 14368
rect 37297 14359 37355 14365
rect 36170 14328 36176 14340
rect 35173 14300 36176 14328
rect 34020 14288 34026 14300
rect 36170 14288 36176 14300
rect 36228 14288 36234 14340
rect 36372 14328 36400 14356
rect 36630 14328 36636 14340
rect 36372 14300 36492 14328
rect 36591 14300 36636 14328
rect 26513 14263 26571 14269
rect 26513 14260 26525 14263
rect 23032 14232 26525 14260
rect 22925 14223 22983 14229
rect 26513 14229 26525 14232
rect 26559 14229 26571 14263
rect 26513 14223 26571 14229
rect 35161 14263 35219 14269
rect 35161 14229 35173 14263
rect 35207 14260 35219 14263
rect 35618 14260 35624 14272
rect 35207 14232 35624 14260
rect 35207 14229 35219 14232
rect 35161 14223 35219 14229
rect 35618 14220 35624 14232
rect 35676 14260 35682 14272
rect 36078 14260 36084 14272
rect 35676 14232 36084 14260
rect 35676 14220 35682 14232
rect 36078 14220 36084 14232
rect 36136 14220 36142 14272
rect 36262 14220 36268 14272
rect 36320 14260 36326 14272
rect 36464 14269 36492 14300
rect 36630 14288 36636 14300
rect 36688 14288 36694 14340
rect 36357 14263 36415 14269
rect 36357 14260 36369 14263
rect 36320 14232 36369 14260
rect 36320 14220 36326 14232
rect 36357 14229 36369 14232
rect 36403 14229 36415 14263
rect 36357 14223 36415 14229
rect 36449 14263 36507 14269
rect 36449 14229 36461 14263
rect 36495 14229 36507 14263
rect 37200 14260 37228 14359
rect 37734 14356 37740 14368
rect 37792 14356 37798 14408
rect 38280 14399 38338 14405
rect 38280 14365 38292 14399
rect 38326 14396 38338 14399
rect 38838 14396 38844 14408
rect 38326 14368 38844 14396
rect 38326 14365 38338 14368
rect 38280 14359 38338 14365
rect 38838 14356 38844 14368
rect 38896 14356 38902 14408
rect 40218 14396 40224 14408
rect 40179 14368 40224 14396
rect 40218 14356 40224 14368
rect 40276 14356 40282 14408
rect 40328 14405 40356 14436
rect 40681 14433 40693 14467
rect 40727 14464 40739 14467
rect 40770 14464 40776 14476
rect 40727 14436 40776 14464
rect 40727 14433 40739 14436
rect 40681 14427 40739 14433
rect 40770 14424 40776 14436
rect 40828 14424 40834 14476
rect 41506 14464 41512 14476
rect 41064 14436 41512 14464
rect 40313 14399 40371 14405
rect 40313 14365 40325 14399
rect 40359 14365 40371 14399
rect 40313 14359 40371 14365
rect 40405 14399 40463 14405
rect 40405 14365 40417 14399
rect 40451 14396 40463 14399
rect 41064 14396 41092 14436
rect 41506 14424 41512 14436
rect 41564 14424 41570 14476
rect 42444 14436 43668 14464
rect 41230 14396 41236 14408
rect 40451 14368 41092 14396
rect 41191 14368 41236 14396
rect 40451 14365 40463 14368
rect 40405 14359 40463 14365
rect 41230 14356 41236 14368
rect 41288 14356 41294 14408
rect 41322 14356 41328 14408
rect 41380 14396 41386 14408
rect 41380 14368 41425 14396
rect 41616 14368 41828 14396
rect 41380 14356 41386 14368
rect 37458 14288 37464 14340
rect 37516 14328 37522 14340
rect 38746 14328 38752 14340
rect 37516 14300 38752 14328
rect 37516 14288 37522 14300
rect 38746 14288 38752 14300
rect 38804 14288 38810 14340
rect 40586 14337 40592 14340
rect 40543 14331 40592 14337
rect 40543 14297 40555 14331
rect 40589 14297 40592 14331
rect 40543 14291 40592 14297
rect 40586 14288 40592 14291
rect 40644 14288 40650 14340
rect 41046 14288 41052 14340
rect 41104 14328 41110 14340
rect 41616 14328 41644 14368
rect 41104 14300 41644 14328
rect 41800 14328 41828 14368
rect 41874 14356 41880 14408
rect 41932 14396 41938 14408
rect 42061 14399 42119 14405
rect 42061 14396 42073 14399
rect 41932 14368 42073 14396
rect 41932 14356 41938 14368
rect 42061 14365 42073 14368
rect 42107 14365 42119 14399
rect 42061 14359 42119 14365
rect 42209 14399 42267 14405
rect 42209 14365 42221 14399
rect 42255 14396 42267 14399
rect 42444 14396 42472 14436
rect 42255 14368 42472 14396
rect 42526 14399 42584 14405
rect 42255 14365 42267 14368
rect 42209 14359 42267 14365
rect 42526 14365 42538 14399
rect 42572 14398 42584 14399
rect 42572 14396 42656 14398
rect 42702 14396 42708 14408
rect 42572 14370 42708 14396
rect 42572 14365 42584 14370
rect 42628 14368 42708 14370
rect 42526 14359 42584 14365
rect 42702 14356 42708 14368
rect 42760 14356 42766 14408
rect 43254 14396 43260 14408
rect 43215 14368 43260 14396
rect 43254 14356 43260 14368
rect 43312 14356 43318 14408
rect 42337 14331 42395 14337
rect 42337 14328 42349 14331
rect 41800 14300 42349 14328
rect 41104 14288 41110 14300
rect 42337 14297 42349 14300
rect 42383 14297 42395 14331
rect 42337 14291 42395 14297
rect 42429 14331 42487 14337
rect 42429 14297 42441 14331
rect 42475 14328 42487 14331
rect 43346 14328 43352 14340
rect 42475 14300 43352 14328
rect 42475 14297 42487 14300
rect 42429 14291 42487 14297
rect 43346 14288 43352 14300
rect 43404 14288 43410 14340
rect 43640 14328 43668 14436
rect 43806 14356 43812 14408
rect 43864 14396 43870 14408
rect 44008 14405 44036 14504
rect 44082 14492 44088 14544
rect 44140 14532 44146 14544
rect 44818 14532 44824 14544
rect 44140 14504 44824 14532
rect 44140 14492 44146 14504
rect 44818 14492 44824 14504
rect 44876 14492 44882 14544
rect 44450 14464 44456 14476
rect 44284 14436 44456 14464
rect 43993 14399 44051 14405
rect 43864 14368 43944 14396
rect 43864 14356 43870 14368
rect 43916 14328 43944 14368
rect 43993 14365 44005 14399
rect 44039 14365 44051 14399
rect 44174 14396 44180 14408
rect 44135 14368 44180 14396
rect 43993 14359 44051 14365
rect 44174 14356 44180 14368
rect 44232 14356 44238 14408
rect 44284 14405 44312 14436
rect 44450 14424 44456 14436
rect 44508 14424 44514 14476
rect 46750 14424 46756 14476
rect 46808 14464 46814 14476
rect 46952 14464 46980 14572
rect 48593 14569 48605 14572
rect 48639 14600 48651 14603
rect 56502 14600 56508 14612
rect 48639 14572 56508 14600
rect 48639 14569 48651 14572
rect 48593 14563 48651 14569
rect 56502 14560 56508 14572
rect 56560 14560 56566 14612
rect 46808 14436 46980 14464
rect 46808 14424 46814 14436
rect 44269 14399 44327 14405
rect 44269 14365 44281 14399
rect 44315 14365 44327 14399
rect 44269 14359 44327 14365
rect 44361 14399 44419 14405
rect 44361 14365 44373 14399
rect 44407 14365 44419 14399
rect 44361 14359 44419 14365
rect 45373 14399 45431 14405
rect 45373 14365 45385 14399
rect 45419 14396 45431 14399
rect 45462 14396 45468 14408
rect 45419 14368 45468 14396
rect 45419 14365 45431 14368
rect 45373 14359 45431 14365
rect 44376 14328 44404 14359
rect 45462 14356 45468 14368
rect 45520 14396 45526 14408
rect 47213 14399 47271 14405
rect 47213 14396 47225 14399
rect 45520 14368 47225 14396
rect 45520 14356 45526 14368
rect 47213 14365 47225 14368
rect 47259 14365 47271 14399
rect 57974 14396 57980 14408
rect 57935 14368 57980 14396
rect 47213 14359 47271 14365
rect 57974 14356 57980 14368
rect 58032 14356 58038 14408
rect 43640 14300 43852 14328
rect 43916 14300 44404 14328
rect 38654 14260 38660 14272
rect 37200 14232 38660 14260
rect 36449 14223 36507 14229
rect 38654 14220 38660 14232
rect 38712 14220 38718 14272
rect 39390 14260 39396 14272
rect 39351 14232 39396 14260
rect 39390 14220 39396 14232
rect 39448 14220 39454 14272
rect 39666 14220 39672 14272
rect 39724 14260 39730 14272
rect 41509 14263 41567 14269
rect 41509 14260 41521 14263
rect 39724 14232 41521 14260
rect 39724 14220 39730 14232
rect 41509 14229 41521 14232
rect 41555 14229 41567 14263
rect 41509 14223 41567 14229
rect 43441 14263 43499 14269
rect 43441 14229 43453 14263
rect 43487 14260 43499 14263
rect 43714 14260 43720 14272
rect 43487 14232 43720 14260
rect 43487 14229 43499 14232
rect 43441 14223 43499 14229
rect 43714 14220 43720 14232
rect 43772 14220 43778 14272
rect 43824 14260 43852 14300
rect 44450 14288 44456 14340
rect 44508 14328 44514 14340
rect 45640 14331 45698 14337
rect 44508 14300 45600 14328
rect 44508 14288 44514 14300
rect 44358 14260 44364 14272
rect 43824 14232 44364 14260
rect 44358 14220 44364 14232
rect 44416 14220 44422 14272
rect 44545 14263 44603 14269
rect 44545 14229 44557 14263
rect 44591 14260 44603 14263
rect 44818 14260 44824 14272
rect 44591 14232 44824 14260
rect 44591 14229 44603 14232
rect 44545 14223 44603 14229
rect 44818 14220 44824 14232
rect 44876 14220 44882 14272
rect 45572 14260 45600 14300
rect 45640 14297 45652 14331
rect 45686 14328 45698 14331
rect 46566 14328 46572 14340
rect 45686 14300 46572 14328
rect 45686 14297 45698 14300
rect 45640 14291 45698 14297
rect 46566 14288 46572 14300
rect 46624 14288 46630 14340
rect 47480 14331 47538 14337
rect 47480 14297 47492 14331
rect 47526 14328 47538 14331
rect 48130 14328 48136 14340
rect 47526 14300 48136 14328
rect 47526 14297 47538 14300
rect 47480 14291 47538 14297
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 46842 14260 46848 14272
rect 45572 14232 46848 14260
rect 46842 14220 46848 14232
rect 46900 14220 46906 14272
rect 58066 14260 58072 14272
rect 58027 14232 58072 14260
rect 58066 14220 58072 14232
rect 58124 14220 58130 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 11054 14056 11060 14068
rect 10520 14028 11060 14056
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 2424 13920 2452 14016
rect 1627 13892 2452 13920
rect 10045 13923 10103 13929
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10520 13920 10548 14028
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 12434 14056 12440 14068
rect 11195 14028 12440 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 15930 14056 15936 14068
rect 13004 14028 15936 14056
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 12158 13988 12164 14000
rect 10744 13960 12164 13988
rect 10744 13948 10750 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 12250 13920 12256 13932
rect 10091 13892 10548 13920
rect 12211 13892 12256 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 13004 13920 13032 14028
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14056 16267 14059
rect 17218 14056 17224 14068
rect 16255 14028 17224 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 28353 14059 28411 14065
rect 28353 14056 28365 14059
rect 17460 14028 28365 14056
rect 17460 14016 17466 14028
rect 28353 14025 28365 14028
rect 28399 14025 28411 14059
rect 28353 14019 28411 14025
rect 31297 14059 31355 14065
rect 31297 14025 31309 14059
rect 31343 14025 31355 14059
rect 36262 14056 36268 14068
rect 31297 14019 31355 14025
rect 31404 14028 36268 14056
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 22732 13991 22790 13997
rect 13136 13960 16988 13988
rect 13136 13948 13142 13960
rect 12483 13892 13032 13920
rect 13173 13923 13231 13929
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13538 13920 13544 13932
rect 13219 13892 13544 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 15286 13920 15292 13932
rect 14047 13892 15292 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 16482 13920 16488 13932
rect 16264 13892 16488 13920
rect 16264 13880 16270 13892
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 16960 13920 16988 13960
rect 22732 13957 22744 13991
rect 22778 13988 22790 13991
rect 26786 13988 26792 14000
rect 22778 13960 26792 13988
rect 22778 13957 22790 13960
rect 22732 13951 22790 13957
rect 26786 13948 26792 13960
rect 26844 13948 26850 14000
rect 30006 13988 30012 14000
rect 27172 13960 30012 13988
rect 19153 13923 19211 13929
rect 19153 13920 19165 13923
rect 16960 13892 19165 13920
rect 19153 13889 19165 13892
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 24302 13920 24308 13932
rect 19300 13892 23520 13920
rect 24263 13892 24308 13920
rect 19300 13880 19306 13892
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 11422 13852 11428 13864
rect 9907 13824 11428 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 11974 13852 11980 13864
rect 11935 13824 11980 13852
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 12124 13824 12173 13852
rect 12124 13812 12130 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13852 12403 13855
rect 12526 13852 12532 13864
rect 12391 13824 12532 13852
rect 12391 13821 12403 13824
rect 12345 13815 12403 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12676 13824 13277 13852
rect 12676 13812 12682 13824
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 14792 13824 17141 13852
rect 14792 13812 14798 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13852 21511 13855
rect 22186 13852 22192 13864
rect 21499 13824 22192 13852
rect 21499 13821 21511 13824
rect 21453 13815 21511 13821
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22462 13852 22468 13864
rect 22423 13824 22468 13852
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 7892 13756 10977 13784
rect 7892 13744 7898 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 10965 13747 11023 13753
rect 13541 13787 13599 13793
rect 13541 13753 13553 13787
rect 13587 13784 13599 13787
rect 13722 13784 13728 13796
rect 13587 13756 13728 13784
rect 13587 13753 13599 13756
rect 13541 13747 13599 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13906 13744 13912 13796
rect 13964 13784 13970 13796
rect 16022 13784 16028 13796
rect 13964 13756 16028 13784
rect 13964 13744 13970 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18104 13756 18460 13784
rect 18104 13744 18110 13756
rect 10042 13676 10048 13728
rect 10100 13716 10106 13728
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 10100 13688 10241 13716
rect 10100 13676 10106 13688
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 14458 13716 14464 13728
rect 12952 13688 14464 13716
rect 12952 13676 12958 13688
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 18230 13716 18236 13728
rect 14700 13688 18236 13716
rect 14700 13676 14706 13688
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18432 13725 18460 13756
rect 21818 13744 21824 13796
rect 21876 13784 21882 13796
rect 22370 13784 22376 13796
rect 21876 13756 22376 13784
rect 21876 13744 21882 13756
rect 22370 13744 22376 13756
rect 22428 13744 22434 13796
rect 23492 13784 23520 13892
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 25222 13880 25228 13932
rect 25280 13920 25286 13932
rect 27172 13929 27200 13960
rect 30006 13948 30012 13960
rect 30064 13948 30070 14000
rect 30190 13997 30196 14000
rect 30184 13988 30196 13997
rect 30151 13960 30196 13988
rect 30184 13951 30196 13960
rect 30190 13948 30196 13951
rect 30248 13948 30254 14000
rect 31018 13948 31024 14000
rect 31076 13988 31082 14000
rect 31312 13988 31340 14019
rect 31076 13960 31340 13988
rect 31076 13948 31082 13960
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 25280 13892 27169 13920
rect 25280 13880 25286 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 29822 13880 29828 13932
rect 29880 13920 29886 13932
rect 29917 13923 29975 13929
rect 29917 13920 29929 13923
rect 29880 13892 29929 13920
rect 29880 13880 29886 13892
rect 29917 13889 29929 13892
rect 29963 13889 29975 13923
rect 31404 13920 31432 14028
rect 36262 14016 36268 14028
rect 36320 14016 36326 14068
rect 36357 14059 36415 14065
rect 36357 14025 36369 14059
rect 36403 14056 36415 14059
rect 37090 14056 37096 14068
rect 36403 14028 37096 14056
rect 36403 14025 36415 14028
rect 36357 14019 36415 14025
rect 37090 14016 37096 14028
rect 37148 14016 37154 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37645 14059 37703 14065
rect 37645 14056 37657 14059
rect 37424 14028 37657 14056
rect 37424 14016 37430 14028
rect 37645 14025 37657 14028
rect 37691 14025 37703 14059
rect 37645 14019 37703 14025
rect 38654 14016 38660 14068
rect 38712 14056 38718 14068
rect 38712 14028 40356 14056
rect 38712 14016 38718 14028
rect 34330 13948 34336 14000
rect 34388 13988 34394 14000
rect 39108 13991 39166 13997
rect 34388 13960 38976 13988
rect 34388 13948 34394 13960
rect 29917 13883 29975 13889
rect 30015 13892 31432 13920
rect 32861 13923 32919 13929
rect 29270 13812 29276 13864
rect 29328 13852 29334 13864
rect 30015 13852 30043 13892
rect 32861 13889 32873 13923
rect 32907 13920 32919 13923
rect 32950 13920 32956 13932
rect 32907 13892 32956 13920
rect 32907 13889 32919 13892
rect 32861 13883 32919 13889
rect 32950 13880 32956 13892
rect 33008 13880 33014 13932
rect 33137 13923 33195 13929
rect 33137 13889 33149 13923
rect 33183 13920 33195 13923
rect 34882 13920 34888 13932
rect 33183 13892 34888 13920
rect 33183 13889 33195 13892
rect 33137 13883 33195 13889
rect 34882 13880 34888 13892
rect 34940 13880 34946 13932
rect 35241 13929 35247 13932
rect 35233 13923 35247 13929
rect 35233 13920 35245 13923
rect 35202 13892 35245 13920
rect 35233 13889 35245 13892
rect 35233 13883 35247 13889
rect 35241 13880 35247 13883
rect 35299 13880 35305 13932
rect 37274 13880 37280 13932
rect 37332 13920 37338 13932
rect 37550 13920 37556 13932
rect 37332 13892 37556 13920
rect 37332 13880 37338 13892
rect 37550 13880 37556 13892
rect 37608 13880 37614 13932
rect 38010 13880 38016 13932
rect 38068 13920 38074 13932
rect 38841 13923 38899 13929
rect 38841 13920 38853 13923
rect 38068 13892 38853 13920
rect 38068 13880 38074 13892
rect 38841 13889 38853 13892
rect 38887 13889 38899 13923
rect 38948 13920 38976 13960
rect 39108 13957 39120 13991
rect 39154 13988 39166 13991
rect 39666 13988 39672 14000
rect 39154 13960 39672 13988
rect 39154 13957 39166 13960
rect 39108 13951 39166 13957
rect 39666 13948 39672 13960
rect 39724 13948 39730 14000
rect 40328 13988 40356 14028
rect 40402 14016 40408 14068
rect 40460 14056 40466 14068
rect 40770 14056 40776 14068
rect 40460 14028 40776 14056
rect 40460 14016 40466 14028
rect 40770 14016 40776 14028
rect 40828 14016 40834 14068
rect 41874 14056 41880 14068
rect 41340 14028 41736 14056
rect 41835 14028 41880 14056
rect 41230 13988 41236 14000
rect 40328 13960 41236 13988
rect 41230 13948 41236 13960
rect 41288 13948 41294 14000
rect 41046 13920 41052 13932
rect 38948 13892 41052 13920
rect 38841 13883 38899 13889
rect 41046 13880 41052 13892
rect 41104 13880 41110 13932
rect 41340 13929 41368 14028
rect 41598 13988 41604 14000
rect 41559 13960 41604 13988
rect 41598 13948 41604 13960
rect 41656 13948 41662 14000
rect 41708 13988 41736 14028
rect 41874 14016 41880 14028
rect 41932 14016 41938 14068
rect 43441 14059 43499 14065
rect 43441 14025 43453 14059
rect 43487 14056 43499 14059
rect 43622 14056 43628 14068
rect 43487 14028 43628 14056
rect 43487 14025 43499 14028
rect 43441 14019 43499 14025
rect 43622 14016 43628 14028
rect 43680 14016 43686 14068
rect 44726 14056 44732 14068
rect 44687 14028 44732 14056
rect 44726 14016 44732 14028
rect 44784 14016 44790 14068
rect 47213 14059 47271 14065
rect 47213 14025 47225 14059
rect 47259 14056 47271 14059
rect 48130 14056 48136 14068
rect 47259 14028 47900 14056
rect 48091 14028 48136 14056
rect 47259 14025 47271 14028
rect 47213 14019 47271 14025
rect 41708 13960 42288 13988
rect 41325 13923 41383 13929
rect 41325 13889 41337 13923
rect 41371 13889 41383 13923
rect 41325 13883 41383 13889
rect 41509 13923 41567 13929
rect 41509 13889 41521 13923
rect 41555 13889 41567 13923
rect 41509 13883 41567 13889
rect 41693 13923 41751 13929
rect 41693 13889 41705 13923
rect 41739 13889 41751 13923
rect 41693 13883 41751 13889
rect 29328 13824 30043 13852
rect 29328 13812 29334 13824
rect 30926 13812 30932 13864
rect 30984 13852 30990 13864
rect 33870 13852 33876 13864
rect 30984 13824 33876 13852
rect 30984 13812 30990 13824
rect 33870 13812 33876 13824
rect 33928 13852 33934 13864
rect 34241 13855 34299 13861
rect 34241 13852 34253 13855
rect 33928 13824 34253 13852
rect 33928 13812 33934 13824
rect 34241 13821 34253 13824
rect 34287 13821 34299 13855
rect 34241 13815 34299 13821
rect 34790 13812 34796 13864
rect 34848 13852 34854 13864
rect 34977 13855 35035 13861
rect 34977 13852 34989 13855
rect 34848 13824 34989 13852
rect 34848 13812 34854 13824
rect 34977 13821 34989 13824
rect 35023 13821 35035 13855
rect 34977 13815 35035 13821
rect 36078 13812 36084 13864
rect 36136 13852 36142 13864
rect 37458 13852 37464 13864
rect 36136 13824 37464 13852
rect 36136 13812 36142 13824
rect 37458 13812 37464 13824
rect 37516 13812 37522 13864
rect 40402 13852 40408 13864
rect 40236 13824 40408 13852
rect 28166 13784 28172 13796
rect 23492 13756 28172 13784
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 40236 13793 40264 13824
rect 40402 13812 40408 13824
rect 40460 13812 40466 13864
rect 40770 13812 40776 13864
rect 40828 13852 40834 13864
rect 41524 13852 41552 13883
rect 40828 13824 41552 13852
rect 40828 13812 40834 13824
rect 40221 13787 40279 13793
rect 35912 13756 36492 13784
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13716 18475 13719
rect 22646 13716 22652 13728
rect 18463 13688 22652 13716
rect 18463 13685 18475 13688
rect 18417 13679 18475 13685
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 23106 13676 23112 13728
rect 23164 13716 23170 13728
rect 23845 13719 23903 13725
rect 23845 13716 23857 13719
rect 23164 13688 23857 13716
rect 23164 13676 23170 13688
rect 23845 13685 23857 13688
rect 23891 13716 23903 13719
rect 25222 13716 25228 13728
rect 23891 13688 25228 13716
rect 23891 13685 23903 13688
rect 23845 13679 23903 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 25498 13716 25504 13728
rect 25459 13688 25504 13716
rect 25498 13676 25504 13688
rect 25556 13676 25562 13728
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 34238 13716 34244 13728
rect 31168 13688 34244 13716
rect 31168 13676 31174 13688
rect 34238 13676 34244 13688
rect 34296 13676 34302 13728
rect 34330 13676 34336 13728
rect 34388 13716 34394 13728
rect 35912 13716 35940 13756
rect 34388 13688 35940 13716
rect 36464 13716 36492 13756
rect 40221 13753 40233 13787
rect 40267 13753 40279 13787
rect 41046 13784 41052 13796
rect 40221 13747 40279 13753
rect 40328 13756 41052 13784
rect 40328 13716 40356 13756
rect 41046 13744 41052 13756
rect 41104 13744 41110 13796
rect 41322 13744 41328 13796
rect 41380 13784 41386 13796
rect 41708 13784 41736 13883
rect 41380 13756 41736 13784
rect 42260 13784 42288 13960
rect 43714 13948 43720 14000
rect 43772 13988 43778 14000
rect 43772 13960 44404 13988
rect 43772 13948 43778 13960
rect 43346 13920 43352 13932
rect 43307 13892 43352 13920
rect 43346 13880 43352 13892
rect 43404 13880 43410 13932
rect 43533 13923 43591 13929
rect 43533 13889 43545 13923
rect 43579 13920 43591 13923
rect 44082 13920 44088 13932
rect 43579 13892 44088 13920
rect 43579 13889 43591 13892
rect 43533 13883 43591 13889
rect 44082 13880 44088 13892
rect 44140 13880 44146 13932
rect 43806 13812 43812 13864
rect 43864 13852 43870 13864
rect 43990 13852 43996 13864
rect 43864 13824 43996 13852
rect 43864 13812 43870 13824
rect 43990 13812 43996 13824
rect 44048 13812 44054 13864
rect 44376 13861 44404 13960
rect 46842 13948 46848 14000
rect 46900 13988 46906 14000
rect 46900 13960 46945 13988
rect 46900 13948 46906 13960
rect 44531 13926 44589 13929
rect 44531 13923 44763 13926
rect 44531 13889 44543 13923
rect 44577 13920 44763 13923
rect 44818 13920 44824 13932
rect 44577 13898 44824 13920
rect 44577 13889 44589 13898
rect 44735 13892 44824 13898
rect 44531 13883 44589 13889
rect 44818 13880 44824 13892
rect 44876 13880 44882 13932
rect 46658 13920 46664 13932
rect 46619 13892 46664 13920
rect 46658 13880 46664 13892
rect 46716 13880 46722 13932
rect 46750 13880 46756 13932
rect 46808 13920 46814 13932
rect 46937 13923 46995 13929
rect 46937 13920 46949 13923
rect 46808 13892 46949 13920
rect 46808 13880 46814 13892
rect 46937 13889 46949 13892
rect 46983 13889 46995 13923
rect 46937 13883 46995 13889
rect 47029 13923 47087 13929
rect 47029 13889 47041 13923
rect 47075 13920 47087 13923
rect 47486 13920 47492 13932
rect 47075 13892 47492 13920
rect 47075 13889 47087 13892
rect 47029 13883 47087 13889
rect 47486 13880 47492 13892
rect 47544 13880 47550 13932
rect 47872 13920 47900 14028
rect 48130 14016 48136 14028
rect 48188 14016 48194 14068
rect 48222 14016 48228 14068
rect 48280 14056 48286 14068
rect 57238 14056 57244 14068
rect 48280 14028 57244 14056
rect 48280 14016 48286 14028
rect 57238 14016 57244 14028
rect 57296 14016 57302 14068
rect 47949 13923 48007 13929
rect 47949 13920 47961 13923
rect 47872 13892 47961 13920
rect 47949 13889 47961 13892
rect 47995 13889 48007 13923
rect 48866 13920 48872 13932
rect 47949 13883 48007 13889
rect 48056 13892 48872 13920
rect 44361 13855 44419 13861
rect 44361 13821 44373 13855
rect 44407 13852 44419 13855
rect 47765 13855 47823 13861
rect 47765 13852 47777 13855
rect 44407 13824 47777 13852
rect 44407 13821 44419 13824
rect 44361 13815 44419 13821
rect 47765 13821 47777 13824
rect 47811 13852 47823 13855
rect 48056 13852 48084 13892
rect 48866 13880 48872 13892
rect 48924 13880 48930 13932
rect 50798 13852 50804 13864
rect 47811 13824 48084 13852
rect 48286 13824 50804 13852
rect 47811 13821 47823 13824
rect 47765 13815 47823 13821
rect 48286 13784 48314 13824
rect 50798 13812 50804 13824
rect 50856 13812 50862 13864
rect 42260 13756 48314 13784
rect 41380 13744 41386 13756
rect 36464 13688 40356 13716
rect 34388 13676 34394 13688
rect 40402 13676 40408 13728
rect 40460 13716 40466 13728
rect 41340 13716 41368 13744
rect 40460 13688 41368 13716
rect 40460 13676 40466 13688
rect 41506 13676 41512 13728
rect 41564 13716 41570 13728
rect 49234 13716 49240 13728
rect 41564 13688 49240 13716
rect 41564 13676 41570 13688
rect 49234 13676 49240 13688
rect 49292 13676 49298 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11287 13484 16160 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 10597 13447 10655 13453
rect 10597 13413 10609 13447
rect 10643 13444 10655 13447
rect 12802 13444 12808 13456
rect 10643 13416 12808 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 12802 13404 12808 13416
rect 12860 13444 12866 13456
rect 16022 13444 16028 13456
rect 12860 13416 14780 13444
rect 15983 13416 16028 13444
rect 12860 13404 12866 13416
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 12253 13379 12311 13385
rect 12253 13376 12265 13379
rect 11664 13348 12265 13376
rect 11664 13336 11670 13348
rect 12253 13345 12265 13348
rect 12299 13345 12311 13379
rect 13538 13376 13544 13388
rect 13499 13348 13544 13376
rect 12253 13339 12311 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 13906 13376 13912 13388
rect 13679 13348 13912 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 14516 13348 14688 13376
rect 14516 13336 14522 13348
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13277 1639 13311
rect 10594 13308 10600 13320
rect 10555 13280 10600 13308
rect 1581 13271 1639 13277
rect 1596 13172 1624 13271
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11701 13311 11759 13317
rect 11480 13280 11525 13308
rect 11480 13268 11486 13280
rect 11701 13277 11713 13311
rect 11747 13308 11759 13311
rect 11882 13308 11888 13320
rect 11747 13280 11888 13308
rect 11747 13277 11759 13280
rect 11701 13271 11759 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 12360 13240 12388 13271
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12952 13280 13369 13308
rect 12952 13268 12958 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13286 13507 13311
rect 14090 13308 14096 13320
rect 13648 13286 14096 13308
rect 13495 13280 14096 13286
rect 13495 13277 13676 13280
rect 13449 13271 13676 13277
rect 13464 13258 13676 13271
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13305 14427 13311
rect 14550 13308 14556 13320
rect 14476 13305 14556 13308
rect 14415 13280 14556 13305
rect 14415 13277 14504 13280
rect 14369 13271 14427 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14660 13317 14688 13348
rect 14752 13317 14780 13416
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 16132 13444 16160 13484
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16264 13484 20484 13512
rect 16264 13472 16270 13484
rect 18966 13444 18972 13456
rect 16132 13416 18972 13444
rect 18966 13404 18972 13416
rect 19024 13404 19030 13456
rect 20456 13444 20484 13484
rect 21910 13472 21916 13524
rect 21968 13512 21974 13524
rect 25498 13512 25504 13524
rect 21968 13484 25504 13512
rect 21968 13472 21974 13484
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 28166 13472 28172 13524
rect 28224 13512 28230 13524
rect 31938 13512 31944 13524
rect 28224 13484 31944 13512
rect 28224 13472 28230 13484
rect 31938 13472 31944 13484
rect 31996 13472 32002 13524
rect 33226 13472 33232 13524
rect 33284 13512 33290 13524
rect 35434 13512 35440 13524
rect 33284 13484 35440 13512
rect 33284 13472 33290 13484
rect 35434 13472 35440 13484
rect 35492 13472 35498 13524
rect 35802 13472 35808 13524
rect 35860 13512 35866 13524
rect 37461 13515 37519 13521
rect 37461 13512 37473 13515
rect 35860 13484 37473 13512
rect 35860 13472 35866 13484
rect 37461 13481 37473 13484
rect 37507 13481 37519 13515
rect 37461 13475 37519 13481
rect 38105 13515 38163 13521
rect 38105 13481 38117 13515
rect 38151 13512 38163 13515
rect 38378 13512 38384 13524
rect 38151 13484 38384 13512
rect 38151 13481 38163 13484
rect 38105 13475 38163 13481
rect 38378 13472 38384 13484
rect 38436 13472 38442 13524
rect 41046 13472 41052 13524
rect 41104 13512 41110 13524
rect 45186 13512 45192 13524
rect 41104 13484 45192 13512
rect 41104 13472 41110 13484
rect 45186 13472 45192 13484
rect 45244 13472 45250 13524
rect 22925 13447 22983 13453
rect 22925 13444 22937 13447
rect 20456 13416 22937 13444
rect 22925 13413 22937 13416
rect 22971 13413 22983 13447
rect 22925 13407 22983 13413
rect 29733 13447 29791 13453
rect 29733 13413 29745 13447
rect 29779 13444 29791 13447
rect 32306 13444 32312 13456
rect 29779 13416 32312 13444
rect 29779 13413 29791 13416
rect 29733 13407 29791 13413
rect 32306 13404 32312 13416
rect 32364 13404 32370 13456
rect 32858 13404 32864 13456
rect 32916 13444 32922 13456
rect 34330 13444 34336 13456
rect 32916 13416 34336 13444
rect 32916 13404 32922 13416
rect 34330 13404 34336 13416
rect 34388 13404 34394 13456
rect 34790 13404 34796 13456
rect 34848 13444 34854 13456
rect 34848 13416 35204 13444
rect 34848 13404 34854 13416
rect 35176 13388 35204 13416
rect 36262 13404 36268 13456
rect 36320 13444 36326 13456
rect 36541 13447 36599 13453
rect 36541 13444 36553 13447
rect 36320 13416 36553 13444
rect 36320 13404 36326 13416
rect 36541 13413 36553 13416
rect 36587 13444 36599 13447
rect 37090 13444 37096 13456
rect 36587 13416 37096 13444
rect 36587 13413 36599 13416
rect 36541 13407 36599 13413
rect 37090 13404 37096 13416
rect 37148 13404 37154 13456
rect 37734 13404 37740 13456
rect 37792 13444 37798 13456
rect 40310 13444 40316 13456
rect 37792 13416 40316 13444
rect 37792 13404 37798 13416
rect 40310 13404 40316 13416
rect 40368 13404 40374 13456
rect 40402 13404 40408 13456
rect 40460 13404 40466 13456
rect 40678 13404 40684 13456
rect 40736 13444 40742 13456
rect 41414 13444 41420 13456
rect 40736 13416 41420 13444
rect 40736 13404 40742 13416
rect 41414 13404 41420 13416
rect 41472 13404 41478 13456
rect 41506 13404 41512 13456
rect 41564 13444 41570 13456
rect 43438 13444 43444 13456
rect 41564 13416 43444 13444
rect 41564 13404 41570 13416
rect 43438 13404 43444 13416
rect 43496 13404 43502 13456
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 19426 13376 19432 13388
rect 14976 13348 15700 13376
rect 14976 13336 14982 13348
rect 15672 13320 15700 13348
rect 15764 13348 19334 13376
rect 19387 13348 19432 13376
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15654 13308 15660 13320
rect 15615 13280 15660 13308
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 15764 13317 15792 13348
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15893 13311 15951 13317
rect 15893 13277 15905 13311
rect 15939 13308 15951 13311
rect 16206 13308 16212 13320
rect 15939 13280 16212 13308
rect 15939 13277 15951 13280
rect 15893 13271 15951 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 12360 13212 13400 13240
rect 2314 13172 2320 13184
rect 1596 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 11112 13144 11621 13172
rect 11112 13132 11118 13144
rect 11609 13141 11621 13144
rect 11655 13172 11667 13175
rect 12342 13172 12348 13184
rect 11655 13144 12348 13172
rect 11655 13141 11667 13144
rect 11609 13135 11667 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12713 13175 12771 13181
rect 12713 13141 12725 13175
rect 12759 13172 12771 13175
rect 12986 13172 12992 13184
rect 12759 13144 12992 13172
rect 12759 13141 12771 13144
rect 12713 13135 12771 13141
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 13170 13172 13176 13184
rect 13131 13144 13176 13172
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13372 13172 13400 13212
rect 13906 13172 13912 13184
rect 13372 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 14553 13175 14611 13181
rect 14553 13172 14565 13175
rect 14148 13144 14565 13172
rect 14148 13132 14154 13144
rect 14553 13141 14565 13144
rect 14599 13172 14611 13175
rect 14826 13172 14832 13184
rect 14599 13144 14832 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 14921 13175 14979 13181
rect 14921 13141 14933 13175
rect 14967 13172 14979 13175
rect 15028 13172 15056 13268
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 16592 13240 16620 13271
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 17494 13308 17500 13320
rect 16908 13280 17500 13308
rect 16908 13268 16914 13280
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18012 13280 18889 13308
rect 18012 13268 18018 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 19306 13308 19334 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 27617 13379 27675 13385
rect 27617 13376 27629 13379
rect 26108 13348 27629 13376
rect 26108 13336 26114 13348
rect 27617 13345 27629 13348
rect 27663 13345 27675 13379
rect 27617 13339 27675 13345
rect 27982 13336 27988 13388
rect 28040 13376 28046 13388
rect 29914 13376 29920 13388
rect 28040 13348 29920 13376
rect 28040 13336 28046 13348
rect 29914 13336 29920 13348
rect 29972 13376 29978 13388
rect 30285 13379 30343 13385
rect 30285 13376 30297 13379
rect 29972 13348 30297 13376
rect 29972 13336 29978 13348
rect 30285 13345 30297 13348
rect 30331 13345 30343 13379
rect 32674 13376 32680 13388
rect 30285 13339 30343 13345
rect 30944 13348 32680 13376
rect 21634 13308 21640 13320
rect 19306 13280 21640 13308
rect 18877 13271 18935 13277
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 21729 13311 21787 13317
rect 21729 13277 21741 13311
rect 21775 13308 21787 13311
rect 21910 13308 21916 13320
rect 21775 13280 21916 13308
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 21910 13268 21916 13280
rect 21968 13268 21974 13320
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 22520 13280 24593 13308
rect 22520 13268 22526 13280
rect 24581 13277 24593 13280
rect 24627 13308 24639 13311
rect 25130 13308 25136 13320
rect 24627 13280 25136 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 26510 13308 26516 13320
rect 26471 13280 26516 13308
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 30101 13311 30159 13317
rect 26752 13280 27844 13308
rect 26752 13268 26758 13280
rect 16080 13212 16620 13240
rect 16080 13200 16086 13212
rect 17402 13200 17408 13252
rect 17460 13240 17466 13252
rect 18046 13240 18052 13252
rect 17460 13212 18052 13240
rect 17460 13200 17466 13212
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 18782 13200 18788 13252
rect 18840 13240 18846 13252
rect 19674 13243 19732 13249
rect 19674 13240 19686 13243
rect 18840 13212 19686 13240
rect 18840 13200 18846 13212
rect 19674 13209 19686 13212
rect 19720 13209 19732 13243
rect 19674 13203 19732 13209
rect 20254 13200 20260 13252
rect 20312 13240 20318 13252
rect 20898 13240 20904 13252
rect 20312 13212 20904 13240
rect 20312 13200 20318 13212
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 24826 13243 24884 13249
rect 24826 13240 24838 13243
rect 22848 13212 24838 13240
rect 20806 13172 20812 13184
rect 14967 13144 15056 13172
rect 20767 13144 20812 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 21450 13132 21456 13184
rect 21508 13172 21514 13184
rect 22848 13172 22876 13212
rect 24826 13209 24838 13212
rect 24872 13209 24884 13243
rect 27816 13240 27844 13280
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30944 13308 30972 13348
rect 32674 13336 32680 13348
rect 32732 13336 32738 13388
rect 32768 13348 33824 13376
rect 30147 13280 30972 13308
rect 31205 13311 31263 13317
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 31205 13277 31217 13311
rect 31251 13308 31263 13311
rect 32768 13308 32796 13348
rect 33594 13308 33600 13320
rect 31251 13280 32796 13308
rect 33555 13280 33600 13308
rect 31251 13277 31263 13280
rect 31205 13271 31263 13277
rect 24826 13203 24884 13209
rect 25976 13212 27660 13240
rect 27816 13212 30328 13240
rect 21508 13144 22876 13172
rect 21508 13132 21514 13144
rect 24302 13132 24308 13184
rect 24360 13172 24366 13184
rect 25976 13181 26004 13212
rect 25961 13175 26019 13181
rect 25961 13172 25973 13175
rect 24360 13144 25973 13172
rect 24360 13132 24366 13144
rect 25961 13141 25973 13144
rect 26007 13141 26019 13175
rect 25961 13135 26019 13141
rect 26142 13132 26148 13184
rect 26200 13172 26206 13184
rect 27522 13172 27528 13184
rect 26200 13144 27528 13172
rect 26200 13132 26206 13144
rect 27522 13132 27528 13144
rect 27580 13132 27586 13184
rect 27632 13172 27660 13212
rect 28258 13172 28264 13184
rect 27632 13144 28264 13172
rect 28258 13132 28264 13144
rect 28316 13132 28322 13184
rect 30098 13132 30104 13184
rect 30156 13172 30162 13184
rect 30193 13175 30251 13181
rect 30193 13172 30205 13175
rect 30156 13144 30205 13172
rect 30156 13132 30162 13144
rect 30193 13141 30205 13144
rect 30239 13141 30251 13175
rect 30300 13172 30328 13212
rect 30374 13200 30380 13252
rect 30432 13240 30438 13252
rect 31220 13240 31248 13271
rect 33594 13268 33600 13280
rect 33652 13268 33658 13320
rect 33796 13308 33824 13348
rect 35158 13336 35164 13388
rect 35216 13376 35222 13388
rect 40126 13376 40132 13388
rect 35216 13348 35261 13376
rect 36179 13348 40132 13376
rect 35216 13336 35222 13348
rect 34992 13308 35112 13310
rect 36179 13308 36207 13348
rect 40126 13336 40132 13348
rect 40184 13336 40190 13388
rect 33796 13302 35112 13308
rect 35173 13302 36207 13308
rect 33796 13282 36207 13302
rect 33796 13280 35020 13282
rect 35084 13280 36207 13282
rect 37093 13311 37151 13317
rect 35084 13274 35201 13280
rect 37093 13277 37105 13311
rect 37139 13277 37151 13311
rect 37274 13308 37280 13320
rect 37235 13280 37280 13308
rect 37093 13271 37151 13277
rect 32950 13240 32956 13252
rect 30432 13212 31248 13240
rect 32911 13212 32956 13240
rect 30432 13200 30438 13212
rect 32950 13200 32956 13212
rect 33008 13200 33014 13252
rect 33410 13240 33416 13252
rect 33371 13212 33416 13240
rect 33410 13200 33416 13212
rect 33468 13200 33474 13252
rect 34974 13240 34980 13252
rect 33704 13212 34980 13240
rect 33704 13181 33732 13212
rect 34974 13200 34980 13212
rect 35032 13200 35038 13252
rect 35406 13243 35464 13249
rect 35406 13209 35418 13243
rect 35452 13240 35464 13243
rect 35526 13240 35532 13252
rect 35452 13212 35532 13240
rect 35452 13209 35464 13212
rect 35406 13203 35464 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 37108 13240 37136 13271
rect 37274 13268 37280 13280
rect 37332 13268 37338 13320
rect 37734 13268 37740 13320
rect 37792 13308 37798 13320
rect 37921 13311 37979 13317
rect 37921 13308 37933 13311
rect 37792 13280 37933 13308
rect 37792 13268 37798 13280
rect 37921 13277 37933 13280
rect 37967 13277 37979 13311
rect 37921 13271 37979 13277
rect 38378 13268 38384 13320
rect 38436 13308 38442 13320
rect 38749 13311 38807 13317
rect 38749 13308 38761 13311
rect 38436 13280 38761 13308
rect 38436 13268 38442 13280
rect 38749 13277 38761 13280
rect 38795 13277 38807 13311
rect 38749 13271 38807 13277
rect 39117 13311 39175 13317
rect 39117 13277 39129 13311
rect 39163 13277 39175 13311
rect 40034 13308 40040 13320
rect 39995 13280 40040 13308
rect 39117 13271 39175 13277
rect 35728 13212 37136 13240
rect 33689 13175 33747 13181
rect 33689 13172 33701 13175
rect 30300 13144 33701 13172
rect 30193 13135 30251 13141
rect 33689 13141 33701 13144
rect 33735 13141 33747 13175
rect 33689 13135 33747 13141
rect 34238 13132 34244 13184
rect 34296 13172 34302 13184
rect 35728 13172 35756 13212
rect 38654 13200 38660 13252
rect 38712 13240 38718 13252
rect 38838 13240 38844 13252
rect 38712 13212 38844 13240
rect 38712 13200 38718 13212
rect 38838 13200 38844 13212
rect 38896 13240 38902 13252
rect 39132 13240 39160 13271
rect 40034 13268 40040 13280
rect 40092 13268 40098 13320
rect 40420 13317 40448 13404
rect 43622 13336 43628 13388
rect 43680 13376 43686 13388
rect 57514 13376 57520 13388
rect 43680 13348 57520 13376
rect 43680 13336 43686 13348
rect 57514 13336 57520 13348
rect 57572 13336 57578 13388
rect 58158 13376 58164 13388
rect 58119 13348 58164 13376
rect 58158 13336 58164 13348
rect 58216 13336 58222 13388
rect 40313 13311 40371 13317
rect 40313 13308 40325 13311
rect 40144 13280 40325 13308
rect 38896 13212 39160 13240
rect 38896 13200 38902 13212
rect 39758 13200 39764 13252
rect 39816 13240 39822 13252
rect 40144 13240 40172 13280
rect 40313 13277 40325 13280
rect 40359 13277 40371 13311
rect 40313 13271 40371 13277
rect 40405 13311 40463 13317
rect 40405 13277 40417 13311
rect 40451 13277 40463 13311
rect 40770 13308 40776 13320
rect 40405 13271 40463 13277
rect 40538 13280 40776 13308
rect 39816 13212 40172 13240
rect 40221 13243 40279 13249
rect 39816 13200 39822 13212
rect 40221 13209 40233 13243
rect 40267 13240 40279 13243
rect 40538 13240 40566 13280
rect 40770 13268 40776 13280
rect 40828 13268 40834 13320
rect 41046 13308 41052 13320
rect 41007 13280 41052 13308
rect 41046 13268 41052 13280
rect 41104 13268 41110 13320
rect 41138 13268 41144 13320
rect 41196 13308 41202 13320
rect 41233 13311 41291 13317
rect 41233 13308 41245 13311
rect 41196 13280 41245 13308
rect 41196 13268 41202 13280
rect 41233 13277 41245 13280
rect 41279 13277 41291 13311
rect 41233 13271 41291 13277
rect 41325 13311 41383 13317
rect 41325 13277 41337 13311
rect 41371 13308 41383 13311
rect 41414 13308 41420 13320
rect 41371 13280 41420 13308
rect 41371 13277 41383 13280
rect 41325 13271 41383 13277
rect 41414 13268 41420 13280
rect 41472 13268 41478 13320
rect 41509 13311 41567 13317
rect 41509 13277 41521 13311
rect 41555 13277 41567 13311
rect 41509 13271 41567 13277
rect 41601 13311 41659 13317
rect 41601 13277 41613 13311
rect 41647 13308 41659 13311
rect 41966 13308 41972 13320
rect 41647 13280 41972 13308
rect 41647 13277 41659 13280
rect 41601 13271 41659 13277
rect 41524 13240 41552 13271
rect 41966 13268 41972 13280
rect 42024 13268 42030 13320
rect 42061 13311 42119 13317
rect 42061 13277 42073 13311
rect 42107 13277 42119 13311
rect 42061 13271 42119 13277
rect 40267 13212 40566 13240
rect 40604 13212 41552 13240
rect 40267 13209 40279 13212
rect 40221 13203 40279 13209
rect 34296 13144 35756 13172
rect 34296 13132 34302 13144
rect 35802 13132 35808 13184
rect 35860 13172 35866 13184
rect 39942 13172 39948 13184
rect 35860 13144 39948 13172
rect 35860 13132 35866 13144
rect 39942 13132 39948 13144
rect 40000 13132 40006 13184
rect 40604 13181 40632 13212
rect 40589 13175 40647 13181
rect 40589 13141 40601 13175
rect 40635 13141 40647 13175
rect 40589 13135 40647 13141
rect 41414 13132 41420 13184
rect 41472 13172 41478 13184
rect 42076 13172 42104 13271
rect 42150 13268 42156 13320
rect 42208 13308 42214 13320
rect 42208 13280 42253 13308
rect 42208 13268 42214 13280
rect 51074 13268 51080 13320
rect 51132 13308 51138 13320
rect 57885 13311 57943 13317
rect 57885 13308 57897 13311
rect 51132 13280 57897 13308
rect 51132 13268 51138 13280
rect 57885 13277 57897 13280
rect 57931 13277 57943 13311
rect 57885 13271 57943 13277
rect 57054 13240 57060 13252
rect 57015 13212 57060 13240
rect 57054 13200 57060 13212
rect 57112 13200 57118 13252
rect 41472 13144 42104 13172
rect 41472 13132 41478 13144
rect 48958 13132 48964 13184
rect 49016 13172 49022 13184
rect 57149 13175 57207 13181
rect 57149 13172 57161 13175
rect 49016 13144 57161 13172
rect 49016 13132 49022 13144
rect 57149 13141 57161 13144
rect 57195 13141 57207 13175
rect 57149 13135 57207 13141
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 12529 12971 12587 12977
rect 12529 12937 12541 12971
rect 12575 12968 12587 12971
rect 12618 12968 12624 12980
rect 12575 12940 12624 12968
rect 12575 12937 12587 12940
rect 12529 12931 12587 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 15654 12968 15660 12980
rect 13228 12940 15660 12968
rect 13228 12928 13234 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 17865 12971 17923 12977
rect 17865 12968 17877 12971
rect 15804 12940 17877 12968
rect 15804 12928 15810 12940
rect 17865 12937 17877 12940
rect 17911 12968 17923 12971
rect 17911 12940 17984 12968
rect 17911 12937 17923 12940
rect 17865 12931 17923 12937
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12900 10195 12903
rect 12710 12900 12716 12912
rect 10183 12872 12716 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 13538 12860 13544 12912
rect 13596 12900 13602 12912
rect 13596 12872 14044 12900
rect 13596 12860 13602 12872
rect 10042 12832 10048 12844
rect 10003 12804 10048 12832
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 11882 12832 11888 12844
rect 10275 12804 11888 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12492 12804 13185 12832
rect 12492 12792 12498 12804
rect 13173 12801 13185 12804
rect 13219 12832 13231 12835
rect 13722 12832 13728 12844
rect 13219 12804 13728 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14016 12841 14044 12872
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 17402 12900 17408 12912
rect 14792 12872 17408 12900
rect 14792 12860 14798 12872
rect 17402 12860 17408 12872
rect 17460 12900 17466 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 17460 12872 17785 12900
rect 17460 12860 17466 12872
rect 17773 12869 17785 12872
rect 17819 12869 17831 12903
rect 17956 12900 17984 12940
rect 18230 12928 18236 12980
rect 18288 12968 18294 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 18288 12940 25237 12968
rect 18288 12928 18294 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 25225 12931 25283 12937
rect 26970 12928 26976 12980
rect 27028 12968 27034 12980
rect 27338 12968 27344 12980
rect 27028 12940 27344 12968
rect 27028 12928 27034 12940
rect 27338 12928 27344 12940
rect 27396 12928 27402 12980
rect 27614 12968 27620 12980
rect 27448 12940 27620 12968
rect 17956 12872 19288 12900
rect 17773 12863 17831 12869
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16908 12804 16957 12832
rect 16908 12792 16914 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17310 12832 17316 12844
rect 17175 12804 17316 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17954 12841 17960 12844
rect 17941 12835 17960 12841
rect 17941 12801 17953 12835
rect 17941 12795 17960 12801
rect 17954 12792 17960 12795
rect 18012 12792 18018 12844
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 18288 12804 19165 12832
rect 18288 12792 18294 12804
rect 19153 12801 19165 12804
rect 19199 12801 19211 12835
rect 19260 12832 19288 12872
rect 20254 12860 20260 12912
rect 20312 12900 20318 12912
rect 22278 12909 22284 12912
rect 20312 12872 21680 12900
rect 20312 12860 20318 12872
rect 21652 12832 21680 12872
rect 22272 12863 22284 12909
rect 22336 12900 22342 12912
rect 22336 12872 22372 12900
rect 22278 12860 22284 12863
rect 22336 12860 22342 12872
rect 25038 12860 25044 12912
rect 25096 12900 25102 12912
rect 26050 12900 26056 12912
rect 25096 12872 26056 12900
rect 25096 12860 25102 12872
rect 26050 12860 26056 12872
rect 26108 12860 26114 12912
rect 26510 12860 26516 12912
rect 26568 12900 26574 12912
rect 27448 12909 27476 12940
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 27709 12971 27767 12977
rect 27709 12937 27721 12971
rect 27755 12968 27767 12971
rect 46658 12968 46664 12980
rect 27755 12940 41276 12968
rect 27755 12937 27767 12940
rect 27709 12931 27767 12937
rect 27433 12903 27491 12909
rect 27433 12900 27445 12903
rect 26568 12872 27445 12900
rect 26568 12860 26574 12872
rect 27433 12869 27445 12872
rect 27479 12869 27491 12903
rect 27798 12900 27804 12912
rect 27433 12863 27491 12869
rect 27586 12872 27804 12900
rect 19260 12804 20944 12832
rect 21652 12804 23060 12832
rect 19153 12795 19211 12801
rect 10686 12764 10692 12776
rect 10647 12736 10692 12764
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 13265 12767 13323 12773
rect 12115 12736 13216 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 10962 12696 10968 12708
rect 10923 12668 10968 12696
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 12342 12696 12348 12708
rect 12303 12668 12348 12696
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 13188 12696 13216 12736
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13538 12764 13544 12776
rect 13311 12736 13544 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14182 12764 14188 12776
rect 13648 12736 14188 12764
rect 13648 12696 13676 12736
rect 14182 12724 14188 12736
rect 14240 12764 14246 12776
rect 14550 12764 14556 12776
rect 14240 12736 14556 12764
rect 14240 12724 14246 12736
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 15102 12764 15108 12776
rect 15063 12736 15108 12764
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17589 12767 17647 12773
rect 17589 12764 17601 12767
rect 17236 12736 17601 12764
rect 13188 12668 13676 12696
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 15838 12696 15844 12708
rect 13780 12668 15844 12696
rect 13780 12656 13786 12668
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 13449 12631 13507 12637
rect 13449 12597 13461 12631
rect 13495 12628 13507 12631
rect 13814 12628 13820 12640
rect 13495 12600 13820 12628
rect 13495 12597 13507 12600
rect 13449 12591 13507 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14734 12628 14740 12640
rect 13964 12600 14740 12628
rect 13964 12588 13970 12600
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 17236 12628 17264 12736
rect 17589 12733 17601 12736
rect 17635 12764 17647 12767
rect 18325 12767 18383 12773
rect 17635 12736 17816 12764
rect 17635 12733 17647 12736
rect 17589 12727 17647 12733
rect 17788 12696 17816 12736
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18598 12764 18604 12776
rect 18371 12736 18604 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 20254 12764 20260 12776
rect 19168 12736 20260 12764
rect 19168 12696 19196 12736
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20346 12724 20352 12776
rect 20404 12764 20410 12776
rect 20806 12764 20812 12776
rect 20404 12736 20812 12764
rect 20404 12724 20410 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 20714 12696 20720 12708
rect 17788 12668 19196 12696
rect 19306 12668 20720 12696
rect 14884 12600 17264 12628
rect 14884 12588 14890 12600
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 19306 12628 19334 12668
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 20346 12628 20352 12640
rect 18104 12600 19334 12628
rect 20307 12600 20352 12628
rect 18104 12588 18110 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20916 12628 20944 12804
rect 22002 12764 22008 12776
rect 21963 12736 22008 12764
rect 22002 12724 22008 12736
rect 22060 12724 22066 12776
rect 23032 12764 23060 12804
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 24084 12804 24129 12832
rect 24084 12792 24090 12804
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 26476 12804 27169 12832
rect 26476 12792 26482 12804
rect 27157 12801 27169 12804
rect 27203 12832 27215 12835
rect 27203 12804 27292 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 24210 12764 24216 12776
rect 23032 12736 24216 12764
rect 24210 12724 24216 12736
rect 24268 12724 24274 12776
rect 27264 12764 27292 12804
rect 27338 12792 27344 12844
rect 27396 12832 27402 12844
rect 27586 12841 27614 12872
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 32490 12900 32496 12912
rect 28000 12872 32352 12900
rect 32451 12872 32496 12900
rect 27571 12835 27629 12841
rect 27396 12804 27441 12832
rect 27396 12792 27402 12804
rect 27571 12801 27583 12835
rect 27617 12801 27629 12835
rect 28000 12832 28028 12872
rect 28166 12832 28172 12844
rect 27571 12795 27629 12801
rect 27715 12804 28028 12832
rect 28127 12804 28172 12832
rect 27715 12764 27743 12804
rect 28166 12792 28172 12804
rect 28224 12792 28230 12844
rect 28258 12792 28264 12844
rect 28316 12832 28322 12844
rect 32324 12841 32352 12872
rect 32490 12860 32496 12872
rect 32548 12860 32554 12912
rect 32582 12860 32588 12912
rect 32640 12900 32646 12912
rect 36446 12900 36452 12912
rect 32640 12872 32685 12900
rect 36407 12872 36452 12900
rect 32640 12860 32646 12872
rect 36446 12860 36452 12872
rect 36504 12900 36510 12912
rect 37090 12900 37096 12912
rect 36504 12872 37096 12900
rect 36504 12860 36510 12872
rect 37090 12860 37096 12872
rect 37148 12860 37154 12912
rect 40954 12900 40960 12912
rect 40915 12872 40960 12900
rect 40954 12860 40960 12872
rect 41012 12860 41018 12912
rect 41248 12900 41276 12940
rect 41386 12940 46664 12968
rect 41386 12900 41414 12940
rect 46658 12928 46664 12940
rect 46716 12928 46722 12980
rect 41248 12872 41414 12900
rect 42981 12903 43039 12909
rect 42981 12869 42993 12903
rect 43027 12900 43039 12903
rect 51902 12900 51908 12912
rect 43027 12872 51908 12900
rect 43027 12869 43039 12872
rect 42981 12863 43039 12869
rect 51902 12860 51908 12872
rect 51960 12860 51966 12912
rect 31297 12835 31355 12841
rect 31297 12832 31309 12835
rect 28316 12804 31309 12832
rect 28316 12792 28322 12804
rect 31297 12801 31309 12804
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 32677 12835 32735 12841
rect 32677 12801 32689 12835
rect 32723 12801 32735 12835
rect 32677 12795 32735 12801
rect 31386 12764 31392 12776
rect 27264 12736 27743 12764
rect 31299 12736 31392 12764
rect 31386 12724 31392 12736
rect 31444 12724 31450 12776
rect 31478 12724 31484 12776
rect 31536 12764 31542 12776
rect 31536 12736 31581 12764
rect 31536 12724 31542 12736
rect 23474 12696 23480 12708
rect 22940 12668 23480 12696
rect 22940 12628 22968 12668
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 27338 12656 27344 12708
rect 27396 12696 27402 12708
rect 29365 12699 29423 12705
rect 29365 12696 29377 12699
rect 27396 12668 29377 12696
rect 27396 12656 27402 12668
rect 29365 12665 29377 12668
rect 29411 12665 29423 12699
rect 29365 12659 29423 12665
rect 29730 12656 29736 12708
rect 29788 12696 29794 12708
rect 30929 12699 30987 12705
rect 30929 12696 30941 12699
rect 29788 12668 30941 12696
rect 29788 12656 29794 12668
rect 30929 12665 30941 12668
rect 30975 12665 30987 12699
rect 30929 12659 30987 12665
rect 20916 12600 22968 12628
rect 23382 12588 23388 12640
rect 23440 12628 23446 12640
rect 23440 12600 23485 12628
rect 23440 12588 23446 12600
rect 27568 12588 27574 12640
rect 27626 12628 27632 12640
rect 31404 12628 31432 12724
rect 32692 12640 32720 12795
rect 32950 12792 32956 12844
rect 33008 12832 33014 12844
rect 33873 12835 33931 12841
rect 33873 12832 33885 12835
rect 33008 12804 33885 12832
rect 33008 12792 33014 12804
rect 33873 12801 33885 12804
rect 33919 12832 33931 12835
rect 34790 12832 34796 12844
rect 33919 12804 34796 12832
rect 33919 12801 33931 12804
rect 33873 12795 33931 12801
rect 34790 12792 34796 12804
rect 34848 12792 34854 12844
rect 35802 12832 35808 12844
rect 34900 12804 35808 12832
rect 34149 12767 34207 12773
rect 34149 12733 34161 12767
rect 34195 12764 34207 12767
rect 34900 12764 34928 12804
rect 35802 12792 35808 12804
rect 35860 12792 35866 12844
rect 36078 12832 36084 12844
rect 35991 12804 36084 12832
rect 36078 12792 36084 12804
rect 36136 12832 36142 12844
rect 36538 12832 36544 12844
rect 36136 12804 36544 12832
rect 36136 12792 36142 12804
rect 36538 12792 36544 12804
rect 36596 12792 36602 12844
rect 36814 12792 36820 12844
rect 36872 12832 36878 12844
rect 39666 12832 39672 12844
rect 36872 12804 38976 12832
rect 39627 12804 39672 12832
rect 36872 12792 36878 12804
rect 38948 12776 38976 12804
rect 39666 12792 39672 12804
rect 39724 12792 39730 12844
rect 39853 12835 39911 12841
rect 39853 12832 39865 12835
rect 39776 12804 39865 12832
rect 39776 12776 39804 12804
rect 39853 12801 39865 12804
rect 39899 12832 39911 12835
rect 39942 12832 39948 12844
rect 39899 12804 39948 12832
rect 39899 12801 39911 12804
rect 39853 12795 39911 12801
rect 39942 12792 39948 12804
rect 40000 12792 40006 12844
rect 40678 12832 40684 12844
rect 40639 12804 40684 12832
rect 40678 12792 40684 12804
rect 40736 12792 40742 12844
rect 40770 12792 40776 12844
rect 40828 12832 40834 12844
rect 40865 12835 40923 12841
rect 40865 12832 40877 12835
rect 40828 12804 40877 12832
rect 40828 12792 40834 12804
rect 40865 12801 40877 12804
rect 40911 12801 40923 12835
rect 40865 12795 40923 12801
rect 41049 12835 41107 12841
rect 41049 12801 41061 12835
rect 41095 12832 41107 12835
rect 41322 12832 41328 12844
rect 41095 12804 41328 12832
rect 41095 12801 41107 12804
rect 41049 12795 41107 12801
rect 41322 12792 41328 12804
rect 41380 12792 41386 12844
rect 41874 12832 41880 12844
rect 41835 12804 41880 12832
rect 41874 12792 41880 12804
rect 41932 12792 41938 12844
rect 34195 12736 34928 12764
rect 34195 12733 34207 12736
rect 34149 12727 34207 12733
rect 35158 12724 35164 12776
rect 35216 12764 35222 12776
rect 37366 12764 37372 12776
rect 35216 12736 37372 12764
rect 35216 12724 35222 12736
rect 37366 12724 37372 12736
rect 37424 12764 37430 12776
rect 37461 12767 37519 12773
rect 37461 12764 37473 12767
rect 37424 12736 37473 12764
rect 37424 12724 37430 12736
rect 37461 12733 37473 12736
rect 37507 12733 37519 12767
rect 37734 12764 37740 12776
rect 37695 12736 37740 12764
rect 37461 12727 37519 12733
rect 37734 12724 37740 12736
rect 37792 12724 37798 12776
rect 38930 12764 38936 12776
rect 38891 12736 38936 12764
rect 38930 12724 38936 12736
rect 38988 12724 38994 12776
rect 39758 12724 39764 12776
rect 39816 12724 39822 12776
rect 41414 12764 41420 12776
rect 39868 12736 41420 12764
rect 32858 12696 32864 12708
rect 32819 12668 32864 12696
rect 32858 12656 32864 12668
rect 32916 12656 32922 12708
rect 37274 12696 37280 12708
rect 34808 12668 37280 12696
rect 32674 12628 32680 12640
rect 27626 12600 31432 12628
rect 32587 12600 32680 12628
rect 27626 12588 27632 12600
rect 32674 12588 32680 12600
rect 32732 12628 32738 12640
rect 34808 12628 34836 12668
rect 37274 12656 37280 12668
rect 37332 12656 37338 12708
rect 39114 12696 39120 12708
rect 38764 12668 39120 12696
rect 35434 12628 35440 12640
rect 32732 12600 34836 12628
rect 35395 12600 35440 12628
rect 32732 12588 32738 12600
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 35802 12588 35808 12640
rect 35860 12628 35866 12640
rect 38764 12628 38792 12668
rect 39114 12656 39120 12668
rect 39172 12656 39178 12708
rect 39574 12656 39580 12708
rect 39632 12696 39638 12708
rect 39868 12696 39896 12736
rect 41414 12724 41420 12736
rect 41472 12724 41478 12776
rect 41693 12767 41751 12773
rect 41693 12733 41705 12767
rect 41739 12764 41751 12767
rect 42058 12764 42064 12776
rect 41739 12736 42064 12764
rect 41739 12733 41751 12736
rect 41693 12727 41751 12733
rect 42058 12724 42064 12736
rect 42116 12724 42122 12776
rect 43070 12764 43076 12776
rect 43031 12736 43076 12764
rect 43070 12724 43076 12736
rect 43128 12724 43134 12776
rect 43162 12724 43168 12776
rect 43220 12764 43226 12776
rect 43346 12764 43352 12776
rect 43220 12736 43352 12764
rect 43220 12724 43226 12736
rect 43346 12724 43352 12736
rect 43404 12724 43410 12776
rect 41233 12699 41291 12705
rect 41233 12696 41245 12699
rect 39632 12668 39896 12696
rect 41156 12668 41245 12696
rect 39632 12656 39638 12668
rect 39942 12628 39948 12640
rect 35860 12600 38792 12628
rect 39903 12600 39948 12628
rect 35860 12588 35866 12600
rect 39942 12588 39948 12600
rect 40000 12588 40006 12640
rect 40494 12588 40500 12640
rect 40552 12628 40558 12640
rect 41156 12628 41184 12668
rect 41233 12665 41245 12668
rect 41279 12665 41291 12699
rect 41233 12659 41291 12665
rect 41506 12656 41512 12708
rect 41564 12696 41570 12708
rect 50062 12696 50068 12708
rect 41564 12668 50068 12696
rect 41564 12656 41570 12668
rect 50062 12656 50068 12668
rect 50120 12656 50126 12708
rect 40552 12600 41184 12628
rect 40552 12588 40558 12600
rect 41782 12588 41788 12640
rect 41840 12628 41846 12640
rect 42061 12631 42119 12637
rect 42061 12628 42073 12631
rect 41840 12600 42073 12628
rect 41840 12588 41846 12600
rect 42061 12597 42073 12600
rect 42107 12597 42119 12631
rect 42061 12591 42119 12597
rect 42613 12631 42671 12637
rect 42613 12597 42625 12631
rect 42659 12628 42671 12631
rect 42886 12628 42892 12640
rect 42659 12600 42892 12628
rect 42659 12597 42671 12600
rect 42613 12591 42671 12597
rect 42886 12588 42892 12600
rect 42944 12588 42950 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 10100 12396 12633 12424
rect 10100 12384 10106 12396
rect 12621 12393 12633 12396
rect 12667 12424 12679 12427
rect 12894 12424 12900 12436
rect 12667 12396 12900 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14056 12396 14381 12424
rect 14056 12384 14062 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 14608 12396 16037 12424
rect 14608 12384 14614 12396
rect 16025 12393 16037 12396
rect 16071 12424 16083 12427
rect 17954 12424 17960 12436
rect 16071 12396 17960 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19444 12396 20668 12424
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 10744 12328 11836 12356
rect 10744 12316 10750 12328
rect 11808 12300 11836 12328
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 19444 12356 19472 12396
rect 12032 12328 14136 12356
rect 12032 12316 12038 12328
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 1596 12260 11437 12288
rect 1596 12229 1624 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11698 12288 11704 12300
rect 11659 12260 11704 12288
rect 11425 12251 11483 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 11848 12260 11941 12288
rect 11848 12248 11854 12260
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12189 1639 12223
rect 1854 12220 1860 12232
rect 1815 12192 1860 12220
rect 1581 12183 1639 12189
rect 1854 12180 1860 12192
rect 1912 12180 1918 12232
rect 11606 12220 11612 12232
rect 11567 12192 11612 12220
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 13265 12223 13323 12229
rect 11940 12192 11985 12220
rect 11940 12180 11946 12192
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13446 12220 13452 12232
rect 13311 12192 13452 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 12434 12152 12440 12164
rect 12395 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 12618 12112 12624 12164
rect 12676 12161 12682 12164
rect 12676 12155 12695 12161
rect 12683 12121 12695 12155
rect 12676 12115 12695 12121
rect 12676 12112 12682 12115
rect 12986 12112 12992 12164
rect 13044 12152 13050 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13044 12124 13553 12152
rect 13044 12112 13050 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 14108 12152 14136 12328
rect 15396 12328 19472 12356
rect 15396 12300 15424 12328
rect 14550 12288 14556 12300
rect 14511 12260 14556 12288
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 14734 12288 14740 12300
rect 14695 12260 14740 12288
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 15378 12288 15384 12300
rect 14884 12260 14929 12288
rect 15291 12260 15384 12288
rect 14884 12248 14890 12260
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 15930 12288 15936 12300
rect 15887 12260 15936 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 16298 12248 16304 12300
rect 16356 12288 16362 12300
rect 17218 12288 17224 12300
rect 16356 12260 17224 12288
rect 16356 12248 16362 12260
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 20640 12288 20668 12396
rect 21266 12384 21272 12436
rect 21324 12424 21330 12436
rect 24578 12424 24584 12436
rect 21324 12396 24584 12424
rect 21324 12384 21330 12396
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 32214 12424 32220 12436
rect 27586 12396 32220 12424
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 22925 12359 22983 12365
rect 22925 12356 22937 12359
rect 20772 12328 22937 12356
rect 20772 12316 20778 12328
rect 22925 12325 22937 12328
rect 22971 12325 22983 12359
rect 27586 12356 27614 12396
rect 32214 12384 32220 12396
rect 32272 12384 32278 12436
rect 33137 12427 33195 12433
rect 33137 12393 33149 12427
rect 33183 12424 33195 12427
rect 33226 12424 33232 12436
rect 33183 12396 33232 12424
rect 33183 12393 33195 12396
rect 33137 12387 33195 12393
rect 33226 12384 33232 12396
rect 33284 12384 33290 12436
rect 34054 12384 34060 12436
rect 34112 12424 34118 12436
rect 36078 12424 36084 12436
rect 34112 12396 36084 12424
rect 34112 12384 34118 12396
rect 36078 12384 36084 12396
rect 36136 12384 36142 12436
rect 36538 12384 36544 12436
rect 36596 12424 36602 12436
rect 39114 12424 39120 12436
rect 36596 12396 38654 12424
rect 39075 12396 39120 12424
rect 36596 12384 36602 12396
rect 22925 12319 22983 12325
rect 23032 12328 27614 12356
rect 23032 12288 23060 12328
rect 28718 12316 28724 12368
rect 28776 12356 28782 12368
rect 32232 12356 32260 12384
rect 28776 12328 30972 12356
rect 32232 12328 34468 12356
rect 28776 12316 28782 12328
rect 20640 12260 23060 12288
rect 23474 12248 23480 12300
rect 23532 12288 23538 12300
rect 25685 12291 25743 12297
rect 25685 12288 25697 12291
rect 23532 12260 25697 12288
rect 23532 12248 23538 12260
rect 25685 12257 25697 12260
rect 25731 12257 25743 12291
rect 25685 12251 25743 12257
rect 29362 12248 29368 12300
rect 29420 12288 29426 12300
rect 30285 12291 30343 12297
rect 30285 12288 30297 12291
rect 29420 12260 30297 12288
rect 29420 12248 29426 12260
rect 30285 12257 30297 12260
rect 30331 12257 30343 12291
rect 30944 12288 30972 12328
rect 31570 12288 31576 12300
rect 30944 12260 31576 12288
rect 30285 12251 30343 12257
rect 31570 12248 31576 12260
rect 31628 12248 31634 12300
rect 31662 12248 31668 12300
rect 31720 12288 31726 12300
rect 33689 12291 33747 12297
rect 33689 12288 33701 12291
rect 31720 12260 33701 12288
rect 31720 12248 31726 12260
rect 33689 12257 33701 12260
rect 33735 12257 33747 12291
rect 33689 12251 33747 12257
rect 33778 12248 33784 12300
rect 33836 12288 33842 12300
rect 34054 12288 34060 12300
rect 33836 12260 34060 12288
rect 33836 12248 33842 12260
rect 34054 12248 34060 12260
rect 34112 12248 34118 12300
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15010 12220 15016 12232
rect 14691 12192 15016 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15160 12192 16344 12220
rect 15160 12180 15166 12192
rect 16316 12164 16344 12192
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16540 12192 16589 12220
rect 16540 12180 16546 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 19242 12220 19248 12232
rect 16908 12192 19248 12220
rect 16908 12180 16914 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 21729 12223 21787 12229
rect 19484 12192 20760 12220
rect 19484 12180 19490 12192
rect 15194 12152 15200 12164
rect 14108 12124 15200 12152
rect 13541 12115 13599 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 15657 12155 15715 12161
rect 15657 12152 15669 12155
rect 15528 12124 15669 12152
rect 15528 12112 15534 12124
rect 15657 12121 15669 12124
rect 15703 12152 15715 12155
rect 15703 12124 16252 12152
rect 15703 12121 15715 12124
rect 15657 12115 15715 12121
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 13814 12084 13820 12096
rect 12851 12056 13820 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 15838 12084 15844 12096
rect 15795 12056 15844 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 15838 12044 15844 12056
rect 15896 12084 15902 12096
rect 16114 12084 16120 12096
rect 15896 12056 16120 12084
rect 15896 12044 15902 12056
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16224 12084 16252 12124
rect 16298 12112 16304 12164
rect 16356 12112 16362 12164
rect 19696 12155 19754 12161
rect 19696 12121 19708 12155
rect 19742 12152 19754 12155
rect 20254 12152 20260 12164
rect 19742 12124 20260 12152
rect 19742 12121 19754 12124
rect 19696 12115 19754 12121
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 20732 12152 20760 12192
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 24578 12220 24584 12232
rect 21775 12192 24440 12220
rect 24539 12192 24584 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22002 12152 22008 12164
rect 20732 12124 22008 12152
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 24412 12152 24440 12192
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 25130 12180 25136 12232
rect 25188 12220 25194 12232
rect 27709 12223 27767 12229
rect 27709 12220 27721 12223
rect 25188 12192 27721 12220
rect 25188 12180 25194 12192
rect 27709 12189 27721 12192
rect 27755 12220 27767 12223
rect 29822 12220 29828 12232
rect 27755 12192 29828 12220
rect 27755 12189 27767 12192
rect 27709 12183 27767 12189
rect 29822 12180 29828 12192
rect 29880 12180 29886 12232
rect 30929 12223 30987 12229
rect 30929 12189 30941 12223
rect 30975 12220 30987 12223
rect 31018 12220 31024 12232
rect 30975 12192 31024 12220
rect 30975 12189 30987 12192
rect 30929 12183 30987 12189
rect 31018 12180 31024 12192
rect 31076 12180 31082 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 33410 12220 33416 12232
rect 31251 12192 33416 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 33410 12180 33416 12192
rect 33468 12180 33474 12232
rect 33505 12223 33563 12229
rect 33505 12189 33517 12223
rect 33551 12220 33563 12223
rect 33870 12220 33876 12232
rect 33551 12192 33876 12220
rect 33551 12189 33563 12192
rect 33505 12183 33563 12189
rect 33870 12180 33876 12192
rect 33928 12220 33934 12232
rect 34238 12220 34244 12232
rect 33928 12192 34244 12220
rect 33928 12180 33934 12192
rect 34238 12180 34244 12192
rect 34296 12180 34302 12232
rect 27338 12152 27344 12164
rect 24412 12124 27344 12152
rect 27338 12112 27344 12124
rect 27396 12112 27402 12164
rect 27976 12155 28034 12161
rect 27976 12121 27988 12155
rect 28022 12152 28034 12155
rect 29914 12152 29920 12164
rect 28022 12124 29920 12152
rect 28022 12121 28034 12124
rect 27976 12115 28034 12121
rect 29914 12112 29920 12124
rect 29972 12112 29978 12164
rect 30006 12112 30012 12164
rect 30064 12152 30070 12164
rect 30101 12155 30159 12161
rect 30101 12152 30113 12155
rect 30064 12124 30113 12152
rect 30064 12112 30070 12124
rect 30101 12121 30113 12124
rect 30147 12121 30159 12155
rect 30101 12115 30159 12121
rect 31864 12124 32904 12152
rect 20438 12084 20444 12096
rect 16224 12056 20444 12084
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12084 20867 12087
rect 23106 12084 23112 12096
rect 20855 12056 23112 12084
rect 20855 12053 20867 12056
rect 20809 12047 20867 12053
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 29089 12087 29147 12093
rect 29089 12084 29101 12087
rect 27764 12056 29101 12084
rect 27764 12044 27770 12056
rect 29089 12053 29101 12056
rect 29135 12053 29147 12087
rect 29089 12047 29147 12053
rect 29178 12044 29184 12096
rect 29236 12084 29242 12096
rect 29733 12087 29791 12093
rect 29733 12084 29745 12087
rect 29236 12056 29745 12084
rect 29236 12044 29242 12056
rect 29733 12053 29745 12056
rect 29779 12053 29791 12087
rect 30190 12084 30196 12096
rect 30151 12056 30196 12084
rect 29733 12047 29791 12053
rect 30190 12044 30196 12056
rect 30248 12044 30254 12096
rect 31478 12044 31484 12096
rect 31536 12084 31542 12096
rect 31864 12084 31892 12124
rect 31536 12056 31892 12084
rect 31536 12044 31542 12056
rect 31938 12044 31944 12096
rect 31996 12084 32002 12096
rect 32490 12084 32496 12096
rect 31996 12056 32496 12084
rect 31996 12044 32002 12056
rect 32490 12044 32496 12056
rect 32548 12044 32554 12096
rect 32876 12084 32904 12124
rect 32950 12112 32956 12164
rect 33008 12152 33014 12164
rect 33597 12155 33655 12161
rect 33597 12152 33609 12155
rect 33008 12124 33609 12152
rect 33008 12112 33014 12124
rect 33597 12121 33609 12124
rect 33643 12121 33655 12155
rect 34440 12152 34468 12328
rect 35158 12316 35164 12368
rect 35216 12356 35222 12368
rect 35434 12356 35440 12368
rect 35216 12328 35440 12356
rect 35216 12316 35222 12328
rect 35434 12316 35440 12328
rect 35492 12316 35498 12368
rect 35526 12316 35532 12368
rect 35584 12356 35590 12368
rect 36262 12356 36268 12368
rect 35584 12328 36268 12356
rect 35584 12316 35590 12328
rect 36262 12316 36268 12328
rect 36320 12316 36326 12368
rect 37274 12316 37280 12368
rect 37332 12356 37338 12368
rect 37553 12359 37611 12365
rect 37553 12356 37565 12359
rect 37332 12328 37565 12356
rect 37332 12316 37338 12328
rect 37553 12325 37565 12328
rect 37599 12325 37611 12359
rect 37553 12319 37611 12325
rect 37642 12316 37648 12368
rect 37700 12356 37706 12368
rect 37700 12328 38139 12356
rect 37700 12316 37706 12328
rect 34514 12248 34520 12300
rect 34572 12288 34578 12300
rect 34572 12260 35572 12288
rect 34572 12248 34578 12260
rect 35222 12223 35280 12229
rect 35222 12189 35234 12223
rect 35268 12220 35280 12223
rect 35434 12220 35440 12232
rect 35268 12192 35440 12220
rect 35268 12189 35280 12192
rect 35222 12183 35280 12189
rect 35434 12180 35440 12192
rect 35492 12180 35498 12232
rect 35544 12152 35572 12260
rect 35618 12248 35624 12300
rect 35676 12288 35682 12300
rect 35676 12260 35721 12288
rect 35676 12248 35682 12260
rect 36078 12248 36084 12300
rect 36136 12288 36142 12300
rect 36173 12291 36231 12297
rect 36173 12288 36185 12291
rect 36136 12260 36185 12288
rect 36136 12248 36142 12260
rect 36173 12257 36185 12260
rect 36219 12257 36231 12291
rect 36541 12291 36599 12297
rect 36541 12288 36553 12291
rect 36173 12251 36231 12257
rect 36280 12260 36553 12288
rect 35710 12220 35716 12232
rect 35671 12192 35716 12220
rect 35710 12180 35716 12192
rect 35768 12180 35774 12232
rect 35802 12180 35808 12232
rect 35860 12220 35866 12232
rect 36280 12220 36308 12260
rect 36541 12257 36553 12260
rect 36587 12257 36599 12291
rect 38010 12288 38016 12300
rect 37971 12260 38016 12288
rect 36541 12251 36599 12257
rect 38010 12248 38016 12260
rect 38068 12248 38074 12300
rect 38111 12232 38139 12328
rect 38197 12291 38255 12297
rect 38197 12257 38209 12291
rect 38243 12257 38255 12291
rect 38626 12288 38654 12396
rect 39114 12384 39120 12396
rect 39172 12384 39178 12436
rect 41414 12384 41420 12436
rect 41472 12424 41478 12436
rect 43073 12427 43131 12433
rect 43073 12424 43085 12427
rect 41472 12396 43085 12424
rect 41472 12384 41478 12396
rect 43073 12393 43085 12396
rect 43119 12424 43131 12427
rect 43622 12424 43628 12436
rect 43119 12396 43628 12424
rect 43119 12393 43131 12396
rect 43073 12387 43131 12393
rect 43622 12384 43628 12396
rect 43680 12384 43686 12436
rect 41509 12291 41567 12297
rect 38626 12260 41414 12288
rect 38197 12251 38255 12257
rect 35860 12192 36308 12220
rect 36357 12223 36415 12229
rect 35860 12180 35866 12192
rect 36357 12189 36369 12223
rect 36403 12220 36415 12223
rect 36446 12220 36452 12232
rect 36403 12192 36452 12220
rect 36403 12189 36415 12192
rect 36357 12183 36415 12189
rect 36446 12180 36452 12192
rect 36504 12180 36510 12232
rect 37918 12220 37924 12232
rect 37879 12192 37924 12220
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 38102 12180 38108 12232
rect 38160 12220 38166 12232
rect 38212 12220 38240 12251
rect 38838 12220 38844 12232
rect 38160 12192 38253 12220
rect 38799 12192 38844 12220
rect 38160 12180 38166 12192
rect 38838 12180 38844 12192
rect 38896 12180 38902 12232
rect 38933 12223 38991 12229
rect 38933 12189 38945 12223
rect 38979 12189 38991 12223
rect 38933 12183 38991 12189
rect 38948 12152 38976 12183
rect 39758 12180 39764 12232
rect 39816 12220 39822 12232
rect 40221 12223 40279 12229
rect 40221 12220 40233 12223
rect 39816 12192 40233 12220
rect 39816 12180 39822 12192
rect 40221 12189 40233 12192
rect 40267 12189 40279 12223
rect 40221 12183 40279 12189
rect 34440 12124 35379 12152
rect 35544 12124 38976 12152
rect 40037 12155 40095 12161
rect 33597 12115 33655 12121
rect 34882 12084 34888 12096
rect 32876 12056 34888 12084
rect 34882 12044 34888 12056
rect 34940 12044 34946 12096
rect 35066 12084 35072 12096
rect 35027 12056 35072 12084
rect 35066 12044 35072 12056
rect 35124 12044 35130 12096
rect 35250 12084 35256 12096
rect 35211 12056 35256 12084
rect 35250 12044 35256 12056
rect 35308 12044 35314 12096
rect 35351 12084 35379 12124
rect 40037 12121 40049 12155
rect 40083 12152 40095 12155
rect 41046 12152 41052 12164
rect 40083 12124 41052 12152
rect 40083 12121 40095 12124
rect 40037 12115 40095 12121
rect 41046 12112 41052 12124
rect 41104 12112 41110 12164
rect 39574 12084 39580 12096
rect 35351 12056 39580 12084
rect 39574 12044 39580 12056
rect 39632 12044 39638 12096
rect 40126 12044 40132 12096
rect 40184 12084 40190 12096
rect 40313 12087 40371 12093
rect 40313 12084 40325 12087
rect 40184 12056 40325 12084
rect 40184 12044 40190 12056
rect 40313 12053 40325 12056
rect 40359 12084 40371 12087
rect 40862 12084 40868 12096
rect 40359 12056 40868 12084
rect 40359 12053 40371 12056
rect 40313 12047 40371 12053
rect 40862 12044 40868 12056
rect 40920 12044 40926 12096
rect 41386 12084 41414 12260
rect 41509 12257 41521 12291
rect 41555 12288 41567 12291
rect 42702 12288 42708 12300
rect 41555 12260 42708 12288
rect 41555 12257 41567 12260
rect 41509 12251 41567 12257
rect 42702 12248 42708 12260
rect 42760 12248 42766 12300
rect 41782 12220 41788 12232
rect 41743 12192 41788 12220
rect 41782 12180 41788 12192
rect 41840 12180 41846 12232
rect 57514 12180 57520 12232
rect 57572 12220 57578 12232
rect 57885 12223 57943 12229
rect 57885 12220 57897 12223
rect 57572 12192 57897 12220
rect 57572 12180 57578 12192
rect 57885 12189 57897 12192
rect 57931 12189 57943 12223
rect 57885 12183 57943 12189
rect 46198 12152 46204 12164
rect 42444 12124 46204 12152
rect 42444 12084 42472 12124
rect 46198 12112 46204 12124
rect 46256 12112 46262 12164
rect 58158 12152 58164 12164
rect 58119 12124 58164 12152
rect 58158 12112 58164 12124
rect 58216 12112 58222 12164
rect 41386 12056 42472 12084
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7616 11852 12112 11880
rect 7616 11840 7622 11852
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 12084 11812 12112 11852
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 15286 11880 15292 11892
rect 12308 11852 14964 11880
rect 15247 11852 15292 11880
rect 12308 11840 12314 11852
rect 14734 11812 14740 11824
rect 11756 11784 11928 11812
rect 12084 11784 14740 11812
rect 11756 11772 11762 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 1627 11716 2774 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 1762 11676 1768 11688
rect 1723 11648 1768 11676
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 2746 11676 2774 11716
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11900 11744 11928 11784
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11664 11716 11836 11744
rect 11900 11716 11989 11744
rect 11664 11704 11670 11716
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 2746 11648 11713 11676
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11808 11676 11836 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 12894 11744 12900 11756
rect 12855 11716 12900 11744
rect 11977 11707 12035 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13814 11744 13820 11756
rect 13775 11716 13820 11744
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14936 11753 14964 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 17034 11880 17040 11892
rect 16995 11852 17040 11880
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 17218 11840 17224 11892
rect 17276 11880 17282 11892
rect 17276 11852 19840 11880
rect 17276 11840 17282 11852
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 15749 11815 15807 11821
rect 15068 11784 15700 11812
rect 15068 11772 15074 11784
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15470 11744 15476 11756
rect 14967 11716 15476 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11808 11648 11897 11676
rect 11701 11639 11759 11645
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 12084 11608 12112 11639
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12989 11679 13047 11685
rect 12216 11648 12261 11676
rect 12216 11636 12222 11648
rect 12989 11645 13001 11679
rect 13035 11676 13047 11679
rect 13906 11676 13912 11688
rect 13035 11648 13912 11676
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15378 11676 15384 11688
rect 15059 11648 15384 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 14182 11608 14188 11620
rect 11848 11580 12112 11608
rect 14143 11580 14188 11608
rect 11848 11568 11854 11580
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14277 11611 14335 11617
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 15562 11608 15568 11620
rect 14323 11580 15568 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 15672 11608 15700 11784
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 18046 11812 18052 11824
rect 15795 11784 18052 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 18046 11772 18052 11784
rect 18104 11772 18110 11824
rect 19334 11812 19340 11824
rect 18156 11784 19340 11812
rect 15930 11744 15936 11756
rect 15891 11716 15936 11744
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16298 11744 16304 11756
rect 16259 11716 16304 11744
rect 16025 11707 16083 11713
rect 16040 11676 16068 11707
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 16942 11744 16948 11756
rect 17000 11753 17006 11756
rect 17000 11747 17036 11753
rect 16632 11716 16948 11744
rect 16632 11704 16638 11716
rect 16942 11704 16948 11716
rect 17024 11713 17036 11747
rect 17000 11707 17036 11713
rect 17000 11704 17006 11707
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 17957 11747 18015 11753
rect 17460 11716 17908 11744
rect 17460 11704 17466 11716
rect 17310 11676 17316 11688
rect 16040 11648 17316 11676
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 17494 11676 17500 11688
rect 17455 11648 17500 11676
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 17880 11676 17908 11716
rect 17957 11713 17969 11747
rect 18003 11744 18015 11747
rect 18156 11744 18184 11784
rect 19334 11772 19340 11784
rect 19392 11772 19398 11824
rect 19812 11812 19840 11852
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 20312 11852 20361 11880
rect 20312 11840 20318 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 23106 11880 23112 11892
rect 20496 11852 23112 11880
rect 20496 11840 20502 11852
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 23385 11883 23443 11889
rect 23385 11849 23397 11883
rect 23431 11880 23443 11883
rect 24026 11880 24032 11892
rect 23431 11852 24032 11880
rect 23431 11849 23443 11852
rect 23385 11843 23443 11849
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 24268 11852 25513 11880
rect 24268 11840 24274 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 27430 11880 27436 11892
rect 26568 11852 27436 11880
rect 26568 11840 26574 11852
rect 27430 11840 27436 11852
rect 27488 11840 27494 11892
rect 27706 11840 27712 11892
rect 27764 11880 27770 11892
rect 27801 11883 27859 11889
rect 27801 11880 27813 11883
rect 27764 11852 27813 11880
rect 27764 11840 27770 11852
rect 27801 11849 27813 11852
rect 27847 11849 27859 11883
rect 29178 11880 29184 11892
rect 27801 11843 27859 11849
rect 27908 11852 29184 11880
rect 21266 11812 21272 11824
rect 19812 11784 21272 11812
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 26142 11812 26148 11824
rect 21876 11784 22968 11812
rect 21876 11772 21882 11784
rect 18003 11716 18184 11744
rect 18233 11747 18291 11753
rect 18003 11713 18015 11716
rect 17957 11707 18015 11713
rect 18233 11713 18245 11747
rect 18279 11744 18291 11747
rect 18782 11744 18788 11756
rect 18279 11716 18788 11744
rect 18279 11713 18291 11716
rect 18233 11707 18291 11713
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 19150 11744 19156 11756
rect 19111 11716 19156 11744
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 21358 11744 21364 11756
rect 19300 11716 21364 11744
rect 19300 11704 19306 11716
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 22002 11744 22008 11756
rect 21963 11716 22008 11744
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22278 11753 22284 11756
rect 22261 11747 22284 11753
rect 22261 11713 22273 11747
rect 22261 11707 22284 11713
rect 22278 11704 22284 11707
rect 22336 11704 22342 11756
rect 22940 11744 22968 11784
rect 24136 11784 26148 11812
rect 24136 11744 24164 11784
rect 26142 11772 26148 11784
rect 26200 11772 26206 11824
rect 27338 11772 27344 11824
rect 27396 11812 27402 11824
rect 27908 11812 27936 11852
rect 29178 11840 29184 11852
rect 29236 11840 29242 11892
rect 30006 11840 30012 11892
rect 30064 11880 30070 11892
rect 30926 11880 30932 11892
rect 30064 11852 30932 11880
rect 30064 11840 30070 11852
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 31294 11840 31300 11892
rect 31352 11880 31358 11892
rect 33318 11880 33324 11892
rect 31352 11852 33324 11880
rect 31352 11840 31358 11852
rect 33318 11840 33324 11852
rect 33376 11840 33382 11892
rect 33410 11840 33416 11892
rect 33468 11880 33474 11892
rect 33597 11883 33655 11889
rect 33597 11880 33609 11883
rect 33468 11852 33609 11880
rect 33468 11840 33474 11852
rect 33597 11849 33609 11852
rect 33643 11849 33655 11883
rect 33597 11843 33655 11849
rect 34057 11883 34115 11889
rect 34057 11849 34069 11883
rect 34103 11880 34115 11883
rect 34514 11880 34520 11892
rect 34103 11852 34520 11880
rect 34103 11849 34115 11852
rect 34057 11843 34115 11849
rect 34514 11840 34520 11852
rect 34572 11840 34578 11892
rect 35066 11840 35072 11892
rect 35124 11880 35130 11892
rect 35124 11852 39344 11880
rect 35124 11840 35130 11852
rect 27396 11784 27936 11812
rect 28629 11815 28687 11821
rect 27396 11772 27402 11784
rect 28629 11781 28641 11815
rect 28675 11812 28687 11815
rect 30374 11812 30380 11824
rect 28675 11784 30380 11812
rect 28675 11781 28687 11784
rect 28629 11775 28687 11781
rect 30374 11772 30380 11784
rect 30432 11772 30438 11824
rect 32398 11812 32404 11824
rect 30484 11784 31340 11812
rect 32359 11784 32404 11812
rect 24302 11744 24308 11756
rect 22940 11716 24164 11744
rect 24263 11716 24308 11744
rect 24302 11704 24308 11716
rect 24360 11704 24366 11756
rect 24486 11704 24492 11756
rect 24544 11744 24550 11756
rect 30484 11744 30512 11784
rect 24544 11716 30512 11744
rect 24544 11704 24550 11716
rect 30558 11704 30564 11756
rect 30616 11744 30622 11756
rect 31205 11747 31263 11753
rect 31205 11744 31217 11747
rect 30616 11716 31217 11744
rect 30616 11704 30622 11716
rect 31205 11713 31217 11716
rect 31251 11713 31263 11747
rect 31312 11744 31340 11784
rect 32398 11772 32404 11784
rect 32456 11772 32462 11824
rect 35713 11815 35771 11821
rect 35713 11812 35725 11815
rect 32508 11784 35725 11812
rect 32508 11744 32536 11784
rect 35713 11781 35725 11784
rect 35759 11781 35771 11815
rect 35713 11775 35771 11781
rect 36170 11772 36176 11824
rect 36228 11812 36234 11824
rect 36541 11815 36599 11821
rect 36541 11812 36553 11815
rect 36228 11784 36553 11812
rect 36228 11772 36234 11784
rect 36541 11781 36553 11784
rect 36587 11781 36599 11815
rect 36541 11775 36599 11781
rect 36633 11815 36691 11821
rect 36633 11781 36645 11815
rect 36679 11812 36691 11815
rect 36814 11812 36820 11824
rect 36679 11784 36820 11812
rect 36679 11781 36691 11784
rect 36633 11775 36691 11781
rect 36814 11772 36820 11784
rect 36872 11772 36878 11824
rect 31312 11716 32536 11744
rect 33413 11747 33471 11753
rect 33413 11742 33425 11747
rect 31205 11707 31263 11713
rect 33336 11714 33425 11742
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 17880 11648 18429 11676
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 21910 11676 21916 11688
rect 18656 11648 21916 11676
rect 18656 11636 18662 11648
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 23106 11636 23112 11688
rect 23164 11676 23170 11688
rect 27614 11676 27620 11688
rect 23164 11648 27620 11676
rect 23164 11636 23170 11648
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 27893 11679 27951 11685
rect 27893 11676 27905 11679
rect 27856 11648 27905 11676
rect 27856 11636 27862 11648
rect 27893 11645 27905 11648
rect 27939 11645 27951 11679
rect 28074 11676 28080 11688
rect 28035 11648 28080 11676
rect 27893 11639 27951 11645
rect 16390 11608 16396 11620
rect 15672 11580 16396 11608
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 16853 11611 16911 11617
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 17862 11608 17868 11620
rect 16899 11580 17868 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 18049 11611 18107 11617
rect 18049 11577 18061 11611
rect 18095 11608 18107 11611
rect 18690 11608 18696 11620
rect 18095 11580 18696 11608
rect 18095 11577 18107 11580
rect 18049 11571 18107 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 20438 11608 20444 11620
rect 18840 11580 20444 11608
rect 18840 11568 18846 11580
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 24302 11568 24308 11620
rect 24360 11608 24366 11620
rect 27908 11608 27936 11639
rect 28074 11636 28080 11648
rect 28132 11636 28138 11688
rect 29178 11636 29184 11688
rect 29236 11676 29242 11688
rect 31294 11676 31300 11688
rect 29236 11648 31300 11676
rect 29236 11636 29242 11648
rect 31294 11636 31300 11648
rect 31352 11636 31358 11688
rect 31386 11636 31392 11688
rect 31444 11676 31450 11688
rect 31444 11648 31489 11676
rect 31444 11636 31450 11648
rect 31570 11636 31576 11688
rect 31628 11676 31634 11688
rect 33042 11676 33048 11688
rect 31628 11648 33048 11676
rect 31628 11636 31634 11648
rect 33042 11636 33048 11648
rect 33100 11676 33106 11688
rect 33229 11679 33287 11685
rect 33229 11676 33241 11679
rect 33100 11648 33241 11676
rect 33100 11636 33106 11648
rect 33229 11645 33241 11648
rect 33275 11645 33287 11679
rect 33229 11639 33287 11645
rect 28534 11608 28540 11620
rect 24360 11580 27844 11608
rect 27908 11580 28540 11608
rect 24360 11568 24366 11580
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12860 11512 12909 11540
rect 12860 11500 12866 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11540 13323 11543
rect 15102 11540 15108 11552
rect 13311 11512 15108 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 16255 11512 17417 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 17405 11509 17417 11512
rect 17451 11540 17463 11543
rect 20070 11540 20076 11552
rect 17451 11512 20076 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 24762 11540 24768 11552
rect 20312 11512 24768 11540
rect 20312 11500 20318 11512
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 27430 11540 27436 11552
rect 27391 11512 27436 11540
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27816 11540 27844 11580
rect 28534 11568 28540 11580
rect 28592 11568 28598 11620
rect 29822 11568 29828 11620
rect 29880 11608 29886 11620
rect 30098 11608 30104 11620
rect 29880 11580 30104 11608
rect 29880 11568 29886 11580
rect 30098 11568 30104 11580
rect 30156 11568 30162 11620
rect 32398 11568 32404 11620
rect 32456 11608 32462 11620
rect 33336 11608 33364 11714
rect 33413 11713 33425 11714
rect 33459 11713 33471 11747
rect 33413 11707 33471 11713
rect 34330 11704 34336 11756
rect 34388 11744 34394 11756
rect 34425 11747 34483 11753
rect 34425 11744 34437 11747
rect 34388 11716 34437 11744
rect 34388 11704 34394 11716
rect 34425 11713 34437 11716
rect 34471 11713 34483 11747
rect 34425 11707 34483 11713
rect 34532 11716 35287 11744
rect 34532 11685 34560 11716
rect 34517 11679 34575 11685
rect 34517 11676 34529 11679
rect 33428 11648 34529 11676
rect 33428 11620 33456 11648
rect 34517 11645 34529 11648
rect 34563 11645 34575 11679
rect 34517 11639 34575 11645
rect 34701 11679 34759 11685
rect 34701 11645 34713 11679
rect 34747 11676 34759 11679
rect 34882 11676 34888 11688
rect 34747 11648 34888 11676
rect 34747 11645 34759 11648
rect 34701 11639 34759 11645
rect 34882 11636 34888 11648
rect 34940 11636 34946 11688
rect 35259 11676 35287 11716
rect 35342 11704 35348 11756
rect 35400 11744 35406 11756
rect 35400 11716 35445 11744
rect 35400 11704 35406 11716
rect 36262 11704 36268 11756
rect 36320 11744 36326 11756
rect 36357 11747 36415 11753
rect 36357 11744 36369 11747
rect 36320 11716 36369 11744
rect 36320 11704 36326 11716
rect 36357 11713 36369 11716
rect 36403 11713 36415 11747
rect 36357 11707 36415 11713
rect 36725 11747 36783 11753
rect 36725 11713 36737 11747
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 36078 11676 36084 11688
rect 35259 11648 36084 11676
rect 36078 11636 36084 11648
rect 36136 11636 36142 11688
rect 32456 11580 33364 11608
rect 32456 11568 32462 11580
rect 33410 11568 33416 11620
rect 33468 11568 33474 11620
rect 34054 11568 34060 11620
rect 34112 11608 34118 11620
rect 36262 11608 36268 11620
rect 34112 11580 36268 11608
rect 34112 11568 34118 11580
rect 36262 11568 36268 11580
rect 36320 11568 36326 11620
rect 30650 11540 30656 11552
rect 27816 11512 30656 11540
rect 30650 11500 30656 11512
rect 30708 11500 30714 11552
rect 30834 11540 30840 11552
rect 30795 11512 30840 11540
rect 30834 11500 30840 11512
rect 30892 11500 30898 11552
rect 30926 11500 30932 11552
rect 30984 11540 30990 11552
rect 32677 11543 32735 11549
rect 32677 11540 32689 11543
rect 30984 11512 32689 11540
rect 30984 11500 30990 11512
rect 32677 11509 32689 11512
rect 32723 11540 32735 11543
rect 33318 11540 33324 11552
rect 32723 11512 33324 11540
rect 32723 11509 32735 11512
rect 32677 11503 32735 11509
rect 33318 11500 33324 11512
rect 33376 11500 33382 11552
rect 33594 11500 33600 11552
rect 33652 11540 33658 11552
rect 35342 11540 35348 11552
rect 33652 11512 35348 11540
rect 33652 11500 33658 11512
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 35434 11500 35440 11552
rect 35492 11540 35498 11552
rect 36740 11540 36768 11707
rect 37274 11704 37280 11756
rect 37332 11744 37338 11756
rect 37717 11747 37775 11753
rect 37717 11744 37729 11747
rect 37332 11716 37729 11744
rect 37332 11704 37338 11716
rect 37717 11713 37729 11716
rect 37763 11713 37775 11747
rect 37717 11707 37775 11713
rect 38562 11704 38568 11756
rect 38620 11744 38626 11756
rect 39316 11753 39344 11852
rect 39666 11840 39672 11892
rect 39724 11880 39730 11892
rect 39945 11883 40003 11889
rect 39945 11880 39957 11883
rect 39724 11852 39957 11880
rect 39724 11840 39730 11852
rect 39945 11849 39957 11852
rect 39991 11849 40003 11883
rect 39945 11843 40003 11849
rect 41509 11883 41567 11889
rect 41509 11849 41521 11883
rect 41555 11880 41567 11883
rect 41874 11880 41880 11892
rect 41555 11852 41880 11880
rect 41555 11849 41567 11852
rect 41509 11843 41567 11849
rect 41874 11840 41880 11852
rect 41932 11840 41938 11892
rect 42334 11840 42340 11892
rect 42392 11880 42398 11892
rect 42978 11880 42984 11892
rect 42392 11852 42984 11880
rect 42392 11840 42398 11852
rect 42978 11840 42984 11852
rect 43036 11840 43042 11892
rect 43070 11840 43076 11892
rect 43128 11880 43134 11892
rect 43993 11883 44051 11889
rect 43993 11880 44005 11883
rect 43128 11852 44005 11880
rect 43128 11840 43134 11852
rect 43993 11849 44005 11852
rect 44039 11849 44051 11883
rect 43993 11843 44051 11849
rect 40678 11812 40684 11824
rect 40236 11784 40684 11812
rect 39301 11747 39359 11753
rect 38620 11716 38700 11744
rect 38620 11704 38626 11716
rect 37366 11636 37372 11688
rect 37424 11676 37430 11688
rect 37461 11679 37519 11685
rect 37461 11676 37473 11679
rect 37424 11648 37473 11676
rect 37424 11636 37430 11648
rect 37461 11645 37473 11648
rect 37507 11645 37519 11679
rect 38672 11676 38700 11716
rect 39301 11713 39313 11747
rect 39347 11713 39359 11747
rect 39301 11707 39359 11713
rect 39485 11747 39543 11753
rect 39485 11713 39497 11747
rect 39531 11744 39543 11747
rect 39574 11744 39580 11756
rect 39531 11716 39580 11744
rect 39531 11713 39543 11716
rect 39485 11707 39543 11713
rect 39574 11704 39580 11716
rect 39632 11704 39638 11756
rect 40126 11744 40132 11756
rect 40087 11716 40132 11744
rect 40126 11704 40132 11716
rect 40184 11704 40190 11756
rect 40236 11753 40264 11784
rect 40678 11772 40684 11784
rect 40736 11772 40742 11824
rect 41233 11815 41291 11821
rect 41233 11781 41245 11815
rect 41279 11812 41291 11815
rect 41414 11812 41420 11824
rect 41279 11784 41420 11812
rect 41279 11781 41291 11784
rect 41233 11775 41291 11781
rect 41414 11772 41420 11784
rect 41472 11772 41478 11824
rect 42886 11821 42892 11824
rect 42880 11812 42892 11821
rect 42847 11784 42892 11812
rect 42880 11775 42892 11784
rect 42886 11772 42892 11775
rect 42944 11772 42950 11824
rect 43162 11772 43168 11824
rect 43220 11812 43226 11824
rect 50890 11812 50896 11824
rect 43220 11784 50896 11812
rect 43220 11772 43226 11784
rect 50890 11772 50896 11784
rect 50948 11772 50954 11824
rect 40221 11747 40279 11753
rect 40221 11713 40233 11747
rect 40267 11713 40279 11747
rect 40221 11707 40279 11713
rect 40310 11704 40316 11756
rect 40368 11744 40374 11756
rect 40405 11747 40463 11753
rect 40405 11744 40417 11747
rect 40368 11716 40417 11744
rect 40368 11704 40374 11716
rect 40405 11713 40417 11716
rect 40451 11713 40463 11747
rect 40405 11707 40463 11713
rect 40494 11704 40500 11756
rect 40552 11744 40558 11756
rect 40957 11747 41015 11753
rect 40957 11744 40969 11747
rect 40552 11716 40597 11744
rect 40696 11716 40969 11744
rect 40552 11704 40558 11716
rect 39393 11679 39451 11685
rect 39393 11676 39405 11679
rect 38672 11648 39405 11676
rect 37461 11639 37519 11645
rect 39393 11645 39405 11648
rect 39439 11645 39451 11679
rect 39393 11639 39451 11645
rect 40586 11636 40592 11688
rect 40644 11676 40650 11688
rect 40696 11676 40724 11716
rect 40957 11713 40969 11716
rect 41003 11713 41015 11747
rect 41138 11744 41144 11756
rect 41099 11716 41144 11744
rect 40957 11707 41015 11713
rect 41138 11704 41144 11716
rect 41196 11704 41202 11756
rect 41325 11747 41383 11753
rect 41325 11713 41337 11747
rect 41371 11744 41383 11747
rect 42334 11744 42340 11756
rect 41371 11716 42340 11744
rect 41371 11713 41383 11716
rect 41325 11707 41383 11713
rect 40644 11648 40724 11676
rect 40644 11636 40650 11648
rect 40770 11636 40776 11688
rect 40828 11676 40834 11688
rect 41340 11676 41368 11707
rect 42334 11704 42340 11716
rect 42392 11704 42398 11756
rect 42613 11747 42671 11753
rect 42613 11713 42625 11747
rect 42659 11744 42671 11747
rect 42702 11744 42708 11756
rect 42659 11716 42708 11744
rect 42659 11713 42671 11716
rect 42613 11707 42671 11713
rect 42702 11704 42708 11716
rect 42760 11704 42766 11756
rect 43438 11704 43444 11756
rect 43496 11744 43502 11756
rect 43714 11744 43720 11756
rect 43496 11716 43720 11744
rect 43496 11704 43502 11716
rect 43714 11704 43720 11716
rect 43772 11704 43778 11756
rect 58066 11744 58072 11756
rect 58027 11716 58072 11744
rect 58066 11704 58072 11716
rect 58124 11704 58130 11756
rect 40828 11648 41368 11676
rect 40828 11636 40834 11648
rect 38562 11568 38568 11620
rect 38620 11608 38626 11620
rect 42334 11608 42340 11620
rect 38620 11580 42340 11608
rect 38620 11568 38626 11580
rect 42334 11568 42340 11580
rect 42392 11568 42398 11620
rect 43548 11580 51074 11608
rect 35492 11512 36768 11540
rect 36909 11543 36967 11549
rect 35492 11500 35498 11512
rect 36909 11509 36921 11543
rect 36955 11540 36967 11543
rect 38746 11540 38752 11552
rect 36955 11512 38752 11540
rect 36955 11509 36967 11512
rect 36909 11503 36967 11509
rect 38746 11500 38752 11512
rect 38804 11500 38810 11552
rect 38838 11500 38844 11552
rect 38896 11540 38902 11552
rect 38896 11512 38941 11540
rect 38896 11500 38902 11512
rect 42610 11500 42616 11552
rect 42668 11540 42674 11552
rect 43548 11540 43576 11580
rect 42668 11512 43576 11540
rect 51046 11540 51074 11580
rect 58253 11543 58311 11549
rect 58253 11540 58265 11543
rect 51046 11512 58265 11540
rect 42668 11500 42674 11512
rect 58253 11509 58265 11512
rect 58299 11509 58311 11543
rect 58253 11503 58311 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 13630 11336 13636 11348
rect 12860 11308 13492 11336
rect 13591 11308 13636 11336
rect 12860 11296 12866 11308
rect 13464 11277 13492 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14734 11336 14740 11348
rect 14695 11308 14740 11336
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 16758 11296 16764 11348
rect 16816 11336 16822 11348
rect 17494 11336 17500 11348
rect 16816 11308 17500 11336
rect 16816 11296 16822 11308
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18874 11336 18880 11348
rect 18835 11308 18880 11336
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 19306 11308 25973 11336
rect 12621 11271 12679 11277
rect 12621 11237 12633 11271
rect 12667 11268 12679 11271
rect 13449 11271 13507 11277
rect 12667 11240 13124 11268
rect 12667 11237 12679 11240
rect 12621 11231 12679 11237
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 13096 11200 13124 11240
rect 13449 11237 13461 11271
rect 13495 11237 13507 11271
rect 19306 11268 19334 11308
rect 25961 11305 25973 11308
rect 26007 11336 26019 11339
rect 27246 11336 27252 11348
rect 26007 11308 27252 11336
rect 26007 11305 26019 11308
rect 25961 11299 26019 11305
rect 27246 11296 27252 11308
rect 27304 11296 27310 11348
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 37182 11336 37188 11348
rect 27488 11308 37188 11336
rect 27488 11296 27494 11308
rect 37182 11296 37188 11308
rect 37240 11296 37246 11348
rect 37366 11336 37372 11348
rect 37327 11308 37372 11336
rect 37366 11296 37372 11308
rect 37424 11296 37430 11348
rect 37734 11296 37740 11348
rect 37792 11336 37798 11348
rect 39025 11339 39083 11345
rect 39025 11336 39037 11339
rect 37792 11308 39037 11336
rect 37792 11296 37798 11308
rect 39025 11305 39037 11308
rect 39071 11305 39083 11339
rect 39025 11299 39083 11305
rect 39390 11296 39396 11348
rect 39448 11336 39454 11348
rect 39448 11308 57928 11336
rect 39448 11296 39454 11308
rect 21726 11268 21732 11280
rect 13449 11231 13507 11237
rect 15028 11240 19334 11268
rect 20732 11240 21732 11268
rect 13538 11200 13544 11212
rect 12308 11172 12756 11200
rect 13096 11172 13544 11200
rect 12308 11160 12314 11172
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 7558 11132 7564 11144
rect 1627 11104 7564 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 12124 11104 12541 11132
rect 12124 11092 12130 11104
rect 12529 11101 12541 11104
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12728 11141 12756 11172
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 15028 11209 15056 11240
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 14608 11172 14933 11200
rect 14608 11160 14614 11172
rect 14921 11169 14933 11172
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11200 15255 11203
rect 16298 11200 16304 11212
rect 15243 11172 16304 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 18380 11172 18521 11200
rect 18380 11160 18386 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 20254 11200 20260 11212
rect 18509 11163 18567 11169
rect 18708 11172 20260 11200
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11132 15163 11135
rect 15151 11104 15240 11132
rect 15151 11101 15163 11104
rect 15105 11095 15163 11101
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 14826 11064 14832 11076
rect 13219 11036 14832 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 15212 11064 15240 11104
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15344 11104 15761 11132
rect 15344 11092 15350 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 18708 11141 18736 11172
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 16264 11104 18705 11132
rect 16264 11092 16270 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19426 11132 19432 11144
rect 18932 11104 19432 11132
rect 18932 11092 18938 11104
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20070 11132 20076 11144
rect 20031 11104 20076 11132
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 20533 11135 20591 11141
rect 20533 11101 20545 11135
rect 20579 11132 20591 11135
rect 20732 11132 20760 11240
rect 21726 11228 21732 11240
rect 21784 11268 21790 11280
rect 24486 11268 24492 11280
rect 21784 11240 24492 11268
rect 21784 11228 21790 11240
rect 24486 11228 24492 11240
rect 24544 11228 24550 11280
rect 27614 11268 27620 11280
rect 27575 11240 27620 11268
rect 27614 11228 27620 11240
rect 27672 11228 27678 11280
rect 30006 11268 30012 11280
rect 28184 11240 30012 11268
rect 22094 11200 22100 11212
rect 21192 11172 22100 11200
rect 20579 11104 20760 11132
rect 20809 11135 20867 11141
rect 20579 11101 20591 11104
rect 20533 11095 20591 11101
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 21082 11132 21088 11144
rect 20855 11104 21088 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21192 11141 21220 11172
rect 22094 11160 22100 11172
rect 22152 11160 22158 11212
rect 25590 11160 25596 11212
rect 25648 11200 25654 11212
rect 27522 11200 27528 11212
rect 25648 11172 27528 11200
rect 25648 11160 25654 11172
rect 27522 11160 27528 11172
rect 27580 11200 27586 11212
rect 28184 11200 28212 11240
rect 30006 11228 30012 11240
rect 30064 11228 30070 11280
rect 33318 11228 33324 11280
rect 33376 11228 33382 11280
rect 33502 11228 33508 11280
rect 33560 11268 33566 11280
rect 33597 11271 33655 11277
rect 33597 11268 33609 11271
rect 33560 11240 33609 11268
rect 33560 11228 33566 11240
rect 33597 11237 33609 11240
rect 33643 11237 33655 11271
rect 33597 11231 33655 11237
rect 33870 11228 33876 11280
rect 33928 11268 33934 11280
rect 34241 11271 34299 11277
rect 34241 11268 34253 11271
rect 33928 11240 34253 11268
rect 33928 11228 33934 11240
rect 34241 11237 34253 11240
rect 34287 11237 34299 11271
rect 34241 11231 34299 11237
rect 36449 11271 36507 11277
rect 36449 11237 36461 11271
rect 36495 11268 36507 11271
rect 36722 11268 36728 11280
rect 36495 11240 36728 11268
rect 36495 11237 36507 11240
rect 36449 11231 36507 11237
rect 36722 11228 36728 11240
rect 36780 11228 36786 11280
rect 37090 11268 37096 11280
rect 37016 11240 37096 11268
rect 27580 11172 28212 11200
rect 27580 11160 27586 11172
rect 28258 11160 28264 11212
rect 28316 11200 28322 11212
rect 28718 11200 28724 11212
rect 28316 11172 28724 11200
rect 28316 11160 28322 11172
rect 28718 11160 28724 11172
rect 28776 11160 28782 11212
rect 33336 11200 33364 11228
rect 33778 11200 33784 11212
rect 33336 11172 33784 11200
rect 33778 11160 33784 11172
rect 33836 11160 33842 11212
rect 34790 11160 34796 11212
rect 34848 11200 34854 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34848 11172 34897 11200
rect 34848 11160 34854 11172
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 35802 11200 35808 11212
rect 34885 11163 34943 11169
rect 34992 11172 35808 11200
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11132 21327 11135
rect 21542 11132 21548 11144
rect 21315 11104 21548 11132
rect 21315 11101 21327 11104
rect 21269 11095 21327 11101
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 21775 11104 22140 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 15378 11064 15384 11076
rect 15212 11036 15384 11064
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 21910 11064 21916 11076
rect 17276 11036 21916 11064
rect 17276 11024 17282 11036
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 22112 11064 22140 11104
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 24486 11132 24492 11144
rect 22244 11104 24492 11132
rect 22244 11092 22250 11104
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 25222 11132 25228 11144
rect 24627 11104 25228 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 26421 11135 26479 11141
rect 26421 11101 26433 11135
rect 26467 11132 26479 11135
rect 28902 11132 28908 11144
rect 26467 11104 28908 11132
rect 26467 11101 26479 11104
rect 26421 11095 26479 11101
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 30098 11092 30104 11144
rect 30156 11132 30162 11144
rect 30285 11135 30343 11141
rect 30285 11132 30297 11135
rect 30156 11104 30297 11132
rect 30156 11092 30162 11104
rect 30285 11101 30297 11104
rect 30331 11132 30343 11135
rect 31018 11132 31024 11144
rect 30331 11104 31024 11132
rect 30331 11101 30343 11104
rect 30285 11095 30343 11101
rect 31018 11092 31024 11104
rect 31076 11132 31082 11144
rect 32217 11135 32275 11141
rect 32217 11132 32229 11135
rect 31076 11104 32229 11132
rect 31076 11092 31082 11104
rect 32217 11101 32229 11104
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 32306 11092 32312 11144
rect 32364 11132 32370 11144
rect 32473 11135 32531 11141
rect 32473 11132 32485 11135
rect 32364 11104 32485 11132
rect 32364 11092 32370 11104
rect 32473 11101 32485 11104
rect 32519 11101 32531 11135
rect 32473 11095 32531 11101
rect 33318 11092 33324 11144
rect 33376 11132 33382 11144
rect 34057 11135 34115 11141
rect 34057 11132 34069 11135
rect 33376 11104 34069 11132
rect 33376 11092 33382 11104
rect 34057 11101 34069 11104
rect 34103 11132 34115 11135
rect 34422 11132 34428 11144
rect 34103 11104 34428 11132
rect 34103 11101 34115 11104
rect 34057 11095 34115 11101
rect 34422 11092 34428 11104
rect 34480 11092 34486 11144
rect 24848 11067 24906 11073
rect 22112 11036 24808 11064
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 16945 10999 17003 11005
rect 16945 10996 16957 10999
rect 14792 10968 16957 10996
rect 14792 10956 14798 10968
rect 16945 10965 16957 10968
rect 16991 10965 17003 10999
rect 16945 10959 17003 10965
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 22925 10999 22983 11005
rect 22925 10996 22937 10999
rect 17092 10968 22937 10996
rect 17092 10956 17098 10968
rect 22925 10965 22937 10968
rect 22971 10965 22983 10999
rect 24780 10996 24808 11036
rect 24848 11033 24860 11067
rect 24894 11064 24906 11067
rect 24946 11064 24952 11076
rect 24894 11036 24952 11064
rect 24894 11033 24906 11036
rect 24848 11027 24906 11033
rect 24946 11024 24952 11036
rect 25004 11024 25010 11076
rect 29086 11064 29092 11076
rect 25332 11036 29092 11064
rect 25332 10996 25360 11036
rect 29086 11024 29092 11036
rect 29144 11024 29150 11076
rect 30552 11067 30610 11073
rect 30552 11033 30564 11067
rect 30598 11064 30610 11067
rect 34992 11064 35020 11172
rect 35802 11160 35808 11172
rect 35860 11160 35866 11212
rect 37016 11209 37044 11240
rect 37090 11228 37096 11240
rect 37148 11228 37154 11280
rect 37274 11228 37280 11280
rect 37332 11268 37338 11280
rect 38010 11268 38016 11280
rect 37332 11240 38016 11268
rect 37332 11228 37338 11240
rect 38010 11228 38016 11240
rect 38068 11268 38074 11280
rect 38838 11268 38844 11280
rect 38068 11240 38844 11268
rect 38068 11228 38074 11240
rect 38838 11228 38844 11240
rect 38896 11228 38902 11280
rect 40678 11268 40684 11280
rect 40512 11240 40684 11268
rect 37001 11203 37059 11209
rect 37001 11169 37013 11203
rect 37047 11169 37059 11203
rect 38197 11203 38255 11209
rect 38197 11200 38209 11203
rect 37001 11163 37059 11169
rect 37108 11172 38209 11200
rect 35161 11135 35219 11141
rect 35161 11101 35173 11135
rect 35207 11132 35219 11135
rect 36906 11132 36912 11144
rect 35207 11104 36912 11132
rect 35207 11101 35219 11104
rect 35161 11095 35219 11101
rect 36906 11092 36912 11104
rect 36964 11092 36970 11144
rect 36722 11064 36728 11076
rect 30598 11036 35020 11064
rect 35820 11036 36728 11064
rect 30598 11033 30610 11036
rect 30552 11027 30610 11033
rect 24780 10968 25360 10996
rect 22925 10959 22983 10965
rect 26602 10956 26608 11008
rect 26660 10996 26666 11008
rect 29362 10996 29368 11008
rect 26660 10968 29368 10996
rect 26660 10956 26666 10968
rect 29362 10956 29368 10968
rect 29420 10956 29426 11008
rect 30650 10956 30656 11008
rect 30708 10996 30714 11008
rect 31110 10996 31116 11008
rect 30708 10968 31116 10996
rect 30708 10956 30714 10968
rect 31110 10956 31116 10968
rect 31168 10996 31174 11008
rect 31665 10999 31723 11005
rect 31665 10996 31677 10999
rect 31168 10968 31677 10996
rect 31168 10956 31174 10968
rect 31665 10965 31677 10968
rect 31711 10996 31723 10999
rect 32674 10996 32680 11008
rect 31711 10968 32680 10996
rect 31711 10965 31723 10968
rect 31665 10959 31723 10965
rect 32674 10956 32680 10968
rect 32732 10956 32738 11008
rect 32950 10956 32956 11008
rect 33008 10996 33014 11008
rect 33318 10996 33324 11008
rect 33008 10968 33324 10996
rect 33008 10956 33014 10968
rect 33318 10956 33324 10968
rect 33376 10956 33382 11008
rect 34514 10956 34520 11008
rect 34572 10996 34578 11008
rect 35820 10996 35848 11036
rect 36722 11024 36728 11036
rect 36780 11024 36786 11076
rect 34572 10968 35848 10996
rect 34572 10956 34578 10968
rect 35986 10956 35992 11008
rect 36044 10996 36050 11008
rect 37108 10996 37136 11172
rect 38197 11169 38209 11172
rect 38243 11169 38255 11203
rect 38197 11163 38255 11169
rect 38286 11160 38292 11212
rect 38344 11200 38350 11212
rect 38657 11203 38715 11209
rect 38657 11200 38669 11203
rect 38344 11172 38669 11200
rect 38344 11160 38350 11172
rect 38657 11169 38669 11172
rect 38703 11169 38715 11203
rect 38657 11163 38715 11169
rect 37182 11092 37188 11144
rect 37240 11132 37246 11144
rect 37829 11135 37887 11141
rect 37240 11104 37285 11132
rect 37240 11092 37246 11104
rect 37829 11101 37841 11135
rect 37875 11101 37887 11135
rect 38010 11132 38016 11144
rect 37971 11104 38016 11132
rect 37829 11095 37887 11101
rect 37844 11064 37872 11095
rect 38010 11092 38016 11104
rect 38068 11092 38074 11144
rect 38746 11092 38752 11144
rect 38804 11132 38810 11144
rect 38841 11135 38899 11141
rect 38841 11132 38853 11135
rect 38804 11104 38853 11132
rect 38804 11092 38810 11104
rect 38841 11101 38853 11104
rect 38887 11101 38899 11135
rect 38841 11095 38899 11101
rect 40405 11135 40463 11141
rect 40405 11101 40417 11135
rect 40451 11132 40463 11135
rect 40512 11132 40540 11240
rect 40678 11228 40684 11240
rect 40736 11228 40742 11280
rect 40957 11271 41015 11277
rect 40957 11237 40969 11271
rect 41003 11268 41015 11271
rect 43622 11268 43628 11280
rect 41003 11240 43628 11268
rect 41003 11237 41015 11240
rect 40957 11231 41015 11237
rect 43622 11228 43628 11240
rect 43680 11228 43686 11280
rect 54202 11268 54208 11280
rect 43916 11240 51074 11268
rect 41138 11200 41144 11212
rect 40451 11104 40540 11132
rect 40604 11172 41144 11200
rect 40451 11101 40463 11104
rect 40405 11095 40463 11101
rect 37246 11036 37872 11064
rect 37246 11008 37274 11036
rect 38930 11024 38936 11076
rect 38988 11064 38994 11076
rect 40604 11073 40632 11172
rect 41138 11160 41144 11172
rect 41196 11160 41202 11212
rect 43916 11200 43944 11240
rect 41708 11172 43944 11200
rect 51046 11200 51074 11240
rect 52656 11240 54208 11268
rect 52454 11200 52460 11212
rect 51046 11172 52460 11200
rect 40770 11132 40776 11144
rect 40731 11104 40776 11132
rect 40770 11092 40776 11104
rect 40828 11092 40834 11144
rect 41708 11141 41736 11172
rect 52454 11160 52460 11172
rect 52512 11160 52518 11212
rect 41693 11135 41751 11141
rect 41693 11101 41705 11135
rect 41739 11101 41751 11135
rect 43162 11132 43168 11144
rect 41693 11095 41751 11101
rect 42720 11104 43168 11132
rect 40589 11067 40647 11073
rect 40589 11064 40601 11067
rect 38988 11036 40601 11064
rect 38988 11024 38994 11036
rect 40589 11033 40601 11036
rect 40635 11033 40647 11067
rect 40589 11027 40647 11033
rect 40681 11067 40739 11073
rect 40681 11033 40693 11067
rect 40727 11064 40739 11067
rect 42720 11064 42748 11104
rect 43162 11092 43168 11104
rect 43220 11092 43226 11144
rect 43254 11092 43260 11144
rect 43312 11132 43318 11144
rect 43901 11135 43959 11141
rect 43901 11132 43913 11135
rect 43312 11104 43913 11132
rect 43312 11092 43318 11104
rect 43901 11101 43913 11104
rect 43947 11101 43959 11135
rect 44082 11132 44088 11144
rect 44043 11104 44088 11132
rect 43901 11095 43959 11101
rect 44082 11092 44088 11104
rect 44140 11092 44146 11144
rect 52656 11141 52684 11240
rect 54202 11228 54208 11240
rect 54260 11228 54266 11280
rect 52730 11160 52736 11212
rect 52788 11200 52794 11212
rect 54478 11200 54484 11212
rect 52788 11172 54484 11200
rect 52788 11160 52794 11172
rect 54478 11160 54484 11172
rect 54536 11160 54542 11212
rect 44269 11135 44327 11141
rect 44269 11132 44281 11135
rect 44192 11104 44281 11132
rect 43438 11064 43444 11076
rect 40727 11036 42748 11064
rect 43399 11036 43444 11064
rect 40727 11033 40739 11036
rect 40681 11027 40739 11033
rect 43438 11024 43444 11036
rect 43496 11024 43502 11076
rect 43622 11024 43628 11076
rect 43680 11064 43686 11076
rect 44192 11064 44220 11104
rect 44269 11101 44281 11104
rect 44315 11101 44327 11135
rect 44269 11095 44327 11101
rect 52641 11135 52699 11141
rect 52641 11101 52653 11135
rect 52687 11101 52699 11135
rect 52641 11095 52699 11101
rect 52822 11092 52828 11144
rect 52880 11132 52886 11144
rect 52880 11104 52925 11132
rect 52880 11092 52886 11104
rect 53006 11092 53012 11144
rect 53064 11132 53070 11144
rect 57900 11141 57928 11308
rect 57885 11135 57943 11141
rect 53064 11104 53109 11132
rect 53064 11092 53070 11104
rect 57885 11101 57897 11135
rect 57931 11101 57943 11135
rect 57885 11095 57943 11101
rect 43680 11036 44220 11064
rect 43680 11024 43686 11036
rect 46198 11024 46204 11076
rect 46256 11064 46262 11076
rect 50614 11064 50620 11076
rect 46256 11036 50620 11064
rect 46256 11024 46262 11036
rect 50614 11024 50620 11036
rect 50672 11024 50678 11076
rect 52913 11067 52971 11073
rect 52913 11033 52925 11067
rect 52959 11064 52971 11067
rect 53098 11064 53104 11076
rect 52959 11036 53104 11064
rect 52959 11033 52971 11036
rect 52913 11027 52971 11033
rect 53098 11024 53104 11036
rect 53156 11024 53162 11076
rect 58161 11067 58219 11073
rect 58161 11064 58173 11067
rect 57900 11036 58173 11064
rect 57900 11008 57928 11036
rect 58161 11033 58173 11036
rect 58207 11033 58219 11067
rect 58161 11027 58219 11033
rect 36044 10968 37136 10996
rect 36044 10956 36050 10968
rect 37182 10956 37188 11008
rect 37240 10968 37274 11008
rect 37240 10956 37246 10968
rect 37366 10956 37372 11008
rect 37424 10996 37430 11008
rect 53193 10999 53251 11005
rect 53193 10996 53205 10999
rect 37424 10968 53205 10996
rect 37424 10956 37430 10968
rect 53193 10965 53205 10968
rect 53239 10965 53251 10999
rect 53193 10959 53251 10965
rect 57882 10956 57888 11008
rect 57940 10956 57946 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 14277 10795 14335 10801
rect 7616 10764 14228 10792
rect 7616 10752 7622 10764
rect 13354 10724 13360 10736
rect 13315 10696 13360 10724
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 13906 10724 13912 10736
rect 13867 10696 13912 10724
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 14090 10684 14096 10736
rect 14148 10733 14154 10736
rect 14148 10727 14167 10733
rect 14155 10693 14167 10727
rect 14148 10687 14167 10693
rect 14148 10684 14154 10687
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 13136 10628 13277 10656
rect 13136 10616 13142 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 13464 10520 13492 10619
rect 14200 10588 14228 10764
rect 14277 10761 14289 10795
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 14292 10724 14320 10755
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15010 10792 15016 10804
rect 14884 10764 15016 10792
rect 14884 10752 14890 10764
rect 15010 10752 15016 10764
rect 15068 10792 15074 10804
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 15068 10764 15117 10792
rect 15068 10752 15074 10764
rect 15105 10761 15117 10764
rect 15151 10792 15163 10795
rect 15378 10792 15384 10804
rect 15151 10764 15384 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 19150 10792 19156 10804
rect 15528 10764 19156 10792
rect 15528 10752 15534 10764
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 22370 10792 22376 10804
rect 19260 10764 22376 10792
rect 19260 10724 19288 10764
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 22830 10752 22836 10804
rect 22888 10792 22894 10804
rect 24949 10795 25007 10801
rect 24949 10792 24961 10795
rect 22888 10764 24961 10792
rect 22888 10752 22894 10764
rect 24949 10761 24961 10764
rect 24995 10761 25007 10795
rect 29086 10792 29092 10804
rect 29047 10764 29092 10792
rect 24949 10755 25007 10761
rect 29086 10752 29092 10764
rect 29144 10752 29150 10804
rect 29362 10752 29368 10804
rect 29420 10792 29426 10804
rect 30558 10792 30564 10804
rect 29420 10764 30564 10792
rect 29420 10752 29426 10764
rect 30558 10752 30564 10764
rect 30616 10752 30622 10804
rect 30837 10795 30895 10801
rect 30837 10761 30849 10795
rect 30883 10761 30895 10795
rect 30837 10755 30895 10761
rect 14292 10696 18092 10724
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14332 10628 14749 10656
rect 14332 10616 14338 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14884 10628 14933 10656
rect 14884 10616 14890 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 15059 10659 15117 10665
rect 15059 10625 15071 10659
rect 15105 10656 15117 10659
rect 15194 10656 15200 10668
rect 15105 10628 15200 10656
rect 15105 10625 15117 10628
rect 15059 10619 15117 10625
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15746 10656 15752 10668
rect 15344 10628 15389 10656
rect 15707 10628 15752 10656
rect 15344 10616 15350 10628
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15896 10628 15945 10656
rect 15896 10616 15902 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16040 10588 16068 10619
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16850 10656 16856 10668
rect 16172 10628 16217 10656
rect 16811 10628 16856 10656
rect 16172 10616 16178 10628
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 18064 10665 18092 10696
rect 18156 10696 19288 10724
rect 18063 10659 18121 10665
rect 17000 10628 17172 10656
rect 17000 10616 17006 10628
rect 14200 10560 16068 10588
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 17034 10588 17040 10600
rect 16264 10560 17040 10588
rect 16264 10548 16270 10560
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17144 10588 17172 10628
rect 18063 10625 18075 10659
rect 18109 10625 18121 10659
rect 18063 10619 18121 10625
rect 18156 10588 18184 10696
rect 20070 10684 20076 10736
rect 20128 10724 20134 10736
rect 20898 10724 20904 10736
rect 20128 10696 20904 10724
rect 20128 10684 20134 10696
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 21324 10696 23612 10724
rect 21324 10684 21330 10696
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 18380 10628 18521 10656
rect 18380 10616 18386 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 19153 10659 19211 10665
rect 19153 10656 19165 10659
rect 19024 10628 19165 10656
rect 19024 10616 19030 10628
rect 19153 10625 19165 10628
rect 19199 10625 19211 10659
rect 19153 10619 19211 10625
rect 19518 10616 19524 10668
rect 19576 10656 19582 10668
rect 20806 10656 20812 10668
rect 19576 10628 20812 10656
rect 19576 10616 19582 10628
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 22186 10656 22192 10668
rect 22099 10628 22192 10656
rect 22186 10616 22192 10628
rect 22244 10656 22250 10668
rect 22646 10656 22652 10668
rect 22244 10628 22652 10656
rect 22244 10616 22250 10628
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 17144 10560 18184 10588
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 18248 10520 18276 10551
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 18472 10560 18613 10588
rect 18472 10548 18478 10560
rect 18601 10557 18613 10560
rect 18647 10588 18659 10591
rect 19702 10588 19708 10600
rect 18647 10560 19708 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 19702 10548 19708 10560
rect 19760 10588 19766 10600
rect 20070 10588 20076 10600
rect 19760 10560 20076 10588
rect 19760 10548 19766 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 22278 10588 22284 10600
rect 20180 10560 22284 10588
rect 20180 10520 20208 10560
rect 22278 10548 22284 10560
rect 22336 10548 22342 10600
rect 22554 10588 22560 10600
rect 22515 10560 22560 10588
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 23474 10520 23480 10532
rect 13464 10492 17724 10520
rect 18248 10492 20208 10520
rect 20272 10492 23480 10520
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10452 14151 10455
rect 15194 10452 15200 10464
rect 14139 10424 15200 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 16301 10455 16359 10461
rect 16301 10452 16313 10455
rect 16264 10424 16313 10452
rect 16264 10412 16270 10424
rect 16301 10421 16313 10424
rect 16347 10421 16359 10455
rect 16301 10415 16359 10421
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17586 10452 17592 10464
rect 17368 10424 17592 10452
rect 17368 10412 17374 10424
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 17696 10452 17724 10492
rect 20272 10452 20300 10492
rect 23474 10480 23480 10492
rect 23532 10480 23538 10532
rect 23584 10520 23612 10696
rect 24026 10684 24032 10736
rect 24084 10724 24090 10736
rect 30852 10724 30880 10755
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31205 10795 31263 10801
rect 31205 10792 31217 10795
rect 31168 10764 31217 10792
rect 31168 10752 31174 10764
rect 31205 10761 31217 10764
rect 31251 10761 31263 10795
rect 31205 10755 31263 10761
rect 31294 10752 31300 10804
rect 31352 10792 31358 10804
rect 32125 10795 32183 10801
rect 31352 10764 31397 10792
rect 31352 10752 31358 10764
rect 32125 10761 32137 10795
rect 32171 10792 32183 10795
rect 32398 10792 32404 10804
rect 32171 10764 32404 10792
rect 32171 10761 32183 10764
rect 32125 10755 32183 10761
rect 32398 10752 32404 10764
rect 32456 10752 32462 10804
rect 33962 10752 33968 10804
rect 34020 10792 34026 10804
rect 34330 10792 34336 10804
rect 34020 10764 34336 10792
rect 34020 10752 34026 10764
rect 34330 10752 34336 10764
rect 34388 10792 34394 10804
rect 34388 10764 34652 10792
rect 34388 10752 34394 10764
rect 32858 10724 32864 10736
rect 24084 10696 28304 10724
rect 30852 10696 32864 10724
rect 24084 10684 24090 10696
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 25038 10656 25044 10668
rect 23799 10628 25044 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 27614 10656 27620 10668
rect 27295 10628 27620 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 28166 10656 28172 10668
rect 27939 10628 28172 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 28166 10616 28172 10628
rect 28224 10616 28230 10668
rect 28276 10656 28304 10696
rect 32858 10684 32864 10696
rect 32916 10684 32922 10736
rect 33134 10724 33140 10736
rect 33095 10696 33140 10724
rect 33134 10684 33140 10696
rect 33192 10724 33198 10736
rect 33873 10727 33931 10733
rect 33873 10724 33885 10727
rect 33192 10696 33885 10724
rect 33192 10684 33198 10696
rect 33873 10693 33885 10696
rect 33919 10693 33931 10727
rect 34514 10724 34520 10736
rect 33873 10687 33931 10693
rect 34348 10696 34520 10724
rect 30558 10656 30564 10668
rect 28276 10628 30564 10656
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 32490 10656 32496 10668
rect 32451 10628 32496 10656
rect 32490 10616 32496 10628
rect 32548 10616 32554 10668
rect 32582 10616 32588 10668
rect 32640 10656 32646 10668
rect 33689 10659 33747 10665
rect 32640 10628 32685 10656
rect 32640 10616 32646 10628
rect 33689 10625 33701 10659
rect 33735 10656 33747 10659
rect 33778 10656 33784 10668
rect 33735 10628 33784 10656
rect 33735 10625 33747 10628
rect 33689 10619 33747 10625
rect 33778 10616 33784 10628
rect 33836 10616 33842 10668
rect 33962 10656 33968 10668
rect 33923 10628 33968 10656
rect 33962 10616 33968 10628
rect 34020 10616 34026 10668
rect 34348 10665 34376 10696
rect 34514 10684 34520 10696
rect 34572 10684 34578 10736
rect 34624 10724 34652 10764
rect 34698 10752 34704 10804
rect 34756 10792 34762 10804
rect 36446 10792 36452 10804
rect 34756 10764 36452 10792
rect 34756 10752 34762 10764
rect 36446 10752 36452 10764
rect 36504 10752 36510 10804
rect 36722 10752 36728 10804
rect 36780 10792 36786 10804
rect 37642 10792 37648 10804
rect 36780 10764 37648 10792
rect 36780 10752 36786 10764
rect 37642 10752 37648 10764
rect 37700 10752 37706 10804
rect 37829 10795 37887 10801
rect 37829 10761 37841 10795
rect 37875 10792 37887 10795
rect 38470 10792 38476 10804
rect 37875 10764 38476 10792
rect 37875 10761 37887 10764
rect 37829 10755 37887 10761
rect 38470 10752 38476 10764
rect 38528 10752 38534 10804
rect 40954 10752 40960 10804
rect 41012 10792 41018 10804
rect 41138 10792 41144 10804
rect 41012 10764 41144 10792
rect 41012 10752 41018 10764
rect 41138 10752 41144 10764
rect 41196 10752 41202 10804
rect 42334 10752 42340 10804
rect 42392 10792 42398 10804
rect 46290 10792 46296 10804
rect 42392 10764 46296 10792
rect 42392 10752 42398 10764
rect 46290 10752 46296 10764
rect 46348 10752 46354 10804
rect 49694 10752 49700 10804
rect 49752 10792 49758 10804
rect 50709 10795 50767 10801
rect 50709 10792 50721 10795
rect 49752 10764 50721 10792
rect 49752 10752 49758 10764
rect 50709 10761 50721 10764
rect 50755 10792 50767 10795
rect 56870 10792 56876 10804
rect 50755 10764 56876 10792
rect 50755 10761 50767 10764
rect 50709 10755 50767 10761
rect 56870 10752 56876 10764
rect 56928 10752 56934 10804
rect 41509 10727 41567 10733
rect 34624 10696 34684 10724
rect 34656 10678 34684 10696
rect 34992 10696 39528 10724
rect 34656 10665 34744 10678
rect 34333 10659 34391 10665
rect 34333 10625 34345 10659
rect 34379 10625 34391 10659
rect 34333 10619 34391 10625
rect 34425 10659 34483 10665
rect 34425 10625 34437 10659
rect 34471 10625 34483 10659
rect 34656 10659 34759 10665
rect 34992 10659 35020 10696
rect 34656 10650 34713 10659
rect 34425 10619 34483 10625
rect 34701 10625 34713 10650
rect 34747 10625 34759 10659
rect 34701 10619 34759 10625
rect 34900 10631 35020 10659
rect 35526 10656 35532 10668
rect 24946 10548 24952 10600
rect 25004 10588 25010 10600
rect 26326 10588 26332 10600
rect 25004 10560 26332 10588
rect 25004 10548 25010 10560
rect 26326 10548 26332 10560
rect 26384 10548 26390 10600
rect 31481 10591 31539 10597
rect 31481 10557 31493 10591
rect 31527 10588 31539 10591
rect 31570 10588 31576 10600
rect 31527 10560 31576 10588
rect 31527 10557 31539 10560
rect 31481 10551 31539 10557
rect 31570 10548 31576 10560
rect 31628 10548 31634 10600
rect 32600 10588 32628 10616
rect 31680 10560 32628 10588
rect 32677 10591 32735 10597
rect 30098 10520 30104 10532
rect 23584 10492 30104 10520
rect 30098 10480 30104 10492
rect 30156 10480 30162 10532
rect 30650 10480 30656 10532
rect 30708 10520 30714 10532
rect 31680 10520 31708 10560
rect 32677 10557 32689 10591
rect 32723 10557 32735 10591
rect 34440 10588 34468 10619
rect 34514 10588 34520 10600
rect 34440 10560 34520 10588
rect 32677 10551 32735 10557
rect 30708 10492 31708 10520
rect 30708 10480 30714 10492
rect 31754 10480 31760 10532
rect 31812 10520 31818 10532
rect 32582 10520 32588 10532
rect 31812 10492 32588 10520
rect 31812 10480 31818 10492
rect 32582 10480 32588 10492
rect 32640 10520 32646 10532
rect 32692 10520 32720 10551
rect 34514 10548 34520 10560
rect 34572 10548 34578 10600
rect 34609 10591 34667 10597
rect 34609 10557 34621 10591
rect 34655 10588 34667 10591
rect 34900 10588 34928 10631
rect 35268 10628 35532 10656
rect 34655 10560 34928 10588
rect 34977 10591 35035 10597
rect 34655 10557 34667 10560
rect 34609 10551 34667 10557
rect 34977 10557 34989 10591
rect 35023 10557 35035 10591
rect 34977 10551 35035 10557
rect 32640 10492 32720 10520
rect 32640 10480 32646 10492
rect 34054 10480 34060 10532
rect 34112 10520 34118 10532
rect 34992 10520 35020 10551
rect 34112 10492 35020 10520
rect 34112 10480 34118 10492
rect 17696 10424 20300 10452
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 20404 10424 20449 10452
rect 20404 10412 20410 10424
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 22278 10452 22284 10464
rect 20772 10424 22284 10452
rect 20772 10412 20778 10424
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 27154 10452 27160 10464
rect 24820 10424 27160 10452
rect 24820 10412 24826 10424
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 27341 10455 27399 10461
rect 27341 10421 27353 10455
rect 27387 10452 27399 10455
rect 28718 10452 28724 10464
rect 27387 10424 28724 10452
rect 27387 10421 27399 10424
rect 27341 10415 27399 10421
rect 28718 10412 28724 10424
rect 28776 10412 28782 10464
rect 33505 10455 33563 10461
rect 33505 10421 33517 10455
rect 33551 10452 33563 10455
rect 35268 10452 35296 10628
rect 35526 10616 35532 10628
rect 35584 10616 35590 10668
rect 35618 10616 35624 10668
rect 35676 10656 35682 10668
rect 35989 10659 36047 10665
rect 35989 10656 36001 10659
rect 35676 10628 36001 10656
rect 35676 10616 35682 10628
rect 35989 10625 36001 10628
rect 36035 10625 36047 10659
rect 36262 10656 36268 10668
rect 36223 10628 36268 10656
rect 35989 10619 36047 10625
rect 36262 10616 36268 10628
rect 36320 10616 36326 10668
rect 38654 10656 38660 10668
rect 36372 10628 37688 10656
rect 38615 10628 38660 10656
rect 35345 10591 35403 10597
rect 35345 10557 35357 10591
rect 35391 10588 35403 10591
rect 35802 10588 35808 10600
rect 35391 10560 35808 10588
rect 35391 10557 35403 10560
rect 35345 10551 35403 10557
rect 35802 10548 35808 10560
rect 35860 10548 35866 10600
rect 35894 10548 35900 10600
rect 35952 10588 35958 10600
rect 36081 10591 36139 10597
rect 36081 10588 36093 10591
rect 35952 10560 36093 10588
rect 35952 10548 35958 10560
rect 36081 10557 36093 10560
rect 36127 10557 36139 10591
rect 36081 10551 36139 10557
rect 36170 10548 36176 10600
rect 36228 10588 36234 10600
rect 36372 10588 36400 10628
rect 37366 10588 37372 10600
rect 36228 10560 36400 10588
rect 36455 10560 37372 10588
rect 36228 10548 36234 10560
rect 35618 10480 35624 10532
rect 35676 10480 35682 10532
rect 35713 10523 35771 10529
rect 35713 10489 35725 10523
rect 35759 10520 35771 10523
rect 36455 10520 36483 10560
rect 37366 10548 37372 10560
rect 37424 10548 37430 10600
rect 35759 10492 36483 10520
rect 35759 10489 35771 10492
rect 35713 10483 35771 10489
rect 33551 10424 35296 10452
rect 35636 10452 35664 10480
rect 35802 10452 35808 10464
rect 35636 10424 35808 10452
rect 33551 10421 33563 10424
rect 33505 10415 33563 10421
rect 35802 10412 35808 10424
rect 35860 10412 35866 10464
rect 36280 10461 36308 10492
rect 36906 10480 36912 10532
rect 36964 10520 36970 10532
rect 37660 10520 37688 10628
rect 38654 10616 38660 10628
rect 38712 10616 38718 10668
rect 38746 10616 38752 10668
rect 38804 10656 38810 10668
rect 39500 10665 39528 10696
rect 39776 10696 41414 10724
rect 38841 10659 38899 10665
rect 38841 10656 38853 10659
rect 38804 10628 38853 10656
rect 38804 10616 38810 10628
rect 38841 10625 38853 10628
rect 38887 10625 38899 10659
rect 38841 10619 38899 10625
rect 39485 10659 39543 10665
rect 39485 10625 39497 10659
rect 39531 10625 39543 10659
rect 39485 10619 39543 10625
rect 39574 10616 39580 10668
rect 39632 10656 39638 10668
rect 39669 10659 39727 10665
rect 39669 10656 39681 10659
rect 39632 10628 39681 10656
rect 39632 10616 39638 10628
rect 39669 10625 39681 10628
rect 39715 10625 39727 10659
rect 39669 10619 39727 10625
rect 37918 10588 37924 10600
rect 37879 10560 37924 10588
rect 37918 10548 37924 10560
rect 37976 10548 37982 10600
rect 38105 10591 38163 10597
rect 38105 10557 38117 10591
rect 38151 10588 38163 10591
rect 39776 10588 39804 10696
rect 40586 10656 40592 10668
rect 40547 10628 40592 10656
rect 40586 10616 40592 10628
rect 40644 10616 40650 10668
rect 40681 10659 40739 10665
rect 40681 10625 40693 10659
rect 40727 10625 40739 10659
rect 40862 10656 40868 10668
rect 40823 10628 40868 10656
rect 40681 10619 40739 10625
rect 38151 10560 39804 10588
rect 38151 10557 38163 10560
rect 38105 10551 38163 10557
rect 38930 10520 38936 10532
rect 36964 10492 37596 10520
rect 37660 10492 38936 10520
rect 36964 10480 36970 10492
rect 36265 10455 36323 10461
rect 36265 10421 36277 10455
rect 36311 10421 36323 10455
rect 36446 10452 36452 10464
rect 36407 10424 36452 10452
rect 36265 10415 36323 10421
rect 36446 10412 36452 10424
rect 36504 10412 36510 10464
rect 37366 10412 37372 10464
rect 37424 10452 37430 10464
rect 37461 10455 37519 10461
rect 37461 10452 37473 10455
rect 37424 10424 37473 10452
rect 37424 10412 37430 10424
rect 37461 10421 37473 10424
rect 37507 10421 37519 10455
rect 37568 10452 37596 10492
rect 38930 10480 38936 10492
rect 38988 10480 38994 10532
rect 40696 10520 40724 10619
rect 40862 10616 40868 10628
rect 40920 10616 40926 10668
rect 40954 10616 40960 10668
rect 41012 10656 41018 10668
rect 41386 10656 41414 10696
rect 41509 10693 41521 10727
rect 41555 10724 41567 10727
rect 41598 10724 41604 10736
rect 41555 10696 41604 10724
rect 41555 10693 41567 10696
rect 41509 10687 41567 10693
rect 41598 10684 41604 10696
rect 41656 10684 41662 10736
rect 43073 10727 43131 10733
rect 43073 10693 43085 10727
rect 43119 10724 43131 10727
rect 43254 10724 43260 10736
rect 43119 10696 43260 10724
rect 43119 10693 43131 10696
rect 43073 10687 43131 10693
rect 43254 10684 43260 10696
rect 43312 10684 43318 10736
rect 43438 10684 43444 10736
rect 43496 10724 43502 10736
rect 44177 10727 44235 10733
rect 44177 10724 44189 10727
rect 43496 10696 44189 10724
rect 43496 10684 43502 10696
rect 44177 10693 44189 10696
rect 44223 10724 44235 10727
rect 47210 10724 47216 10736
rect 44223 10696 47216 10724
rect 44223 10693 44235 10696
rect 44177 10687 44235 10693
rect 47210 10684 47216 10696
rect 47268 10724 47274 10736
rect 49421 10727 49479 10733
rect 49421 10724 49433 10727
rect 47268 10696 49433 10724
rect 47268 10684 47274 10696
rect 49421 10693 49433 10696
rect 49467 10693 49479 10727
rect 49421 10687 49479 10693
rect 49510 10684 49516 10736
rect 49568 10724 49574 10736
rect 53282 10724 53288 10736
rect 49568 10696 53288 10724
rect 49568 10684 49574 10696
rect 53282 10684 53288 10696
rect 53340 10684 53346 10736
rect 42794 10656 42800 10668
rect 41012 10628 41057 10656
rect 41386 10628 42800 10656
rect 41012 10616 41018 10628
rect 42794 10616 42800 10628
rect 42852 10616 42858 10668
rect 42981 10659 43039 10665
rect 42981 10625 42993 10659
rect 43027 10656 43039 10659
rect 57238 10656 57244 10668
rect 43027 10628 51074 10656
rect 57199 10628 57244 10656
rect 43027 10625 43039 10628
rect 42981 10619 43039 10625
rect 43257 10591 43315 10597
rect 43257 10557 43269 10591
rect 43303 10588 43315 10591
rect 43346 10588 43352 10600
rect 43303 10560 43352 10588
rect 43303 10557 43315 10560
rect 43257 10551 43315 10557
rect 43346 10548 43352 10560
rect 43404 10548 43410 10600
rect 51046 10588 51074 10628
rect 57238 10616 57244 10628
rect 57296 10616 57302 10668
rect 57425 10659 57483 10665
rect 57425 10625 57437 10659
rect 57471 10656 57483 10659
rect 57514 10656 57520 10668
rect 57471 10628 57520 10656
rect 57471 10625 57483 10628
rect 57425 10619 57483 10625
rect 57514 10616 57520 10628
rect 57572 10616 57578 10668
rect 51994 10588 52000 10600
rect 51046 10560 52000 10588
rect 51994 10548 52000 10560
rect 52052 10548 52058 10600
rect 40696 10492 46244 10520
rect 39485 10455 39543 10461
rect 39485 10452 39497 10455
rect 37568 10424 39497 10452
rect 37461 10415 37519 10421
rect 39485 10421 39497 10424
rect 39531 10421 39543 10455
rect 39485 10415 39543 10421
rect 40310 10412 40316 10464
rect 40368 10452 40374 10464
rect 40405 10455 40463 10461
rect 40405 10452 40417 10455
rect 40368 10424 40417 10452
rect 40368 10412 40374 10424
rect 40405 10421 40417 10424
rect 40451 10452 40463 10455
rect 40494 10452 40500 10464
rect 40451 10424 40500 10452
rect 40451 10421 40463 10424
rect 40405 10415 40463 10421
rect 40494 10412 40500 10424
rect 40552 10412 40558 10464
rect 40770 10412 40776 10464
rect 40828 10452 40834 10464
rect 41322 10452 41328 10464
rect 40828 10424 41328 10452
rect 40828 10412 40834 10424
rect 41322 10412 41328 10424
rect 41380 10412 41386 10464
rect 41782 10452 41788 10464
rect 41743 10424 41788 10452
rect 41782 10412 41788 10424
rect 41840 10452 41846 10464
rect 42058 10452 42064 10464
rect 41840 10424 42064 10452
rect 41840 10412 41846 10424
rect 42058 10412 42064 10424
rect 42116 10412 42122 10464
rect 42613 10455 42671 10461
rect 42613 10421 42625 10455
rect 42659 10452 42671 10455
rect 42886 10452 42892 10464
rect 42659 10424 42892 10452
rect 42659 10421 42671 10424
rect 42613 10415 42671 10421
rect 42886 10412 42892 10424
rect 42944 10412 42950 10464
rect 45462 10452 45468 10464
rect 45423 10424 45468 10452
rect 45462 10412 45468 10424
rect 45520 10412 45526 10464
rect 46216 10452 46244 10492
rect 46290 10480 46296 10532
rect 46348 10520 46354 10532
rect 58250 10520 58256 10532
rect 46348 10492 58256 10520
rect 46348 10480 46354 10492
rect 58250 10480 58256 10492
rect 58308 10480 58314 10532
rect 51718 10452 51724 10464
rect 46216 10424 51724 10452
rect 51718 10412 51724 10424
rect 51776 10412 51782 10464
rect 57330 10452 57336 10464
rect 57291 10424 57336 10452
rect 57330 10412 57336 10424
rect 57388 10412 57394 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 7558 10248 7564 10260
rect 2004 10220 7564 10248
rect 2004 10208 2010 10220
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 11793 10251 11851 10257
rect 11793 10217 11805 10251
rect 11839 10248 11851 10251
rect 11882 10248 11888 10260
rect 11839 10220 11888 10248
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 16022 10248 16028 10260
rect 14507 10220 16028 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 24026 10248 24032 10260
rect 16172 10220 24032 10248
rect 16172 10208 16178 10220
rect 24026 10208 24032 10220
rect 24084 10248 24090 10260
rect 24394 10248 24400 10260
rect 24084 10220 24400 10248
rect 24084 10208 24090 10220
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 24670 10248 24676 10260
rect 24631 10220 24676 10248
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 24946 10208 24952 10260
rect 25004 10248 25010 10260
rect 25314 10248 25320 10260
rect 25004 10220 25320 10248
rect 25004 10208 25010 10220
rect 25314 10208 25320 10220
rect 25372 10248 25378 10260
rect 25498 10248 25504 10260
rect 25372 10220 25504 10248
rect 25372 10208 25378 10220
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 28997 10251 29055 10257
rect 28997 10248 29009 10251
rect 25608 10220 29009 10248
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 11609 10183 11667 10189
rect 11609 10180 11621 10183
rect 7708 10152 11621 10180
rect 7708 10140 7714 10152
rect 11609 10149 11621 10152
rect 11655 10149 11667 10183
rect 11609 10143 11667 10149
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 14734 10180 14740 10192
rect 12400 10152 14740 10180
rect 12400 10140 12406 10152
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 20346 10180 20352 10192
rect 15304 10152 20352 10180
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11790 10112 11796 10124
rect 11379 10084 11796 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 12584 10084 15117 10112
rect 12584 10072 12590 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13872 10016 14473 10044
rect 13872 10004 13878 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14642 10044 14648 10056
rect 14603 10016 14648 10044
rect 14461 10007 14519 10013
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 15304 10053 15332 10152
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 20806 10140 20812 10192
rect 20864 10180 20870 10192
rect 25608 10180 25636 10220
rect 28997 10217 29009 10220
rect 29043 10248 29055 10251
rect 34057 10251 34115 10257
rect 34057 10248 34069 10251
rect 29043 10220 30236 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 20864 10152 25636 10180
rect 20864 10140 20870 10152
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 17681 10115 17739 10121
rect 17083 10084 17448 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 16114 10044 16120 10056
rect 16075 10016 16120 10044
rect 15289 10007 15347 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 16229 10047 16287 10053
rect 16229 10013 16241 10047
rect 16275 10044 16287 10047
rect 16942 10044 16948 10056
rect 16275 10016 16804 10044
rect 16903 10016 16948 10044
rect 16275 10013 16287 10016
rect 16229 10007 16287 10013
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 15933 9979 15991 9985
rect 15933 9976 15945 9979
rect 13780 9948 15945 9976
rect 13780 9936 13786 9948
rect 15933 9945 15945 9948
rect 15979 9945 15991 9979
rect 15933 9939 15991 9945
rect 16022 9936 16028 9988
rect 16080 9976 16086 9988
rect 16319 9979 16377 9985
rect 16319 9976 16331 9979
rect 16080 9948 16331 9976
rect 16080 9936 16086 9948
rect 16319 9945 16331 9948
rect 16365 9945 16377 9979
rect 16482 9976 16488 9988
rect 16443 9948 16488 9976
rect 16319 9939 16377 9945
rect 16482 9936 16488 9948
rect 16540 9936 16546 9988
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 16666 9908 16672 9920
rect 14148 9880 16672 9908
rect 14148 9868 14154 9880
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 16776 9908 16804 10016
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17218 10044 17224 10056
rect 17179 10016 17224 10044
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 17420 10044 17448 10084
rect 17681 10081 17693 10115
rect 17727 10112 17739 10115
rect 17770 10112 17776 10124
rect 17727 10084 17776 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18233 10115 18291 10121
rect 17920 10084 18106 10112
rect 17920 10072 17926 10084
rect 17420 10016 17724 10044
rect 17696 9988 17724 10016
rect 18078 10038 18106 10084
rect 18233 10081 18245 10115
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 18141 10047 18199 10053
rect 18141 10038 18153 10047
rect 18078 10013 18153 10038
rect 18187 10013 18199 10047
rect 18078 10010 18199 10013
rect 18141 10007 18199 10010
rect 17678 9936 17684 9988
rect 17736 9976 17742 9988
rect 18248 9976 18276 10075
rect 18506 10072 18512 10124
rect 18564 10112 18570 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18564 10084 18613 10112
rect 18564 10072 18570 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18690 10072 18696 10124
rect 18748 10112 18754 10124
rect 20714 10112 20720 10124
rect 18748 10084 20720 10112
rect 18748 10072 18754 10084
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21542 10112 21548 10124
rect 20916 10084 21548 10112
rect 20916 10056 20944 10084
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 21910 10072 21916 10124
rect 21968 10112 21974 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 21968 10084 23213 10112
rect 21968 10072 21974 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23201 10075 23259 10081
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23753 10115 23811 10121
rect 23753 10112 23765 10115
rect 23440 10084 23765 10112
rect 23440 10072 23446 10084
rect 23753 10081 23765 10084
rect 23799 10112 23811 10115
rect 24670 10112 24676 10124
rect 23799 10084 24676 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 25130 10112 25136 10124
rect 25043 10084 25136 10112
rect 25130 10072 25136 10084
rect 25188 10112 25194 10124
rect 25777 10115 25835 10121
rect 25777 10112 25789 10115
rect 25188 10084 25789 10112
rect 25188 10072 25194 10084
rect 25777 10081 25789 10084
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 28626 10072 28632 10124
rect 28684 10112 28690 10124
rect 30208 10121 30236 10220
rect 33888 10220 34069 10248
rect 33134 10140 33140 10192
rect 33192 10180 33198 10192
rect 33888 10180 33916 10220
rect 34057 10217 34069 10220
rect 34103 10217 34115 10251
rect 34057 10211 34115 10217
rect 35437 10251 35495 10257
rect 35437 10217 35449 10251
rect 35483 10248 35495 10251
rect 35802 10248 35808 10260
rect 35483 10220 35808 10248
rect 35483 10217 35495 10220
rect 35437 10211 35495 10217
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 49510 10248 49516 10260
rect 36004 10220 49516 10248
rect 33192 10152 33916 10180
rect 33192 10140 33198 10152
rect 34330 10140 34336 10192
rect 34388 10180 34394 10192
rect 35894 10180 35900 10192
rect 34388 10152 35900 10180
rect 34388 10140 34394 10152
rect 35894 10140 35900 10152
rect 35952 10140 35958 10192
rect 30193 10115 30251 10121
rect 28684 10084 30144 10112
rect 28684 10072 28690 10084
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18417 10047 18475 10053
rect 18417 10044 18429 10047
rect 18380 10016 18429 10044
rect 18380 10004 18386 10016
rect 18417 10013 18429 10016
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 19518 10004 19524 10056
rect 19576 10004 19582 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19794 10004 19800 10056
rect 19852 10053 19858 10056
rect 19852 10047 19914 10053
rect 19852 10013 19868 10047
rect 19902 10046 19914 10047
rect 19981 10047 20039 10053
rect 19902 10016 19932 10046
rect 19902 10013 19914 10016
rect 19852 10007 19914 10013
rect 19981 10013 19993 10047
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10046 20131 10047
rect 20119 10044 20199 10046
rect 20530 10044 20536 10056
rect 20119 10018 20536 10044
rect 20119 10013 20131 10018
rect 20171 10016 20536 10018
rect 20073 10007 20131 10013
rect 19852 10004 19858 10007
rect 19536 9976 19564 10004
rect 17736 9948 18276 9976
rect 19352 9948 19564 9976
rect 19996 9976 20024 10007
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 20898 10044 20904 10056
rect 20855 10016 20904 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 21177 10047 21235 10053
rect 21177 10013 21189 10047
rect 21223 10013 21235 10047
rect 21177 10007 21235 10013
rect 20438 9976 20444 9988
rect 19996 9948 20444 9976
rect 17736 9936 17742 9948
rect 19352 9908 19380 9948
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 21192 9976 21220 10007
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 21324 10016 21373 10044
rect 21324 10004 21330 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 22152 10016 22197 10044
rect 22152 10004 22158 10016
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23290 10044 23296 10056
rect 23164 10016 23296 10044
rect 23164 10004 23170 10016
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 23658 10044 23664 10056
rect 23619 10016 23664 10044
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 27617 10047 27675 10053
rect 27617 10044 27629 10047
rect 25372 10016 27629 10044
rect 25372 10004 25378 10016
rect 27617 10013 27629 10016
rect 27663 10013 27675 10047
rect 28994 10044 29000 10056
rect 27617 10007 27675 10013
rect 27816 10016 29000 10044
rect 21192 9948 21404 9976
rect 21376 9920 21404 9948
rect 22278 9936 22284 9988
rect 22336 9976 22342 9988
rect 22649 9979 22707 9985
rect 22649 9976 22661 9979
rect 22336 9948 22661 9976
rect 22336 9936 22342 9948
rect 22649 9945 22661 9948
rect 22695 9976 22707 9979
rect 23750 9976 23756 9988
rect 22695 9948 23756 9976
rect 22695 9945 22707 9948
rect 22649 9939 22707 9945
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 25225 9979 25283 9985
rect 25225 9945 25237 9979
rect 25271 9945 25283 9979
rect 25225 9939 25283 9945
rect 26044 9979 26102 9985
rect 26044 9945 26056 9979
rect 26090 9976 26102 9979
rect 27816 9976 27844 10016
rect 28994 10004 29000 10016
rect 29052 10004 29058 10056
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 30116 10053 30144 10084
rect 30193 10081 30205 10115
rect 30239 10081 30251 10115
rect 30193 10075 30251 10081
rect 30282 10072 30288 10124
rect 30340 10112 30346 10124
rect 30340 10084 30385 10112
rect 30340 10072 30346 10084
rect 31202 10072 31208 10124
rect 31260 10112 31266 10124
rect 31846 10112 31852 10124
rect 31260 10084 31852 10112
rect 31260 10072 31266 10084
rect 31312 10053 31340 10084
rect 31846 10072 31852 10084
rect 31904 10072 31910 10124
rect 32398 10072 32404 10124
rect 32456 10112 32462 10124
rect 32766 10112 32772 10124
rect 32456 10084 32772 10112
rect 32456 10072 32462 10084
rect 32766 10072 32772 10084
rect 32824 10072 32830 10124
rect 33042 10072 33048 10124
rect 33100 10112 33106 10124
rect 33100 10084 34652 10112
rect 33100 10072 33106 10084
rect 30101 10047 30159 10053
rect 29144 10016 29868 10044
rect 29144 10004 29150 10016
rect 26090 9948 27844 9976
rect 27884 9979 27942 9985
rect 26090 9945 26102 9948
rect 26044 9939 26102 9945
rect 27884 9945 27896 9979
rect 27930 9976 27942 9979
rect 29840 9976 29868 10016
rect 30101 10013 30113 10047
rect 30147 10013 30159 10047
rect 30101 10007 30159 10013
rect 31297 10047 31355 10053
rect 31297 10013 31309 10047
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 33962 10004 33968 10056
rect 34020 10044 34026 10056
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 34020 10016 34069 10044
rect 34020 10004 34026 10016
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34333 10047 34391 10053
rect 34333 10041 34345 10047
rect 34057 10007 34115 10013
rect 34256 10013 34345 10041
rect 34379 10041 34391 10047
rect 34514 10044 34520 10056
rect 34440 10041 34520 10044
rect 34379 10016 34520 10041
rect 34379 10013 34468 10016
rect 27930 9948 29776 9976
rect 29840 9948 32536 9976
rect 27930 9945 27942 9948
rect 27884 9939 27942 9945
rect 16776 9880 19380 9908
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19521 9911 19579 9917
rect 19521 9908 19533 9911
rect 19484 9880 19533 9908
rect 19484 9868 19490 9880
rect 19521 9877 19533 9880
rect 19567 9877 19579 9911
rect 19521 9871 19579 9877
rect 20625 9911 20683 9917
rect 20625 9877 20637 9911
rect 20671 9908 20683 9911
rect 20990 9908 20996 9920
rect 20671 9880 20996 9908
rect 20671 9877 20683 9880
rect 20625 9871 20683 9877
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 21082 9868 21088 9920
rect 21140 9908 21146 9920
rect 21266 9908 21272 9920
rect 21140 9880 21272 9908
rect 21140 9868 21146 9880
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21358 9868 21364 9920
rect 21416 9868 21422 9920
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 24946 9908 24952 9920
rect 22244 9880 24952 9908
rect 22244 9868 22250 9880
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 25133 9911 25191 9917
rect 25133 9908 25145 9911
rect 25096 9880 25145 9908
rect 25096 9868 25102 9880
rect 25133 9877 25145 9880
rect 25179 9877 25191 9911
rect 25240 9908 25268 9939
rect 27157 9911 27215 9917
rect 27157 9908 27169 9911
rect 25240 9880 27169 9908
rect 25133 9871 25191 9877
rect 27157 9877 27169 9880
rect 27203 9908 27215 9911
rect 27614 9908 27620 9920
rect 27203 9880 27620 9908
rect 27203 9877 27215 9880
rect 27157 9871 27215 9877
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 29748 9917 29776 9948
rect 32508 9917 32536 9948
rect 33778 9936 33784 9988
rect 33836 9976 33842 9988
rect 34256 9976 34284 10013
rect 34333 10007 34391 10013
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 33836 9948 34284 9976
rect 34624 9976 34652 10084
rect 34790 10072 34796 10124
rect 34848 10112 34854 10124
rect 34848 10084 35204 10112
rect 34848 10072 34854 10084
rect 34882 10044 34888 10056
rect 34843 10016 34888 10044
rect 34882 10004 34888 10016
rect 34940 10004 34946 10056
rect 35066 10044 35072 10056
rect 35027 10016 35072 10044
rect 35066 10004 35072 10016
rect 35124 10004 35130 10056
rect 35176 10053 35204 10084
rect 35161 10047 35219 10053
rect 35161 10013 35173 10047
rect 35207 10013 35219 10047
rect 35161 10007 35219 10013
rect 35250 10004 35256 10056
rect 35308 10044 35314 10056
rect 36004 10053 36032 10220
rect 49510 10208 49516 10220
rect 49568 10208 49574 10260
rect 57514 10208 57520 10260
rect 57572 10248 57578 10260
rect 58253 10251 58311 10257
rect 58253 10248 58265 10251
rect 57572 10220 58265 10248
rect 57572 10208 57578 10220
rect 58253 10217 58265 10220
rect 58299 10217 58311 10251
rect 58253 10211 58311 10217
rect 36262 10140 36268 10192
rect 36320 10180 36326 10192
rect 36541 10183 36599 10189
rect 36541 10180 36553 10183
rect 36320 10152 36553 10180
rect 36320 10140 36326 10152
rect 36541 10149 36553 10152
rect 36587 10149 36599 10183
rect 36541 10143 36599 10149
rect 38102 10140 38108 10192
rect 38160 10180 38166 10192
rect 39206 10180 39212 10192
rect 38160 10152 39212 10180
rect 38160 10140 38166 10152
rect 39206 10140 39212 10152
rect 39264 10140 39270 10192
rect 40402 10140 40408 10192
rect 40460 10140 40466 10192
rect 36630 10112 36636 10124
rect 36280 10084 36636 10112
rect 35989 10047 36047 10053
rect 35308 10016 35353 10044
rect 35308 10004 35314 10016
rect 35989 10013 36001 10047
rect 36035 10013 36047 10047
rect 36170 10044 36176 10056
rect 36131 10016 36176 10044
rect 35989 10007 36047 10013
rect 36170 10004 36176 10016
rect 36228 10004 36234 10056
rect 36280 10053 36308 10084
rect 36630 10072 36636 10084
rect 36688 10072 36694 10124
rect 40420 10112 40448 10140
rect 41417 10115 41475 10121
rect 39960 10084 40448 10112
rect 40512 10084 41184 10112
rect 39960 10056 39988 10084
rect 36265 10047 36323 10053
rect 36265 10013 36277 10047
rect 36311 10013 36323 10047
rect 36265 10007 36323 10013
rect 36357 10047 36415 10053
rect 36357 10013 36369 10047
rect 36403 10013 36415 10047
rect 37090 10044 37096 10056
rect 37051 10016 37096 10044
rect 36357 10007 36415 10013
rect 36372 9976 36400 10007
rect 37090 10004 37096 10016
rect 37148 10004 37154 10056
rect 37366 10053 37372 10056
rect 37360 10044 37372 10053
rect 37327 10016 37372 10044
rect 37360 10007 37372 10016
rect 37366 10004 37372 10007
rect 37424 10004 37430 10056
rect 38654 10004 38660 10056
rect 38712 10044 38718 10056
rect 39942 10044 39948 10056
rect 38712 10016 39948 10044
rect 38712 10004 38718 10016
rect 39942 10004 39948 10016
rect 40000 10004 40006 10056
rect 40034 10004 40040 10056
rect 40092 10044 40098 10056
rect 40512 10053 40540 10084
rect 40313 10047 40371 10053
rect 40313 10044 40325 10047
rect 40092 10016 40325 10044
rect 40092 10004 40098 10016
rect 40313 10013 40325 10016
rect 40359 10013 40371 10047
rect 40313 10007 40371 10013
rect 40461 10047 40540 10053
rect 40461 10013 40473 10047
rect 40507 10016 40540 10047
rect 40678 10044 40684 10056
rect 40639 10016 40684 10044
rect 40507 10013 40519 10016
rect 40461 10007 40519 10013
rect 40678 10004 40684 10016
rect 40736 10004 40742 10056
rect 40770 10004 40776 10056
rect 40828 10053 40834 10056
rect 40828 10044 40836 10053
rect 40828 10016 40873 10044
rect 40828 10007 40836 10016
rect 40828 10004 40834 10007
rect 34624 9948 36400 9976
rect 33836 9936 33842 9948
rect 36446 9936 36452 9988
rect 36504 9976 36510 9988
rect 38933 9979 38991 9985
rect 38933 9976 38945 9979
rect 36504 9948 38945 9976
rect 36504 9936 36510 9948
rect 38933 9945 38945 9948
rect 38979 9945 38991 9979
rect 39114 9976 39120 9988
rect 39075 9948 39120 9976
rect 38933 9939 38991 9945
rect 39114 9936 39120 9948
rect 39172 9936 39178 9988
rect 39206 9936 39212 9988
rect 39264 9976 39270 9988
rect 39301 9979 39359 9985
rect 39301 9976 39313 9979
rect 39264 9948 39313 9976
rect 39264 9936 39270 9948
rect 39301 9945 39313 9948
rect 39347 9945 39359 9979
rect 39301 9939 39359 9945
rect 40589 9979 40647 9985
rect 40589 9945 40601 9979
rect 40635 9976 40647 9979
rect 41046 9976 41052 9988
rect 40635 9948 41052 9976
rect 40635 9945 40647 9948
rect 40589 9939 40647 9945
rect 29733 9911 29791 9917
rect 29733 9877 29745 9911
rect 29779 9877 29791 9911
rect 29733 9871 29791 9877
rect 32493 9911 32551 9917
rect 32493 9877 32505 9911
rect 32539 9877 32551 9911
rect 32493 9871 32551 9877
rect 32674 9868 32680 9920
rect 32732 9908 32738 9920
rect 34241 9911 34299 9917
rect 34241 9908 34253 9911
rect 32732 9880 34253 9908
rect 32732 9868 32738 9880
rect 34241 9877 34253 9880
rect 34287 9877 34299 9911
rect 34241 9871 34299 9877
rect 34790 9868 34796 9920
rect 34848 9908 34854 9920
rect 37918 9908 37924 9920
rect 34848 9880 37924 9908
rect 34848 9868 34854 9880
rect 37918 9868 37924 9880
rect 37976 9908 37982 9920
rect 38473 9911 38531 9917
rect 38473 9908 38485 9911
rect 37976 9880 38485 9908
rect 37976 9868 37982 9880
rect 38473 9877 38485 9880
rect 38519 9877 38531 9911
rect 38473 9871 38531 9877
rect 38654 9868 38660 9920
rect 38712 9908 38718 9920
rect 40604 9908 40632 9939
rect 41046 9936 41052 9948
rect 41104 9936 41110 9988
rect 41156 9976 41184 10084
rect 41417 10081 41429 10115
rect 41463 10112 41475 10115
rect 42702 10112 42708 10124
rect 41463 10084 42708 10112
rect 41463 10081 41475 10084
rect 41417 10075 41475 10081
rect 42702 10072 42708 10084
rect 42760 10072 42766 10124
rect 43073 10115 43131 10121
rect 43073 10081 43085 10115
rect 43119 10112 43131 10115
rect 43162 10112 43168 10124
rect 43119 10084 43168 10112
rect 43119 10081 43131 10084
rect 43073 10075 43131 10081
rect 43162 10072 43168 10084
rect 43220 10072 43226 10124
rect 43346 10072 43352 10124
rect 43404 10112 43410 10124
rect 44177 10115 44235 10121
rect 44177 10112 44189 10115
rect 43404 10084 44189 10112
rect 43404 10072 43410 10084
rect 44177 10081 44189 10084
rect 44223 10081 44235 10115
rect 56870 10112 56876 10124
rect 56831 10084 56876 10112
rect 44177 10075 44235 10081
rect 56870 10072 56876 10084
rect 56928 10072 56934 10124
rect 41693 10047 41751 10053
rect 41693 10013 41705 10047
rect 41739 10044 41751 10047
rect 43622 10044 43628 10056
rect 41739 10016 43628 10044
rect 41739 10013 41751 10016
rect 41693 10007 41751 10013
rect 43622 10004 43628 10016
rect 43680 10004 43686 10056
rect 43901 10047 43959 10053
rect 43901 10013 43913 10047
rect 43947 10013 43959 10047
rect 43901 10007 43959 10013
rect 41156 9948 41552 9976
rect 38712 9880 40632 9908
rect 40957 9911 41015 9917
rect 38712 9868 38718 9880
rect 40957 9877 40969 9911
rect 41003 9908 41015 9911
rect 41414 9908 41420 9920
rect 41003 9880 41420 9908
rect 41003 9877 41015 9880
rect 40957 9871 41015 9877
rect 41414 9868 41420 9880
rect 41472 9868 41478 9920
rect 41524 9908 41552 9948
rect 42794 9936 42800 9988
rect 42852 9976 42858 9988
rect 43916 9976 43944 10007
rect 45094 9976 45100 9988
rect 42852 9948 45100 9976
rect 42852 9936 42858 9948
rect 45094 9936 45100 9948
rect 45152 9936 45158 9988
rect 56778 9936 56784 9988
rect 56836 9976 56842 9988
rect 57118 9979 57176 9985
rect 57118 9976 57130 9979
rect 56836 9948 57130 9976
rect 56836 9936 56842 9948
rect 57118 9945 57130 9948
rect 57164 9945 57176 9979
rect 57118 9939 57176 9945
rect 45186 9908 45192 9920
rect 41524 9880 45192 9908
rect 45186 9868 45192 9880
rect 45244 9868 45250 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 17770 9704 17776 9716
rect 17000 9676 17776 9704
rect 17000 9664 17006 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 22554 9704 22560 9716
rect 18708 9676 22560 9704
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 17218 9636 17224 9648
rect 14424 9608 15240 9636
rect 14424 9596 14430 9608
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11974 9568 11980 9580
rect 11747 9540 11980 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 14550 9568 14556 9580
rect 14511 9540 14556 9568
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15212 9577 15240 9608
rect 15764 9608 17224 9636
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 12158 9500 12164 9512
rect 12119 9472 12164 9500
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 15764 9500 15792 9608
rect 17218 9596 17224 9608
rect 17276 9636 17282 9648
rect 17276 9608 17908 9636
rect 17276 9596 17282 9608
rect 16390 9528 16396 9580
rect 16448 9528 16454 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17126 9568 17132 9580
rect 16899 9540 17132 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17770 9568 17776 9580
rect 17731 9540 17776 9568
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17880 9577 17908 9608
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 14691 9472 15792 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16298 9500 16304 9512
rect 15896 9472 15941 9500
rect 16259 9472 16304 9500
rect 15896 9460 15902 9472
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16408 9500 16436 9528
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16408 9472 16957 9500
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 18064 9500 18092 9531
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18708 9577 18736 9676
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 24397 9707 24455 9713
rect 24397 9673 24409 9707
rect 24443 9704 24455 9707
rect 24443 9676 24624 9704
rect 24443 9673 24455 9676
rect 24397 9667 24455 9673
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 19153 9639 19211 9645
rect 19153 9636 19165 9639
rect 18932 9608 19165 9636
rect 18932 9596 18938 9608
rect 19153 9605 19165 9608
rect 19199 9636 19211 9639
rect 20806 9636 20812 9648
rect 19199 9608 20812 9636
rect 19199 9605 19211 9608
rect 19153 9599 19211 9605
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 20898 9596 20904 9648
rect 20956 9636 20962 9648
rect 20993 9639 21051 9645
rect 20993 9636 21005 9639
rect 20956 9608 21005 9636
rect 20956 9596 20962 9608
rect 20993 9605 21005 9608
rect 21039 9605 21051 9639
rect 24596 9636 24624 9676
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 26602 9704 26608 9716
rect 25004 9676 26608 9704
rect 25004 9664 25010 9676
rect 26602 9664 26608 9676
rect 26660 9664 26666 9716
rect 26694 9664 26700 9716
rect 26752 9704 26758 9716
rect 28626 9704 28632 9716
rect 26752 9676 28632 9704
rect 26752 9664 26758 9676
rect 28626 9664 28632 9676
rect 28684 9664 28690 9716
rect 28994 9704 29000 9716
rect 28955 9676 29000 9704
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 29730 9664 29736 9716
rect 29788 9704 29794 9716
rect 30282 9704 30288 9716
rect 29788 9676 30288 9704
rect 29788 9664 29794 9676
rect 30282 9664 30288 9676
rect 30340 9664 30346 9716
rect 30466 9664 30472 9716
rect 30524 9704 30530 9716
rect 30561 9707 30619 9713
rect 30561 9704 30573 9707
rect 30524 9676 30573 9704
rect 30524 9664 30530 9676
rect 30561 9673 30573 9676
rect 30607 9704 30619 9707
rect 30926 9704 30932 9716
rect 30607 9676 30932 9704
rect 30607 9673 30619 9676
rect 30561 9667 30619 9673
rect 30926 9664 30932 9676
rect 30984 9704 30990 9716
rect 31573 9707 31631 9713
rect 31573 9704 31585 9707
rect 30984 9676 31585 9704
rect 30984 9664 30990 9676
rect 31573 9673 31585 9676
rect 31619 9673 31631 9707
rect 31573 9667 31631 9673
rect 32309 9707 32367 9713
rect 32309 9673 32321 9707
rect 32355 9704 32367 9707
rect 32398 9704 32404 9716
rect 32355 9676 32404 9704
rect 32355 9673 32367 9676
rect 32309 9667 32367 9673
rect 32398 9664 32404 9676
rect 32456 9664 32462 9716
rect 32674 9704 32680 9716
rect 32635 9676 32680 9704
rect 32674 9664 32680 9676
rect 32732 9664 32738 9716
rect 32950 9664 32956 9716
rect 33008 9704 33014 9716
rect 34790 9704 34796 9716
rect 33008 9676 34796 9704
rect 33008 9664 33014 9676
rect 34790 9664 34796 9676
rect 34848 9664 34854 9716
rect 34882 9664 34888 9716
rect 34940 9704 34946 9716
rect 40313 9707 40371 9713
rect 34940 9676 40264 9704
rect 34940 9664 34946 9676
rect 25038 9636 25044 9648
rect 24596 9608 25044 9636
rect 20993 9599 21051 9605
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 25133 9639 25191 9645
rect 25133 9605 25145 9639
rect 25179 9636 25191 9639
rect 25866 9636 25872 9648
rect 25179 9608 25872 9636
rect 25179 9605 25191 9608
rect 25133 9599 25191 9605
rect 25866 9596 25872 9608
rect 25924 9596 25930 9648
rect 27614 9596 27620 9648
rect 27672 9636 27678 9648
rect 29365 9639 29423 9645
rect 29365 9636 29377 9639
rect 27672 9608 29377 9636
rect 27672 9596 27678 9608
rect 29365 9605 29377 9608
rect 29411 9605 29423 9639
rect 29365 9599 29423 9605
rect 29454 9596 29460 9648
rect 29512 9636 29518 9648
rect 29512 9608 29557 9636
rect 29512 9596 29518 9608
rect 29638 9596 29644 9648
rect 29696 9636 29702 9648
rect 30745 9639 30803 9645
rect 30745 9636 30757 9639
rect 29696 9608 30757 9636
rect 29696 9596 29702 9608
rect 30745 9605 30757 9608
rect 30791 9605 30803 9639
rect 30745 9599 30803 9605
rect 31110 9596 31116 9648
rect 31168 9636 31174 9648
rect 31389 9639 31447 9645
rect 31389 9636 31401 9639
rect 31168 9608 31401 9636
rect 31168 9596 31174 9608
rect 31389 9605 31401 9608
rect 31435 9605 31447 9639
rect 33778 9636 33784 9648
rect 31389 9599 31447 9605
rect 32508 9608 33784 9636
rect 18693 9571 18751 9577
rect 18196 9540 18241 9568
rect 18196 9528 18202 9540
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19702 9568 19708 9580
rect 19024 9540 19708 9568
rect 19024 9528 19030 9540
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 19886 9568 19892 9580
rect 19847 9540 19892 9568
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9537 20315 9571
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20257 9531 20315 9537
rect 17644 9472 18092 9500
rect 17644 9460 17650 9472
rect 18322 9460 18328 9512
rect 18380 9500 18386 9512
rect 20272 9500 20300 9531
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21416 9540 21465 9568
rect 21416 9528 21422 9540
rect 21453 9537 21465 9540
rect 21499 9568 21511 9571
rect 21910 9568 21916 9580
rect 21499 9540 21916 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22186 9568 22192 9580
rect 22147 9540 22192 9568
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 23845 9571 23903 9577
rect 23845 9537 23857 9571
rect 23891 9568 23903 9571
rect 24210 9568 24216 9580
rect 23891 9540 24216 9568
rect 23891 9537 23903 9540
rect 23845 9531 23903 9537
rect 24210 9528 24216 9540
rect 24268 9528 24274 9580
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9537 24547 9571
rect 24489 9531 24547 9537
rect 24581 9571 24639 9577
rect 24581 9537 24593 9571
rect 24627 9566 24639 9571
rect 25590 9568 25596 9580
rect 24688 9566 25596 9568
rect 24627 9540 25596 9566
rect 24627 9538 24716 9540
rect 24627 9537 24639 9538
rect 24581 9531 24639 9537
rect 20898 9500 20904 9512
rect 18380 9472 20904 9500
rect 18380 9460 18386 9472
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22738 9500 22744 9512
rect 22152 9472 22744 9500
rect 22152 9460 22158 9472
rect 22738 9460 22744 9472
rect 22796 9500 22802 9512
rect 23201 9503 23259 9509
rect 23201 9500 23213 9503
rect 22796 9472 23213 9500
rect 22796 9460 22802 9472
rect 23201 9469 23213 9472
rect 23247 9500 23259 9503
rect 23382 9500 23388 9512
rect 23247 9472 23388 9500
rect 23247 9469 23259 9472
rect 23201 9463 23259 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9469 24087 9503
rect 24504 9500 24532 9531
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 25961 9571 26019 9577
rect 25961 9537 25973 9571
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 25038 9500 25044 9512
rect 24504 9472 25044 9500
rect 24029 9463 24087 9469
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 11977 9435 12035 9441
rect 11977 9432 11989 9435
rect 5868 9404 11989 9432
rect 5868 9392 5874 9404
rect 11977 9401 11989 9404
rect 12023 9401 12035 9435
rect 11977 9395 12035 9401
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 12124 9404 16129 9432
rect 12124 9392 12130 9404
rect 16117 9401 16129 9404
rect 16163 9401 16175 9435
rect 16117 9395 16175 9401
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 20714 9432 20720 9444
rect 16448 9404 20720 9432
rect 16448 9392 16454 9404
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 20806 9392 20812 9444
rect 20864 9432 20870 9444
rect 23658 9432 23664 9444
rect 20864 9404 23664 9432
rect 20864 9392 20870 9404
rect 23658 9392 23664 9404
rect 23716 9392 23722 9444
rect 24044 9432 24072 9463
rect 25038 9460 25044 9472
rect 25096 9460 25102 9512
rect 25130 9460 25136 9512
rect 25188 9500 25194 9512
rect 25792 9500 25820 9531
rect 25188 9472 25820 9500
rect 25188 9460 25194 9472
rect 25866 9460 25872 9512
rect 25924 9500 25930 9512
rect 25976 9500 26004 9531
rect 26050 9528 26056 9580
rect 26108 9568 26114 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26108 9540 27169 9568
rect 26108 9528 26114 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27430 9528 27436 9580
rect 27488 9568 27494 9580
rect 27488 9540 28488 9568
rect 27488 9528 27494 9540
rect 26418 9500 26424 9512
rect 25924 9472 26004 9500
rect 26379 9472 26424 9500
rect 25924 9460 25930 9472
rect 26418 9460 26424 9472
rect 26476 9460 26482 9512
rect 26513 9503 26571 9509
rect 26513 9469 26525 9503
rect 26559 9469 26571 9503
rect 26513 9463 26571 9469
rect 26142 9432 26148 9444
rect 24044 9404 26148 9432
rect 26142 9392 26148 9404
rect 26200 9432 26206 9444
rect 26528 9432 26556 9463
rect 26970 9460 26976 9512
rect 27028 9500 27034 9512
rect 28258 9500 28264 9512
rect 27028 9472 28264 9500
rect 27028 9460 27034 9472
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 28353 9503 28411 9509
rect 28353 9469 28365 9503
rect 28399 9469 28411 9503
rect 28353 9463 28411 9469
rect 27430 9432 27436 9444
rect 26200 9404 27436 9432
rect 26200 9392 26206 9404
rect 27430 9392 27436 9404
rect 27488 9392 27494 9444
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 14918 9364 14924 9376
rect 10928 9336 14924 9364
rect 10928 9324 10934 9336
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 16758 9364 16764 9376
rect 15335 9336 16764 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 16908 9336 17601 9364
rect 16908 9324 16914 9336
rect 17589 9333 17601 9336
rect 17635 9364 17647 9367
rect 18874 9364 18880 9376
rect 17635 9336 18880 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 19886 9364 19892 9376
rect 19024 9336 19892 9364
rect 19024 9324 19030 9336
rect 19886 9324 19892 9336
rect 19944 9364 19950 9376
rect 21358 9364 21364 9376
rect 19944 9336 21364 9364
rect 19944 9324 19950 9336
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 25130 9364 25136 9376
rect 24544 9336 25136 9364
rect 24544 9324 24550 9336
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 25774 9324 25780 9376
rect 25832 9364 25838 9376
rect 28368 9364 28396 9463
rect 28460 9432 28488 9540
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 30193 9571 30251 9577
rect 30193 9568 30205 9571
rect 29052 9540 30205 9568
rect 29052 9528 29058 9540
rect 30193 9537 30205 9540
rect 30239 9537 30251 9571
rect 30193 9531 30251 9537
rect 30282 9528 30288 9580
rect 30340 9568 30346 9580
rect 30377 9571 30435 9577
rect 30377 9568 30389 9571
rect 30340 9540 30389 9568
rect 30340 9528 30346 9540
rect 30377 9537 30389 9540
rect 30423 9537 30435 9571
rect 30377 9531 30435 9537
rect 30515 9571 30573 9577
rect 30515 9537 30527 9571
rect 30561 9568 30573 9571
rect 31018 9568 31024 9580
rect 30561 9540 31024 9568
rect 30561 9537 30573 9540
rect 30515 9531 30573 9537
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31202 9568 31208 9580
rect 31163 9540 31208 9568
rect 31202 9528 31208 9540
rect 31260 9528 31266 9580
rect 31570 9577 31576 9580
rect 31527 9571 31576 9577
rect 31527 9537 31539 9571
rect 31573 9537 31576 9571
rect 31527 9531 31576 9537
rect 31570 9528 31576 9531
rect 31628 9528 31634 9580
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 32508 9577 32536 9608
rect 33778 9596 33784 9608
rect 33836 9596 33842 9648
rect 33965 9639 34023 9645
rect 33965 9605 33977 9639
rect 34011 9636 34023 9639
rect 34238 9636 34244 9648
rect 34011 9608 34244 9636
rect 34011 9605 34023 9608
rect 33965 9599 34023 9605
rect 34238 9596 34244 9608
rect 34296 9596 34302 9648
rect 35066 9596 35072 9648
rect 35124 9636 35130 9648
rect 35897 9639 35955 9645
rect 35897 9636 35909 9639
rect 35124 9608 35909 9636
rect 35124 9596 35130 9608
rect 32493 9571 32551 9577
rect 31812 9540 31855 9568
rect 31812 9528 31818 9540
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 32766 9568 32772 9580
rect 32727 9540 32772 9568
rect 32493 9531 32551 9537
rect 32766 9528 32772 9540
rect 32824 9528 32830 9580
rect 33410 9528 33416 9580
rect 33468 9568 33474 9580
rect 33689 9571 33747 9577
rect 33689 9568 33701 9571
rect 33468 9540 33701 9568
rect 33468 9528 33474 9540
rect 33689 9537 33701 9540
rect 33735 9537 33747 9571
rect 33689 9531 33747 9537
rect 33870 9528 33876 9580
rect 33928 9568 33934 9580
rect 33928 9540 33973 9568
rect 33928 9528 33934 9540
rect 34054 9528 34060 9580
rect 34112 9568 34118 9580
rect 34112 9540 34157 9568
rect 34112 9528 34118 9540
rect 34606 9528 34612 9580
rect 34664 9568 34670 9580
rect 34793 9571 34851 9577
rect 34793 9568 34805 9571
rect 34664 9540 34805 9568
rect 34664 9528 34670 9540
rect 34793 9537 34805 9540
rect 34839 9537 34851 9571
rect 34793 9531 34851 9537
rect 34882 9528 34888 9580
rect 34940 9568 34946 9580
rect 35434 9568 35440 9580
rect 34940 9540 35440 9568
rect 34940 9528 34946 9540
rect 35434 9528 35440 9540
rect 35492 9528 35498 9580
rect 28534 9460 28540 9512
rect 28592 9500 28598 9512
rect 29549 9503 29607 9509
rect 29549 9500 29561 9503
rect 28592 9472 29561 9500
rect 28592 9460 28598 9472
rect 29549 9469 29561 9472
rect 29595 9500 29607 9503
rect 29595 9472 30420 9500
rect 29595 9469 29607 9472
rect 29549 9463 29607 9469
rect 29822 9432 29828 9444
rect 28460 9404 29828 9432
rect 29822 9392 29828 9404
rect 29880 9392 29886 9444
rect 30392 9432 30420 9472
rect 33962 9460 33968 9512
rect 34020 9500 34026 9512
rect 34330 9500 34336 9512
rect 34020 9472 34336 9500
rect 34020 9460 34026 9472
rect 34330 9460 34336 9472
rect 34388 9460 34394 9512
rect 35544 9500 35572 9608
rect 35897 9605 35909 9608
rect 35943 9605 35955 9639
rect 39298 9636 39304 9648
rect 35897 9599 35955 9605
rect 37246 9608 39304 9636
rect 35713 9571 35771 9577
rect 35713 9537 35725 9571
rect 35759 9537 35771 9571
rect 35713 9531 35771 9537
rect 35452 9472 35572 9500
rect 35728 9500 35756 9531
rect 35802 9528 35808 9580
rect 35860 9568 35866 9580
rect 35981 9571 36039 9577
rect 35981 9568 35993 9571
rect 35860 9540 35993 9568
rect 35860 9528 35866 9540
rect 35981 9537 35993 9540
rect 36027 9537 36039 9571
rect 35981 9531 36039 9537
rect 36078 9528 36084 9580
rect 36136 9568 36142 9580
rect 36538 9568 36544 9580
rect 36136 9540 36544 9568
rect 36136 9528 36142 9540
rect 36538 9528 36544 9540
rect 36596 9528 36602 9580
rect 36630 9528 36636 9580
rect 36688 9568 36694 9580
rect 36725 9571 36783 9577
rect 36725 9568 36737 9571
rect 36688 9540 36737 9568
rect 36688 9528 36694 9540
rect 36725 9537 36737 9540
rect 36771 9537 36783 9571
rect 36906 9568 36912 9580
rect 36867 9540 36912 9568
rect 36725 9531 36783 9537
rect 36906 9528 36912 9540
rect 36964 9528 36970 9580
rect 37246 9500 37274 9608
rect 39298 9596 39304 9608
rect 39356 9596 39362 9648
rect 39850 9596 39856 9648
rect 39908 9636 39914 9648
rect 40037 9639 40095 9645
rect 40037 9636 40049 9639
rect 39908 9608 40049 9636
rect 39908 9596 39914 9608
rect 40037 9605 40049 9608
rect 40083 9605 40095 9639
rect 40236 9636 40264 9676
rect 40313 9673 40325 9707
rect 40359 9704 40371 9707
rect 40954 9704 40960 9716
rect 40359 9676 40960 9704
rect 40359 9673 40371 9676
rect 40313 9667 40371 9673
rect 40954 9664 40960 9676
rect 41012 9664 41018 9716
rect 41874 9704 41880 9716
rect 41064 9676 41880 9704
rect 41064 9636 41092 9676
rect 41874 9664 41880 9676
rect 41932 9664 41938 9716
rect 43346 9664 43352 9716
rect 43404 9704 43410 9716
rect 43993 9707 44051 9713
rect 43993 9704 44005 9707
rect 43404 9676 44005 9704
rect 43404 9664 43410 9676
rect 43993 9673 44005 9676
rect 44039 9673 44051 9707
rect 43993 9667 44051 9673
rect 56965 9707 57023 9713
rect 56965 9673 56977 9707
rect 57011 9704 57023 9707
rect 57330 9704 57336 9716
rect 57011 9676 57336 9704
rect 57011 9673 57023 9676
rect 56965 9667 57023 9673
rect 57330 9664 57336 9676
rect 57388 9664 57394 9716
rect 58250 9704 58256 9716
rect 58211 9676 58256 9704
rect 58250 9664 58256 9676
rect 58308 9664 58314 9716
rect 42886 9645 42892 9648
rect 40236 9608 41092 9636
rect 40037 9599 40095 9605
rect 42880 9599 42892 9645
rect 42944 9636 42950 9648
rect 44910 9636 44916 9648
rect 42944 9608 42980 9636
rect 44871 9608 44916 9636
rect 42886 9596 42892 9599
rect 42944 9596 42950 9608
rect 44910 9596 44916 9608
rect 44968 9596 44974 9648
rect 37826 9568 37832 9580
rect 37787 9540 37832 9568
rect 37826 9528 37832 9540
rect 37884 9528 37890 9580
rect 38381 9571 38439 9577
rect 38381 9537 38393 9571
rect 38427 9568 38439 9571
rect 38654 9568 38660 9580
rect 38427 9540 38660 9568
rect 38427 9537 38439 9540
rect 38381 9531 38439 9537
rect 38654 9528 38660 9540
rect 38712 9528 38718 9580
rect 38930 9568 38936 9580
rect 38891 9540 38936 9568
rect 38930 9528 38936 9540
rect 38988 9528 38994 9580
rect 39117 9571 39175 9577
rect 39117 9537 39129 9571
rect 39163 9537 39175 9571
rect 39117 9531 39175 9537
rect 39209 9571 39267 9577
rect 39209 9537 39221 9571
rect 39255 9537 39267 9571
rect 39209 9531 39267 9537
rect 39669 9571 39727 9577
rect 39669 9537 39681 9571
rect 39715 9537 39727 9571
rect 39669 9531 39727 9537
rect 35728 9472 37274 9500
rect 35452 9444 35480 9472
rect 31294 9432 31300 9444
rect 30392 9404 31300 9432
rect 31294 9392 31300 9404
rect 31352 9392 31358 9444
rect 31570 9392 31576 9444
rect 31628 9432 31634 9444
rect 32950 9432 32956 9444
rect 31628 9404 32956 9432
rect 31628 9392 31634 9404
rect 32950 9392 32956 9404
rect 33008 9392 33014 9444
rect 33612 9404 35406 9432
rect 31938 9364 31944 9376
rect 25832 9336 31944 9364
rect 25832 9324 25838 9336
rect 31938 9324 31944 9336
rect 31996 9324 32002 9376
rect 32122 9324 32128 9376
rect 32180 9364 32186 9376
rect 33612 9364 33640 9404
rect 32180 9336 33640 9364
rect 32180 9324 32186 9336
rect 33686 9324 33692 9376
rect 33744 9364 33750 9376
rect 34241 9367 34299 9373
rect 34241 9364 34253 9367
rect 33744 9336 34253 9364
rect 33744 9324 33750 9336
rect 34241 9333 34253 9336
rect 34287 9333 34299 9367
rect 34974 9364 34980 9376
rect 34935 9336 34980 9364
rect 34241 9327 34299 9333
rect 34974 9324 34980 9336
rect 35032 9324 35038 9376
rect 35378 9364 35406 9404
rect 35434 9392 35440 9444
rect 35492 9392 35498 9444
rect 35986 9392 35992 9444
rect 36044 9432 36050 9444
rect 36725 9435 36783 9441
rect 36725 9432 36737 9435
rect 36044 9404 36737 9432
rect 36044 9392 36050 9404
rect 36725 9401 36737 9404
rect 36771 9401 36783 9435
rect 36725 9395 36783 9401
rect 35618 9364 35624 9376
rect 35378 9336 35624 9364
rect 35618 9324 35624 9336
rect 35676 9324 35682 9376
rect 35802 9324 35808 9376
rect 35860 9364 35866 9376
rect 36265 9367 36323 9373
rect 36265 9364 36277 9367
rect 35860 9336 36277 9364
rect 35860 9324 35866 9336
rect 36265 9333 36277 9336
rect 36311 9333 36323 9367
rect 36265 9327 36323 9333
rect 38654 9324 38660 9376
rect 38712 9364 38718 9376
rect 38933 9367 38991 9373
rect 38933 9364 38945 9367
rect 38712 9336 38945 9364
rect 38712 9324 38718 9336
rect 38933 9333 38945 9336
rect 38979 9333 38991 9367
rect 39132 9364 39160 9531
rect 39224 9432 39252 9531
rect 39684 9500 39712 9531
rect 39758 9528 39764 9580
rect 39816 9568 39822 9580
rect 39945 9571 40003 9577
rect 39816 9540 39861 9568
rect 39816 9528 39822 9540
rect 39945 9537 39957 9571
rect 39991 9537 40003 9571
rect 39945 9531 40003 9537
rect 40175 9571 40233 9577
rect 40175 9537 40187 9571
rect 40221 9568 40233 9571
rect 40494 9568 40500 9580
rect 40221 9540 40500 9568
rect 40221 9537 40233 9540
rect 40175 9531 40233 9537
rect 39684 9472 39804 9500
rect 39666 9432 39672 9444
rect 39224 9404 39672 9432
rect 39666 9392 39672 9404
rect 39724 9392 39730 9444
rect 39776 9432 39804 9472
rect 39850 9460 39856 9512
rect 39908 9500 39914 9512
rect 39960 9500 39988 9531
rect 40494 9528 40500 9540
rect 40552 9568 40558 9580
rect 40770 9568 40776 9580
rect 40552 9540 40776 9568
rect 40552 9528 40558 9540
rect 40770 9528 40776 9540
rect 40828 9528 40834 9580
rect 41414 9528 41420 9580
rect 41472 9568 41478 9580
rect 41785 9571 41843 9577
rect 41472 9540 41517 9568
rect 41472 9528 41478 9540
rect 41785 9537 41797 9571
rect 41831 9568 41843 9571
rect 42613 9571 42671 9577
rect 41831 9540 42564 9568
rect 41831 9537 41843 9540
rect 41785 9531 41843 9537
rect 40310 9500 40316 9512
rect 39908 9472 40316 9500
rect 39908 9460 39914 9472
rect 40310 9460 40316 9472
rect 40368 9460 40374 9512
rect 41509 9503 41567 9509
rect 41509 9469 41521 9503
rect 41555 9469 41567 9503
rect 41509 9463 41567 9469
rect 40034 9432 40040 9444
rect 39776 9404 40040 9432
rect 40034 9392 40040 9404
rect 40092 9392 40098 9444
rect 41524 9432 41552 9463
rect 41598 9460 41604 9512
rect 41656 9500 41662 9512
rect 41877 9503 41935 9509
rect 41877 9500 41889 9503
rect 41656 9472 41889 9500
rect 41656 9460 41662 9472
rect 41877 9469 41889 9472
rect 41923 9469 41935 9503
rect 41877 9463 41935 9469
rect 42242 9432 42248 9444
rect 41524 9404 42248 9432
rect 42242 9392 42248 9404
rect 42300 9392 42306 9444
rect 40770 9364 40776 9376
rect 39132 9336 40776 9364
rect 38933 9327 38991 9333
rect 40770 9324 40776 9336
rect 40828 9324 40834 9376
rect 40865 9367 40923 9373
rect 40865 9333 40877 9367
rect 40911 9364 40923 9367
rect 40954 9364 40960 9376
rect 40911 9336 40960 9364
rect 40911 9333 40923 9336
rect 40865 9327 40923 9333
rect 40954 9324 40960 9336
rect 41012 9364 41018 9376
rect 41230 9364 41236 9376
rect 41012 9336 41236 9364
rect 41012 9324 41018 9336
rect 41230 9324 41236 9336
rect 41288 9324 41294 9376
rect 42536 9364 42564 9540
rect 42613 9537 42625 9571
rect 42659 9568 42671 9571
rect 42702 9568 42708 9580
rect 42659 9540 42708 9568
rect 42659 9537 42671 9540
rect 42613 9531 42671 9537
rect 42702 9528 42708 9540
rect 42760 9528 42766 9580
rect 56686 9528 56692 9580
rect 56744 9568 56750 9580
rect 56781 9571 56839 9577
rect 56781 9568 56793 9571
rect 56744 9540 56793 9568
rect 56744 9528 56750 9540
rect 56781 9537 56793 9540
rect 56827 9537 56839 9571
rect 56781 9531 56839 9537
rect 57057 9571 57115 9577
rect 57057 9537 57069 9571
rect 57103 9537 57115 9571
rect 58066 9568 58072 9580
rect 58027 9540 58072 9568
rect 57057 9531 57115 9537
rect 43990 9460 43996 9512
rect 44048 9500 44054 9512
rect 45005 9503 45063 9509
rect 45005 9500 45017 9503
rect 44048 9472 45017 9500
rect 44048 9460 44054 9472
rect 45005 9469 45017 9472
rect 45051 9469 45063 9503
rect 45005 9463 45063 9469
rect 45094 9460 45100 9512
rect 45152 9500 45158 9512
rect 45152 9472 45197 9500
rect 45152 9460 45158 9472
rect 55398 9460 55404 9512
rect 55456 9500 55462 9512
rect 57072 9500 57100 9531
rect 58066 9528 58072 9540
rect 58124 9528 58130 9580
rect 55456 9472 57100 9500
rect 55456 9460 55462 9472
rect 44726 9432 44732 9444
rect 43916 9404 44732 9432
rect 43916 9364 43944 9404
rect 44726 9392 44732 9404
rect 44784 9392 44790 9444
rect 56778 9432 56784 9444
rect 56739 9404 56784 9432
rect 56778 9392 56784 9404
rect 56836 9392 56842 9444
rect 44542 9364 44548 9376
rect 42536 9336 43944 9364
rect 44503 9336 44548 9364
rect 44542 9324 44548 9336
rect 44600 9324 44606 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 16850 9160 16856 9172
rect 14884 9132 16856 9160
rect 14884 9120 14890 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17402 9160 17408 9172
rect 17363 9132 17408 9160
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 18966 9160 18972 9172
rect 18748 9132 18972 9160
rect 18748 9120 18754 9132
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 20073 9163 20131 9169
rect 20073 9160 20085 9163
rect 19392 9132 20085 9160
rect 19392 9120 19398 9132
rect 20073 9129 20085 9132
rect 20119 9129 20131 9163
rect 20073 9123 20131 9129
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 21600 9132 23888 9160
rect 21600 9120 21606 9132
rect 15010 9052 15016 9104
rect 15068 9092 15074 9104
rect 15838 9092 15844 9104
rect 15068 9064 15844 9092
rect 15068 9052 15074 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 16393 9095 16451 9101
rect 16393 9061 16405 9095
rect 16439 9092 16451 9095
rect 17954 9092 17960 9104
rect 16439 9064 17960 9092
rect 16439 9061 16451 9064
rect 16393 9055 16451 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 19058 9052 19064 9104
rect 19116 9092 19122 9104
rect 19116 9064 23796 9092
rect 19116 9052 19122 9064
rect 18046 9024 18052 9036
rect 15672 8996 18052 9024
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 13722 8956 13728 8968
rect 1627 8928 13728 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 15672 8965 15700 8996
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 18524 8996 18920 9024
rect 15657 8959 15715 8965
rect 15657 8925 15669 8959
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16390 8956 16396 8968
rect 16347 8928 16396 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17586 8956 17592 8968
rect 17543 8928 17592 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 16206 8888 16212 8900
rect 13740 8860 16212 8888
rect 13740 8832 13768 8860
rect 16206 8848 16212 8860
rect 16264 8888 16270 8900
rect 16500 8888 16528 8919
rect 16264 8860 16528 8888
rect 17052 8888 17080 8919
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 18322 8956 18328 8968
rect 18064 8928 18328 8956
rect 17402 8888 17408 8900
rect 17052 8860 17408 8888
rect 16264 8848 16270 8860
rect 17402 8848 17408 8860
rect 17460 8888 17466 8900
rect 17678 8888 17684 8900
rect 17460 8860 17684 8888
rect 17460 8848 17466 8860
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 18064 8897 18092 8928
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18524 8965 18552 8996
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18597 8959 18655 8965
rect 18597 8946 18609 8959
rect 18643 8946 18655 8959
rect 18892 8956 18920 8996
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 20346 9024 20352 9036
rect 19024 8996 19472 9024
rect 19024 8984 19030 8996
rect 19334 8956 19340 8968
rect 18597 8919 18604 8946
rect 18049 8891 18107 8897
rect 18049 8857 18061 8891
rect 18095 8857 18107 8891
rect 18049 8851 18107 8857
rect 18141 8891 18199 8897
rect 18141 8857 18153 8891
rect 18187 8888 18199 8891
rect 18230 8888 18236 8900
rect 18187 8860 18236 8888
rect 18187 8857 18199 8860
rect 18141 8851 18199 8857
rect 13722 8780 13728 8832
rect 13780 8780 13786 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 15746 8820 15752 8832
rect 13964 8792 15752 8820
rect 13964 8780 13970 8792
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 18064 8820 18092 8851
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 18598 8894 18604 8919
rect 18656 8894 18662 8946
rect 18892 8928 19340 8956
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19444 8965 19472 8996
rect 19628 8996 20352 9024
rect 19628 8965 19656 8996
rect 20346 8984 20352 8996
rect 20404 8984 20410 9036
rect 20622 9024 20628 9036
rect 20456 8996 20628 9024
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19577 8959 19656 8965
rect 19577 8925 19589 8959
rect 19623 8928 19656 8959
rect 19794 8956 19800 8968
rect 19755 8928 19800 8956
rect 19623 8925 19635 8928
rect 19577 8919 19635 8925
rect 19794 8916 19800 8928
rect 19852 8916 19858 8968
rect 19935 8959 19993 8965
rect 19935 8925 19947 8959
rect 19981 8956 19993 8959
rect 20456 8956 20484 8996
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 21910 8984 21916 9036
rect 21968 9024 21974 9036
rect 21968 8996 23336 9024
rect 21968 8984 21974 8996
rect 19981 8928 20484 8956
rect 20533 8959 20591 8965
rect 19981 8925 19993 8928
rect 19935 8919 19993 8925
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 22094 8956 22100 8968
rect 20579 8928 22100 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 22094 8916 22100 8928
rect 22152 8916 22158 8968
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 22922 8956 22928 8968
rect 22520 8928 22928 8956
rect 22520 8916 22526 8928
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23308 8965 23336 8996
rect 23293 8959 23351 8965
rect 23293 8925 23305 8959
rect 23339 8925 23351 8959
rect 23293 8919 23351 8925
rect 18693 8891 18751 8897
rect 18693 8857 18705 8891
rect 18739 8888 18751 8891
rect 18782 8888 18788 8900
rect 18739 8860 18788 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 19702 8888 19708 8900
rect 19663 8860 19708 8888
rect 19702 8848 19708 8860
rect 19760 8848 19766 8900
rect 20438 8888 20444 8900
rect 19812 8860 20444 8888
rect 16448 8792 18092 8820
rect 16448 8780 16454 8792
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 19812 8820 19840 8860
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 20898 8848 20904 8900
rect 20956 8888 20962 8900
rect 22833 8891 22891 8897
rect 22833 8888 22845 8891
rect 20956 8860 22845 8888
rect 20956 8848 20962 8860
rect 22833 8857 22845 8860
rect 22879 8857 22891 8891
rect 22833 8851 22891 8857
rect 23385 8891 23443 8897
rect 23385 8857 23397 8891
rect 23431 8857 23443 8891
rect 23385 8851 23443 8857
rect 20346 8820 20352 8832
rect 19116 8792 19840 8820
rect 20307 8792 20352 8820
rect 19116 8780 19122 8792
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 21821 8823 21879 8829
rect 21821 8820 21833 8823
rect 20864 8792 21833 8820
rect 20864 8780 20870 8792
rect 21821 8789 21833 8792
rect 21867 8820 21879 8823
rect 22094 8820 22100 8832
rect 21867 8792 22100 8820
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22094 8780 22100 8792
rect 22152 8780 22158 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 23400 8820 23428 8851
rect 22336 8792 23428 8820
rect 23768 8820 23796 9064
rect 23860 9033 23888 9132
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 23992 9132 24593 9160
rect 23992 9120 23998 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 24946 9120 24952 9172
rect 25004 9160 25010 9172
rect 26602 9160 26608 9172
rect 25004 9132 26464 9160
rect 26563 9132 26608 9160
rect 25004 9120 25010 9132
rect 26436 9092 26464 9132
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 27488 9132 28457 9160
rect 27488 9120 27494 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 28445 9123 28503 9129
rect 28997 9163 29055 9169
rect 28997 9129 29009 9163
rect 29043 9160 29055 9163
rect 32766 9160 32772 9172
rect 29043 9132 32772 9160
rect 29043 9129 29055 9132
rect 28997 9123 29055 9129
rect 32766 9120 32772 9132
rect 32824 9120 32830 9172
rect 32950 9120 32956 9172
rect 33008 9160 33014 9172
rect 33594 9160 33600 9172
rect 33008 9132 33600 9160
rect 33008 9120 33014 9132
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 33870 9120 33876 9172
rect 33928 9160 33934 9172
rect 37826 9160 37832 9172
rect 33928 9132 37832 9160
rect 33928 9120 33934 9132
rect 37826 9120 37832 9132
rect 37884 9120 37890 9172
rect 38657 9163 38715 9169
rect 38657 9129 38669 9163
rect 38703 9160 38715 9163
rect 39114 9160 39120 9172
rect 38703 9132 39120 9160
rect 38703 9129 38715 9132
rect 38657 9123 38715 9129
rect 39114 9120 39120 9132
rect 39172 9120 39178 9172
rect 39592 9132 40086 9160
rect 26970 9092 26976 9104
rect 26436 9064 26976 9092
rect 26970 9052 26976 9064
rect 27028 9052 27034 9104
rect 28166 9052 28172 9104
rect 28224 9092 28230 9104
rect 30742 9092 30748 9104
rect 28224 9064 30748 9092
rect 28224 9052 28230 9064
rect 30742 9052 30748 9064
rect 30800 9052 30806 9104
rect 31754 9052 31760 9104
rect 31812 9092 31818 9104
rect 32125 9095 32183 9101
rect 32125 9092 32137 9095
rect 31812 9064 32137 9092
rect 31812 9052 31818 9064
rect 32125 9061 32137 9064
rect 32171 9092 32183 9095
rect 32674 9092 32680 9104
rect 32171 9064 32680 9092
rect 32171 9061 32183 9064
rect 32125 9055 32183 9061
rect 32674 9052 32680 9064
rect 32732 9052 32738 9104
rect 32784 9092 32812 9120
rect 32784 9064 33364 9092
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 8993 23903 9027
rect 25222 9024 25228 9036
rect 25183 8996 25228 9024
rect 23845 8987 23903 8993
rect 25222 8984 25228 8996
rect 25280 8984 25286 9036
rect 26418 8984 26424 9036
rect 26476 9024 26482 9036
rect 32950 9024 32956 9036
rect 26476 8996 27200 9024
rect 26476 8984 26482 8996
rect 23934 8916 23940 8968
rect 23992 8956 23998 8968
rect 24578 8956 24584 8968
rect 23992 8928 24584 8956
rect 23992 8916 23998 8928
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 24762 8956 24768 8968
rect 24723 8928 24768 8956
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 25240 8956 25268 8984
rect 27172 8968 27200 8996
rect 28092 8996 29684 9024
rect 32911 8996 32956 9024
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 25240 8928 27077 8956
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 27154 8916 27160 8968
rect 27212 8956 27218 8968
rect 28092 8956 28120 8996
rect 29656 8968 29684 8996
rect 32950 8984 32956 8996
rect 33008 8984 33014 9036
rect 33336 9024 33364 9064
rect 33410 9052 33416 9104
rect 33468 9092 33474 9104
rect 35802 9092 35808 9104
rect 33468 9064 35808 9092
rect 33468 9052 33474 9064
rect 35802 9052 35808 9064
rect 35860 9052 35866 9104
rect 37182 9052 37188 9104
rect 37240 9092 37246 9104
rect 39592 9092 39620 9132
rect 37240 9064 39620 9092
rect 40058 9092 40086 9132
rect 41414 9092 41420 9104
rect 40058 9064 41420 9092
rect 37240 9052 37246 9064
rect 41414 9052 41420 9064
rect 41472 9052 41478 9104
rect 43990 9092 43996 9104
rect 43951 9064 43996 9092
rect 43990 9052 43996 9064
rect 44048 9052 44054 9104
rect 34149 9027 34207 9033
rect 33336 8996 34100 9024
rect 27212 8928 28120 8956
rect 27212 8916 27218 8928
rect 28718 8916 28724 8968
rect 28776 8956 28782 8968
rect 28997 8959 29055 8965
rect 28997 8956 29009 8959
rect 28776 8928 29009 8956
rect 28776 8916 28782 8928
rect 28997 8925 29009 8928
rect 29043 8956 29055 8959
rect 29086 8956 29092 8968
rect 29043 8928 29092 8956
rect 29043 8925 29055 8928
rect 28997 8919 29055 8925
rect 29086 8916 29092 8928
rect 29144 8916 29150 8968
rect 29181 8959 29239 8965
rect 29181 8925 29193 8959
rect 29227 8925 29239 8959
rect 29181 8919 29239 8925
rect 25492 8891 25550 8897
rect 25492 8857 25504 8891
rect 25538 8888 25550 8891
rect 27332 8891 27390 8897
rect 25538 8860 27292 8888
rect 25538 8857 25550 8860
rect 25492 8851 25550 8857
rect 26694 8820 26700 8832
rect 23768 8792 26700 8820
rect 22336 8780 22342 8792
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 27264 8820 27292 8860
rect 27332 8857 27344 8891
rect 27378 8888 27390 8891
rect 28350 8888 28356 8900
rect 27378 8860 28356 8888
rect 27378 8857 27390 8860
rect 27332 8851 27390 8857
rect 28350 8848 28356 8860
rect 28408 8848 28414 8900
rect 28902 8848 28908 8900
rect 28960 8888 28966 8900
rect 29196 8888 29224 8919
rect 29638 8916 29644 8968
rect 29696 8956 29702 8968
rect 29733 8959 29791 8965
rect 29733 8956 29745 8959
rect 29696 8928 29745 8956
rect 29696 8916 29702 8928
rect 29733 8925 29745 8928
rect 29779 8925 29791 8959
rect 29733 8919 29791 8925
rect 29822 8916 29828 8968
rect 29880 8956 29886 8968
rect 30742 8956 30748 8968
rect 29880 8928 29925 8956
rect 30703 8928 30748 8956
rect 29880 8916 29886 8928
rect 30742 8916 30748 8928
rect 30800 8916 30806 8968
rect 31021 8959 31079 8965
rect 31021 8925 31033 8959
rect 31067 8956 31079 8959
rect 31386 8956 31392 8968
rect 31067 8928 31392 8956
rect 31067 8925 31079 8928
rect 31021 8919 31079 8925
rect 31386 8916 31392 8928
rect 31444 8916 31450 8968
rect 33137 8959 33195 8965
rect 33137 8925 33149 8959
rect 33183 8956 33195 8959
rect 33502 8956 33508 8968
rect 33183 8928 33508 8956
rect 33183 8925 33195 8928
rect 33137 8919 33195 8925
rect 33502 8916 33508 8928
rect 33560 8916 33566 8968
rect 33778 8916 33784 8968
rect 33836 8956 33842 8968
rect 33873 8959 33931 8965
rect 33873 8956 33885 8959
rect 33836 8928 33885 8956
rect 33836 8916 33842 8928
rect 33873 8925 33885 8928
rect 33919 8925 33931 8959
rect 33873 8919 33931 8925
rect 28960 8860 29224 8888
rect 28960 8848 28966 8860
rect 29362 8848 29368 8900
rect 29420 8888 29426 8900
rect 29546 8888 29552 8900
rect 29420 8860 29552 8888
rect 29420 8848 29426 8860
rect 29546 8848 29552 8860
rect 29604 8888 29610 8900
rect 30285 8891 30343 8897
rect 30285 8888 30297 8891
rect 29604 8860 30297 8888
rect 29604 8848 29610 8860
rect 30285 8857 30297 8860
rect 30331 8857 30343 8891
rect 30285 8851 30343 8857
rect 33413 8891 33471 8897
rect 33413 8857 33425 8891
rect 33459 8857 33471 8891
rect 34072 8888 34100 8996
rect 34149 8993 34161 9027
rect 34195 9024 34207 9027
rect 35897 9027 35955 9033
rect 35897 9024 35909 9027
rect 34195 8996 34652 9024
rect 34195 8993 34207 8996
rect 34149 8987 34207 8993
rect 34624 8888 34652 8996
rect 34716 8996 35909 9024
rect 34716 8968 34744 8996
rect 35897 8993 35909 8996
rect 35943 9024 35955 9027
rect 37090 9024 37096 9036
rect 35943 8996 37096 9024
rect 35943 8993 35955 8996
rect 35897 8987 35955 8993
rect 37090 8984 37096 8996
rect 37148 8984 37154 9036
rect 37826 8984 37832 9036
rect 37884 9024 37890 9036
rect 39574 9024 39580 9036
rect 37884 8996 39580 9024
rect 37884 8984 37890 8996
rect 39574 8984 39580 8996
rect 39632 8984 39638 9036
rect 40586 8984 40592 9036
rect 40644 9024 40650 9036
rect 41049 9027 41107 9033
rect 41049 9024 41061 9027
rect 40644 8996 41061 9024
rect 40644 8984 40650 8996
rect 41049 8993 41061 8996
rect 41095 9024 41107 9027
rect 41322 9024 41328 9036
rect 41095 8996 41328 9024
rect 41095 8993 41107 8996
rect 41049 8987 41107 8993
rect 41322 8984 41328 8996
rect 41380 9024 41386 9036
rect 41598 9024 41604 9036
rect 41380 8996 41604 9024
rect 41380 8984 41386 8996
rect 41598 8984 41604 8996
rect 41656 8984 41662 9036
rect 34698 8916 34704 8968
rect 34756 8916 34762 8968
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 34848 8928 34897 8956
rect 34848 8916 34854 8928
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 34974 8916 34980 8968
rect 35032 8956 35038 8968
rect 35161 8959 35219 8965
rect 35161 8956 35173 8959
rect 35032 8928 35173 8956
rect 35032 8916 35038 8928
rect 35161 8925 35173 8928
rect 35207 8925 35219 8959
rect 35161 8919 35219 8925
rect 35434 8916 35440 8968
rect 35492 8956 35498 8968
rect 35618 8956 35624 8968
rect 35492 8928 35624 8956
rect 35492 8916 35498 8928
rect 35618 8916 35624 8928
rect 35676 8916 35682 8968
rect 35986 8956 35992 8968
rect 35866 8928 35992 8956
rect 35866 8888 35894 8928
rect 35986 8916 35992 8928
rect 36044 8916 36050 8968
rect 36173 8959 36231 8965
rect 36173 8925 36185 8959
rect 36219 8956 36231 8959
rect 38010 8956 38016 8968
rect 36219 8928 37872 8956
rect 37971 8928 38016 8956
rect 36219 8925 36231 8928
rect 36173 8919 36231 8925
rect 37550 8888 37556 8900
rect 34072 8860 34560 8888
rect 34624 8860 35894 8888
rect 37511 8860 37556 8888
rect 33413 8851 33471 8857
rect 30834 8820 30840 8832
rect 27264 8792 30840 8820
rect 30834 8780 30840 8792
rect 30892 8780 30898 8832
rect 31754 8780 31760 8832
rect 31812 8820 31818 8832
rect 33321 8823 33379 8829
rect 33321 8820 33333 8823
rect 31812 8792 33333 8820
rect 31812 8780 31818 8792
rect 33321 8789 33333 8792
rect 33367 8789 33379 8823
rect 33428 8820 33456 8851
rect 34054 8820 34060 8832
rect 33428 8792 34060 8820
rect 33321 8783 33379 8789
rect 34054 8780 34060 8792
rect 34112 8780 34118 8832
rect 34532 8820 34560 8860
rect 37550 8848 37556 8860
rect 37608 8848 37614 8900
rect 35158 8820 35164 8832
rect 34532 8792 35164 8820
rect 35158 8780 35164 8792
rect 35216 8780 35222 8832
rect 35434 8780 35440 8832
rect 35492 8820 35498 8832
rect 37642 8820 37648 8832
rect 35492 8792 37648 8820
rect 35492 8780 35498 8792
rect 37642 8780 37648 8792
rect 37700 8780 37706 8832
rect 37844 8820 37872 8928
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 38102 8916 38108 8968
rect 38160 8956 38166 8968
rect 38378 8956 38384 8968
rect 38160 8928 38205 8956
rect 38339 8928 38384 8956
rect 38160 8916 38166 8928
rect 38378 8916 38384 8928
rect 38436 8916 38442 8968
rect 38470 8916 38476 8968
rect 38528 8965 38534 8968
rect 38528 8956 38536 8965
rect 38528 8928 38573 8956
rect 38528 8919 38536 8928
rect 38528 8916 38534 8919
rect 38930 8916 38936 8968
rect 38988 8956 38994 8968
rect 39485 8959 39543 8965
rect 39485 8956 39497 8959
rect 38988 8928 39497 8956
rect 38988 8916 38994 8928
rect 39485 8925 39497 8928
rect 39531 8925 39543 8959
rect 39485 8919 39543 8925
rect 39758 8916 39764 8968
rect 39816 8956 39822 8968
rect 40037 8959 40095 8965
rect 40037 8956 40049 8959
rect 39816 8928 40049 8956
rect 39816 8916 39822 8928
rect 40037 8925 40049 8928
rect 40083 8925 40095 8959
rect 40037 8919 40095 8925
rect 40233 8959 40291 8965
rect 40233 8925 40245 8959
rect 40279 8956 40291 8959
rect 40402 8956 40408 8968
rect 40279 8928 40408 8956
rect 40279 8925 40291 8928
rect 40233 8919 40291 8925
rect 40402 8916 40408 8928
rect 40460 8916 40466 8968
rect 40678 8916 40684 8968
rect 40736 8956 40742 8968
rect 40773 8959 40831 8965
rect 40773 8956 40785 8959
rect 40736 8928 40785 8956
rect 40736 8916 40742 8928
rect 40773 8925 40785 8928
rect 40819 8956 40831 8959
rect 41138 8956 41144 8968
rect 40819 8928 41144 8956
rect 40819 8925 40831 8928
rect 40773 8919 40831 8925
rect 41138 8916 41144 8928
rect 41196 8916 41202 8968
rect 42613 8959 42671 8965
rect 42613 8925 42625 8959
rect 42659 8956 42671 8959
rect 42702 8956 42708 8968
rect 42659 8928 42708 8956
rect 42659 8925 42671 8928
rect 42613 8919 42671 8925
rect 42702 8916 42708 8928
rect 42760 8916 42766 8968
rect 42880 8959 42938 8965
rect 42880 8925 42892 8959
rect 42926 8956 42938 8959
rect 44542 8956 44548 8968
rect 42926 8928 44548 8956
rect 42926 8925 42938 8928
rect 42880 8919 42938 8925
rect 44542 8916 44548 8928
rect 44600 8916 44606 8968
rect 57057 8959 57115 8965
rect 57057 8925 57069 8959
rect 57103 8956 57115 8959
rect 57146 8956 57152 8968
rect 57103 8928 57152 8956
rect 57103 8925 57115 8928
rect 57057 8919 57115 8925
rect 57146 8916 57152 8928
rect 57204 8916 57210 8968
rect 57241 8959 57299 8965
rect 57241 8925 57253 8959
rect 57287 8956 57299 8959
rect 57885 8959 57943 8965
rect 57885 8956 57897 8959
rect 57287 8928 57897 8956
rect 57287 8925 57299 8928
rect 57241 8919 57299 8925
rect 57885 8925 57897 8928
rect 57931 8956 57943 8959
rect 58250 8956 58256 8968
rect 57931 8928 58256 8956
rect 57931 8925 57943 8928
rect 57885 8919 57943 8925
rect 58250 8916 58256 8928
rect 58308 8916 58314 8968
rect 37918 8848 37924 8900
rect 37976 8888 37982 8900
rect 38289 8891 38347 8897
rect 38289 8888 38301 8891
rect 37976 8860 38301 8888
rect 37976 8848 37982 8860
rect 38289 8857 38301 8860
rect 38335 8888 38347 8891
rect 39114 8888 39120 8900
rect 38335 8860 38976 8888
rect 39075 8860 39120 8888
rect 38335 8857 38347 8860
rect 38289 8851 38347 8857
rect 38838 8820 38844 8832
rect 37844 8792 38844 8820
rect 38838 8780 38844 8792
rect 38896 8780 38902 8832
rect 38948 8820 38976 8860
rect 39114 8848 39120 8860
rect 39172 8848 39178 8900
rect 39301 8891 39359 8897
rect 39301 8857 39313 8891
rect 39347 8888 39359 8891
rect 39574 8888 39580 8900
rect 39347 8860 39580 8888
rect 39347 8857 39359 8860
rect 39301 8851 39359 8857
rect 39574 8848 39580 8860
rect 39632 8848 39638 8900
rect 39850 8848 39856 8900
rect 39908 8888 39914 8900
rect 40129 8891 40187 8897
rect 40129 8888 40141 8891
rect 39908 8860 40141 8888
rect 39908 8848 39914 8860
rect 40129 8857 40141 8860
rect 40175 8857 40187 8891
rect 40129 8851 40187 8857
rect 42978 8848 42984 8900
rect 43036 8888 43042 8900
rect 44082 8888 44088 8900
rect 43036 8860 44088 8888
rect 43036 8848 43042 8860
rect 44082 8848 44088 8860
rect 44140 8848 44146 8900
rect 58158 8888 58164 8900
rect 58119 8860 58164 8888
rect 58158 8848 58164 8860
rect 58216 8848 58222 8900
rect 40678 8820 40684 8832
rect 38948 8792 40684 8820
rect 40678 8780 40684 8792
rect 40736 8780 40742 8832
rect 56594 8780 56600 8832
rect 56652 8820 56658 8832
rect 57149 8823 57207 8829
rect 57149 8820 57161 8823
rect 56652 8792 57161 8820
rect 56652 8780 56658 8792
rect 57149 8789 57161 8792
rect 57195 8789 57207 8823
rect 57149 8783 57207 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15252 8588 16221 8616
rect 15252 8576 15258 8588
rect 16209 8585 16221 8588
rect 16255 8616 16267 8619
rect 16390 8616 16396 8628
rect 16255 8588 16396 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 18598 8616 18604 8628
rect 18156 8588 18604 8616
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 8662 8548 8668 8560
rect 2556 8520 8668 8548
rect 2556 8508 2562 8520
rect 8662 8508 8668 8520
rect 8720 8548 8726 8560
rect 17313 8551 17371 8557
rect 8720 8520 17080 8548
rect 8720 8508 8726 8520
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 10413 8483 10471 8489
rect 1627 8452 2774 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2746 8412 2774 8452
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 13630 8480 13636 8492
rect 10459 8452 13636 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 17052 8489 17080 8520
rect 17313 8517 17325 8551
rect 17359 8548 17371 8551
rect 17402 8548 17408 8560
rect 17359 8520 17408 8548
rect 17359 8517 17371 8520
rect 17313 8511 17371 8517
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 2746 8384 10149 8412
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10318 8412 10324 8424
rect 10279 8384 10324 8412
rect 10137 8375 10195 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 10652 8384 10697 8412
rect 10652 8372 10658 8384
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12066 8412 12072 8424
rect 11296 8384 12072 8412
rect 11296 8372 11302 8384
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 16040 8276 16068 8443
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 18156 8489 18184 8588
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18693 8619 18751 8625
rect 18693 8585 18705 8619
rect 18739 8616 18751 8619
rect 19242 8616 19248 8628
rect 18739 8588 19248 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 21450 8616 21456 8628
rect 19392 8588 19932 8616
rect 21411 8588 21456 8616
rect 19392 8576 19398 8588
rect 18509 8551 18567 8557
rect 18509 8517 18521 8551
rect 18555 8548 18567 8551
rect 18782 8548 18788 8560
rect 18555 8520 18788 8548
rect 18555 8517 18567 8520
rect 18509 8511 18567 8517
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 17184 8452 18153 8480
rect 17184 8440 17190 8452
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 19334 8480 19340 8492
rect 18380 8452 19340 8480
rect 18380 8440 18386 8452
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19904 8489 19932 8588
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 24946 8616 24952 8628
rect 22066 8588 24952 8616
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 20806 8548 20812 8560
rect 20128 8520 20812 8548
rect 20128 8508 20134 8520
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19444 8452 19625 8480
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 19444 8412 19472 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19613 8443 19671 8449
rect 19812 8452 19901 8480
rect 19812 8424 19840 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20254 8480 20260 8492
rect 20036 8452 20081 8480
rect 20215 8452 20260 8480
rect 20036 8440 20042 8452
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20456 8489 20484 8520
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 22066 8548 22094 8588
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25406 8616 25412 8628
rect 25148 8588 25412 8616
rect 25148 8557 25176 8588
rect 25406 8576 25412 8588
rect 25464 8616 25470 8628
rect 26970 8616 26976 8628
rect 25464 8588 26976 8616
rect 25464 8576 25470 8588
rect 26970 8576 26976 8588
rect 27028 8576 27034 8628
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27525 8619 27583 8625
rect 27525 8616 27537 8619
rect 27120 8588 27537 8616
rect 27120 8576 27126 8588
rect 27525 8585 27537 8588
rect 27571 8585 27583 8619
rect 28350 8616 28356 8628
rect 28311 8588 28356 8616
rect 27525 8579 27583 8585
rect 28350 8576 28356 8588
rect 28408 8576 28414 8628
rect 28442 8576 28448 8628
rect 28500 8616 28506 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 28500 8588 28733 8616
rect 28500 8576 28506 8588
rect 28721 8585 28733 8588
rect 28767 8585 28779 8619
rect 28721 8579 28779 8585
rect 29086 8576 29092 8628
rect 29144 8616 29150 8628
rect 31294 8616 31300 8628
rect 29144 8588 31300 8616
rect 29144 8576 29150 8588
rect 31294 8576 31300 8588
rect 31352 8576 31358 8628
rect 33226 8616 33232 8628
rect 33187 8588 33232 8616
rect 33226 8576 33232 8588
rect 33284 8576 33290 8628
rect 35713 8619 35771 8625
rect 35713 8616 35725 8619
rect 33336 8588 35725 8616
rect 21192 8520 22094 8548
rect 25133 8551 25191 8557
rect 21192 8489 21220 8520
rect 25133 8517 25145 8551
rect 25179 8517 25191 8551
rect 27154 8548 27160 8560
rect 25133 8511 25191 8517
rect 25976 8520 27160 8548
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21818 8480 21824 8492
rect 21315 8452 21824 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 23750 8480 23756 8492
rect 23711 8452 23756 8480
rect 22097 8443 22155 8449
rect 16724 8384 19472 8412
rect 16724 8372 16730 8384
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 22112 8412 22140 8443
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8480 25651 8483
rect 25774 8480 25780 8492
rect 25639 8452 25780 8480
rect 25639 8449 25651 8452
rect 25593 8443 25651 8449
rect 25774 8440 25780 8452
rect 25832 8440 25838 8492
rect 25976 8489 26004 8520
rect 27154 8508 27160 8520
rect 27212 8508 27218 8560
rect 27246 8508 27252 8560
rect 27304 8548 27310 8560
rect 27617 8551 27675 8557
rect 27617 8548 27629 8551
rect 27304 8520 27629 8548
rect 27304 8508 27310 8520
rect 27617 8517 27629 8520
rect 27663 8517 27675 8551
rect 32306 8548 32312 8560
rect 27617 8511 27675 8517
rect 29840 8520 32312 8548
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8480 26111 8483
rect 26142 8480 26148 8492
rect 26099 8452 26148 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 27430 8440 27436 8492
rect 27488 8480 27494 8492
rect 28813 8483 28871 8489
rect 28813 8480 28825 8483
rect 27488 8452 28825 8480
rect 27488 8440 27494 8452
rect 28813 8449 28825 8452
rect 28859 8449 28871 8483
rect 29730 8480 29736 8492
rect 28813 8443 28871 8449
rect 28920 8452 29736 8480
rect 22830 8412 22836 8424
rect 21048 8384 22140 8412
rect 22791 8384 22836 8412
rect 21048 8372 21054 8384
rect 22830 8372 22836 8384
rect 22888 8372 22894 8424
rect 24026 8372 24032 8424
rect 24084 8412 24090 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 24084 8384 24501 8412
rect 24084 8372 24090 8384
rect 24489 8381 24501 8384
rect 24535 8412 24547 8415
rect 24946 8412 24952 8424
rect 24535 8384 24952 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25866 8412 25872 8424
rect 25096 8384 25872 8412
rect 25096 8372 25102 8384
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 27801 8415 27859 8421
rect 26252 8384 27292 8412
rect 16758 8304 16764 8356
rect 16816 8344 16822 8356
rect 26252 8344 26280 8384
rect 16816 8316 26280 8344
rect 16816 8304 16822 8316
rect 26326 8304 26332 8356
rect 26384 8344 26390 8356
rect 27157 8347 27215 8353
rect 27157 8344 27169 8347
rect 26384 8316 27169 8344
rect 26384 8304 26390 8316
rect 27157 8313 27169 8316
rect 27203 8313 27215 8347
rect 27264 8344 27292 8384
rect 27801 8381 27813 8415
rect 27847 8412 27859 8415
rect 27982 8412 27988 8424
rect 27847 8384 27988 8412
rect 27847 8381 27859 8384
rect 27801 8375 27859 8381
rect 27982 8372 27988 8384
rect 28040 8372 28046 8424
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 28920 8421 28948 8452
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 29840 8489 29868 8520
rect 32306 8508 32312 8520
rect 32364 8508 32370 8560
rect 32582 8548 32588 8560
rect 32543 8520 32588 8548
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 32950 8508 32956 8560
rect 33008 8548 33014 8560
rect 33336 8548 33364 8588
rect 35713 8585 35725 8588
rect 35759 8585 35771 8619
rect 35713 8579 35771 8585
rect 37642 8576 37648 8628
rect 37700 8616 37706 8628
rect 39390 8616 39396 8628
rect 37700 8588 38424 8616
rect 39351 8588 39396 8616
rect 37700 8576 37706 8588
rect 33008 8520 33364 8548
rect 33008 8508 33014 8520
rect 33410 8508 33416 8560
rect 33468 8548 33474 8560
rect 33505 8551 33563 8557
rect 33505 8548 33517 8551
rect 33468 8520 33517 8548
rect 33468 8508 33474 8520
rect 33505 8517 33517 8520
rect 33551 8517 33563 8551
rect 35066 8548 35072 8560
rect 33505 8511 33563 8517
rect 34532 8520 35072 8548
rect 30098 8489 30104 8492
rect 29825 8483 29883 8489
rect 29825 8449 29837 8483
rect 29871 8449 29883 8483
rect 30092 8480 30104 8489
rect 30059 8452 30104 8480
rect 29825 8443 29883 8449
rect 30092 8443 30104 8452
rect 30098 8440 30104 8443
rect 30156 8440 30162 8492
rect 31478 8440 31484 8492
rect 31536 8480 31542 8492
rect 32217 8483 32275 8489
rect 32217 8480 32229 8483
rect 31536 8452 32229 8480
rect 31536 8440 31542 8452
rect 32217 8449 32229 8452
rect 32263 8449 32275 8483
rect 33686 8480 33692 8492
rect 33647 8452 33692 8480
rect 32217 8443 32275 8449
rect 33686 8440 33692 8452
rect 33744 8440 33750 8492
rect 34532 8489 34560 8520
rect 35066 8508 35072 8520
rect 35124 8508 35130 8560
rect 36078 8508 36084 8560
rect 36136 8548 36142 8560
rect 36906 8548 36912 8560
rect 36136 8520 36773 8548
rect 36136 8508 36142 8520
rect 33781 8483 33839 8489
rect 33781 8449 33793 8483
rect 33827 8449 33839 8483
rect 33781 8443 33839 8449
rect 34425 8483 34483 8489
rect 34425 8449 34437 8483
rect 34471 8449 34483 8483
rect 34425 8443 34483 8449
rect 34517 8483 34575 8489
rect 34517 8449 34529 8483
rect 34563 8449 34575 8483
rect 34517 8443 34575 8449
rect 34641 8483 34699 8489
rect 34641 8449 34653 8483
rect 34687 8449 34699 8483
rect 34641 8443 34699 8449
rect 28905 8415 28963 8421
rect 28905 8412 28917 8415
rect 28776 8384 28917 8412
rect 28776 8372 28782 8384
rect 28905 8381 28917 8384
rect 28951 8381 28963 8415
rect 28905 8375 28963 8381
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 32398 8412 32404 8424
rect 31076 8384 32404 8412
rect 31076 8372 31082 8384
rect 32398 8372 32404 8384
rect 32456 8372 32462 8424
rect 33318 8372 33324 8424
rect 33376 8412 33382 8424
rect 33796 8412 33824 8443
rect 34440 8412 34468 8443
rect 33376 8384 33824 8412
rect 33980 8384 34468 8412
rect 33376 8372 33382 8384
rect 29454 8344 29460 8356
rect 27264 8316 29460 8344
rect 27157 8307 27215 8313
rect 29454 8304 29460 8316
rect 29512 8304 29518 8356
rect 33980 8353 34008 8384
rect 33965 8347 34023 8353
rect 33965 8313 33977 8347
rect 34011 8313 34023 8347
rect 34656 8344 34684 8443
rect 35158 8440 35164 8492
rect 35216 8480 35222 8492
rect 35621 8483 35679 8489
rect 35621 8480 35633 8483
rect 35216 8452 35633 8480
rect 35216 8440 35222 8452
rect 35621 8449 35633 8452
rect 35667 8449 35679 8483
rect 36262 8480 36268 8492
rect 36223 8452 36268 8480
rect 35621 8443 35679 8449
rect 36262 8440 36268 8452
rect 36320 8440 36326 8492
rect 36446 8489 36452 8492
rect 36413 8483 36452 8489
rect 36413 8449 36425 8483
rect 36413 8443 36452 8449
rect 36446 8440 36452 8443
rect 36504 8440 36510 8492
rect 36745 8489 36773 8520
rect 36832 8520 36912 8548
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8449 36599 8483
rect 36541 8443 36599 8449
rect 36633 8483 36691 8489
rect 36633 8449 36645 8483
rect 36679 8449 36691 8483
rect 36633 8443 36691 8449
rect 36730 8483 36788 8489
rect 36730 8449 36742 8483
rect 36776 8449 36788 8483
rect 36730 8443 36788 8449
rect 34882 8372 34888 8424
rect 34940 8412 34946 8424
rect 34940 8384 34985 8412
rect 34940 8372 34946 8384
rect 35710 8372 35716 8424
rect 35768 8412 35774 8424
rect 36556 8412 36584 8443
rect 35768 8384 36584 8412
rect 36648 8412 36676 8443
rect 36832 8412 36860 8520
rect 36906 8508 36912 8520
rect 36964 8508 36970 8560
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38258 8551 38316 8557
rect 38258 8548 38270 8551
rect 37516 8520 38270 8548
rect 37516 8508 37522 8520
rect 38258 8517 38270 8520
rect 38304 8517 38316 8551
rect 38258 8511 38316 8517
rect 37090 8440 37096 8492
rect 37148 8480 37154 8492
rect 38013 8483 38071 8489
rect 38013 8480 38025 8483
rect 37148 8452 38025 8480
rect 37148 8440 37154 8452
rect 38013 8449 38025 8452
rect 38059 8449 38071 8483
rect 38396 8480 38424 8588
rect 39390 8576 39396 8588
rect 39448 8576 39454 8628
rect 39574 8576 39580 8628
rect 39632 8616 39638 8628
rect 40586 8616 40592 8628
rect 39632 8588 40592 8616
rect 39632 8576 39638 8588
rect 40586 8576 40592 8588
rect 40644 8576 40650 8628
rect 41230 8616 41236 8628
rect 41191 8588 41236 8616
rect 41230 8576 41236 8588
rect 41288 8576 41294 8628
rect 52638 8616 52644 8628
rect 41524 8588 52644 8616
rect 38470 8508 38476 8560
rect 38528 8548 38534 8560
rect 39666 8548 39672 8560
rect 38528 8520 39672 8548
rect 38528 8508 38534 8520
rect 39666 8508 39672 8520
rect 39724 8508 39730 8560
rect 40405 8551 40463 8557
rect 40405 8517 40417 8551
rect 40451 8548 40463 8551
rect 40862 8548 40868 8560
rect 40451 8520 40868 8548
rect 40451 8517 40463 8520
rect 40405 8511 40463 8517
rect 40862 8508 40868 8520
rect 40920 8508 40926 8560
rect 40034 8480 40040 8492
rect 38396 8452 40040 8480
rect 38013 8443 38071 8449
rect 40034 8440 40040 8452
rect 40092 8440 40098 8492
rect 40130 8483 40188 8489
rect 40130 8449 40142 8483
rect 40176 8449 40188 8483
rect 40310 8480 40316 8492
rect 40271 8452 40316 8480
rect 40130 8443 40188 8449
rect 36648 8384 36860 8412
rect 35768 8372 35774 8384
rect 34974 8344 34980 8356
rect 34656 8316 34980 8344
rect 33965 8307 34023 8313
rect 34974 8304 34980 8316
rect 35032 8304 35038 8356
rect 35066 8304 35072 8356
rect 35124 8344 35130 8356
rect 37182 8344 37188 8356
rect 35124 8316 37188 8344
rect 35124 8304 35130 8316
rect 37182 8304 37188 8316
rect 37240 8304 37246 8356
rect 40034 8304 40040 8356
rect 40092 8344 40098 8356
rect 40145 8344 40173 8443
rect 40310 8440 40316 8452
rect 40368 8440 40374 8492
rect 40499 8440 40505 8492
rect 40557 8480 40563 8492
rect 40557 8452 40602 8480
rect 40557 8440 40563 8452
rect 41322 8440 41328 8492
rect 41380 8480 41386 8492
rect 41524 8489 41552 8588
rect 52638 8576 52644 8588
rect 52696 8576 52702 8628
rect 41417 8483 41475 8489
rect 41417 8480 41429 8483
rect 41380 8452 41429 8480
rect 41380 8440 41386 8452
rect 41417 8449 41429 8452
rect 41463 8449 41475 8483
rect 41417 8443 41475 8449
rect 41509 8483 41567 8489
rect 41509 8449 41521 8483
rect 41555 8449 41567 8483
rect 41690 8480 41696 8492
rect 41651 8452 41696 8480
rect 41509 8443 41567 8449
rect 41690 8440 41696 8452
rect 41748 8440 41754 8492
rect 41785 8483 41843 8489
rect 41785 8449 41797 8483
rect 41831 8449 41843 8483
rect 41785 8443 41843 8449
rect 42705 8483 42763 8489
rect 42705 8449 42717 8483
rect 42751 8480 42763 8483
rect 43622 8480 43628 8492
rect 42751 8452 43484 8480
rect 43583 8452 43628 8480
rect 42751 8449 42763 8452
rect 42705 8443 42763 8449
rect 40092 8316 40173 8344
rect 40681 8347 40739 8353
rect 40092 8304 40098 8316
rect 40681 8313 40693 8347
rect 40727 8344 40739 8347
rect 41800 8344 41828 8443
rect 42978 8412 42984 8424
rect 42939 8384 42984 8412
rect 42978 8372 42984 8384
rect 43036 8372 43042 8424
rect 43456 8412 43484 8452
rect 43622 8440 43628 8452
rect 43680 8440 43686 8492
rect 44082 8440 44088 8492
rect 44140 8480 44146 8492
rect 44545 8483 44603 8489
rect 44545 8480 44557 8483
rect 44140 8452 44557 8480
rect 44140 8440 44146 8452
rect 44545 8449 44557 8452
rect 44591 8449 44603 8483
rect 57146 8480 57152 8492
rect 57107 8452 57152 8480
rect 44545 8443 44603 8449
rect 57146 8440 57152 8452
rect 57204 8440 57210 8492
rect 43806 8412 43812 8424
rect 43456 8384 43812 8412
rect 43806 8372 43812 8384
rect 43864 8372 43870 8424
rect 44174 8372 44180 8424
rect 44232 8412 44238 8424
rect 44729 8415 44787 8421
rect 44729 8412 44741 8415
rect 44232 8384 44741 8412
rect 44232 8372 44238 8384
rect 44729 8381 44741 8384
rect 44775 8381 44787 8415
rect 44729 8375 44787 8381
rect 40727 8316 41828 8344
rect 40727 8313 40739 8316
rect 40681 8307 40739 8313
rect 42610 8304 42616 8356
rect 42668 8344 42674 8356
rect 57333 8347 57391 8353
rect 57333 8344 57345 8347
rect 42668 8316 57345 8344
rect 42668 8304 42674 8316
rect 57333 8313 57345 8316
rect 57379 8313 57391 8347
rect 57333 8307 57391 8313
rect 18230 8276 18236 8288
rect 16040 8248 18236 8276
rect 18230 8236 18236 8248
rect 18288 8276 18294 8288
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 18288 8248 18521 8276
rect 18288 8236 18294 8248
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 19242 8276 19248 8288
rect 19203 8248 19248 8276
rect 18509 8239 18567 8245
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 27522 8276 27528 8288
rect 19760 8248 27528 8276
rect 19760 8236 19766 8248
rect 27522 8236 27528 8248
rect 27580 8236 27586 8288
rect 28626 8236 28632 8288
rect 28684 8276 28690 8288
rect 29086 8276 29092 8288
rect 28684 8248 29092 8276
rect 28684 8236 28690 8248
rect 29086 8236 29092 8248
rect 29144 8236 29150 8288
rect 31202 8276 31208 8288
rect 31163 8248 31208 8276
rect 31202 8236 31208 8248
rect 31260 8236 31266 8288
rect 33226 8236 33232 8288
rect 33284 8276 33290 8288
rect 33505 8279 33563 8285
rect 33505 8276 33517 8279
rect 33284 8248 33517 8276
rect 33284 8236 33290 8248
rect 33505 8245 33517 8248
rect 33551 8276 33563 8279
rect 34333 8279 34391 8285
rect 34333 8276 34345 8279
rect 33551 8248 34345 8276
rect 33551 8245 33563 8248
rect 33505 8239 33563 8245
rect 34333 8245 34345 8248
rect 34379 8245 34391 8279
rect 34333 8239 34391 8245
rect 35802 8236 35808 8288
rect 35860 8276 35866 8288
rect 36170 8276 36176 8288
rect 35860 8248 36176 8276
rect 35860 8236 35866 8248
rect 36170 8236 36176 8248
rect 36228 8236 36234 8288
rect 36262 8236 36268 8288
rect 36320 8276 36326 8288
rect 36909 8279 36967 8285
rect 36909 8276 36921 8279
rect 36320 8248 36921 8276
rect 36320 8236 36326 8248
rect 36909 8245 36921 8248
rect 36955 8245 36967 8279
rect 36909 8239 36967 8245
rect 37826 8236 37832 8288
rect 37884 8276 37890 8288
rect 39114 8276 39120 8288
rect 37884 8248 39120 8276
rect 37884 8236 37890 8248
rect 39114 8236 39120 8248
rect 39172 8276 39178 8288
rect 40126 8276 40132 8288
rect 39172 8248 40132 8276
rect 39172 8236 39178 8248
rect 40126 8236 40132 8248
rect 40184 8276 40190 8288
rect 41690 8276 41696 8288
rect 40184 8248 41696 8276
rect 40184 8236 40190 8248
rect 41690 8236 41696 8248
rect 41748 8276 41754 8288
rect 44174 8276 44180 8288
rect 41748 8248 44180 8276
rect 41748 8236 41754 8248
rect 44174 8236 44180 8248
rect 44232 8236 44238 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10594 8072 10600 8084
rect 10275 8044 10600 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 16666 8072 16672 8084
rect 16623 8044 16672 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17129 8075 17187 8081
rect 17129 8041 17141 8075
rect 17175 8072 17187 8075
rect 20714 8072 20720 8084
rect 17175 8044 20720 8072
rect 17175 8041 17187 8044
rect 17129 8035 17187 8041
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 21082 8072 21088 8084
rect 21008 8044 21088 8072
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 11146 8004 11152 8016
rect 10183 7976 11152 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 15746 7964 15752 8016
rect 15804 8004 15810 8016
rect 15804 7976 17540 8004
rect 15804 7964 15810 7976
rect 17126 7936 17132 7948
rect 16500 7908 17132 7936
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 10134 7868 10140 7880
rect 1627 7840 10140 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 16500 7877 16528 7908
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17512 7945 17540 7976
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 20530 8004 20536 8016
rect 18840 7976 20536 8004
rect 18840 7964 18846 7976
rect 20530 7964 20536 7976
rect 20588 8004 20594 8016
rect 21008 8004 21036 8044
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 22462 8072 22468 8084
rect 21876 8044 22468 8072
rect 21876 8032 21882 8044
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 25590 8032 25596 8084
rect 25648 8072 25654 8084
rect 25774 8072 25780 8084
rect 25648 8044 25780 8072
rect 25648 8032 25654 8044
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 27709 8075 27767 8081
rect 27709 8072 27721 8075
rect 26108 8044 27721 8072
rect 26108 8032 26114 8044
rect 27709 8041 27721 8044
rect 27755 8041 27767 8075
rect 29825 8075 29883 8081
rect 29825 8072 29837 8075
rect 27709 8035 27767 8041
rect 27908 8044 29837 8072
rect 23750 8004 23756 8016
rect 20588 7976 21036 8004
rect 21100 7976 23756 8004
rect 20588 7964 20594 7976
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17276 7908 17417 7936
rect 17276 7896 17282 7908
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 19702 7936 19708 7948
rect 17644 7908 19708 7936
rect 17644 7896 17650 7908
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 20254 7896 20260 7948
rect 20312 7896 20318 7948
rect 20898 7896 20904 7948
rect 20956 7936 20962 7948
rect 21100 7945 21128 7976
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 27908 8004 27936 8044
rect 29825 8041 29837 8044
rect 29871 8072 29883 8075
rect 32030 8072 32036 8084
rect 29871 8044 32036 8072
rect 29871 8041 29883 8044
rect 29825 8035 29883 8041
rect 32030 8032 32036 8044
rect 32088 8032 32094 8084
rect 32950 8072 32956 8084
rect 32692 8044 32956 8072
rect 26896 7976 27936 8004
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20956 7908 21005 7936
rect 20956 7896 20962 7908
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 21726 7936 21732 7948
rect 21085 7899 21143 7905
rect 21192 7908 21732 7936
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 13044 7840 16497 7868
rect 13044 7828 13050 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 17313 7871 17371 7877
rect 17313 7868 17325 7871
rect 16724 7840 17325 7868
rect 16724 7828 16730 7840
rect 17313 7837 17325 7840
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 17954 7828 17960 7880
rect 18012 7868 18018 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 18012 7840 18153 7868
rect 18012 7828 18018 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18322 7868 18328 7880
rect 18283 7840 18328 7868
rect 18141 7831 18199 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 18598 7877 18604 7880
rect 18555 7871 18604 7877
rect 18472 7840 18517 7868
rect 18472 7828 18478 7840
rect 18555 7837 18567 7871
rect 18601 7837 18604 7871
rect 18555 7831 18604 7837
rect 18598 7828 18604 7831
rect 18656 7828 18662 7880
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 18748 7840 18920 7868
rect 18748 7828 18754 7840
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 9769 7803 9827 7809
rect 9769 7800 9781 7803
rect 9732 7772 9781 7800
rect 9732 7760 9738 7772
rect 9769 7769 9781 7772
rect 9815 7800 9827 7803
rect 10502 7800 10508 7812
rect 9815 7772 10508 7800
rect 9815 7769 9827 7772
rect 9769 7763 9827 7769
rect 10502 7760 10508 7772
rect 10560 7760 10566 7812
rect 18782 7800 18788 7812
rect 18524 7772 18788 7800
rect 17126 7692 17132 7744
rect 17184 7732 17190 7744
rect 18524 7732 18552 7772
rect 18782 7760 18788 7772
rect 18840 7760 18846 7812
rect 18892 7800 18920 7840
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19024 7840 20085 7868
rect 19024 7828 19030 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20272 7868 20300 7896
rect 20211 7840 20300 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21192 7868 21220 7908
rect 21726 7896 21732 7908
rect 21784 7936 21790 7948
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21784 7908 22017 7936
rect 21784 7896 21790 7908
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22152 7908 22508 7936
rect 22152 7896 22158 7908
rect 21450 7868 21456 7880
rect 20864 7840 21220 7868
rect 21363 7840 21456 7868
rect 20864 7828 20870 7840
rect 21450 7828 21456 7840
rect 21508 7868 21514 7880
rect 22480 7877 22508 7908
rect 22554 7896 22560 7948
rect 22612 7936 22618 7948
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 22612 7908 22845 7936
rect 22612 7896 22618 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 25130 7936 25136 7948
rect 25091 7908 25136 7936
rect 22833 7899 22891 7905
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 25222 7896 25228 7948
rect 25280 7936 25286 7948
rect 25590 7936 25596 7948
rect 25280 7908 25596 7936
rect 25280 7896 25286 7908
rect 25590 7896 25596 7908
rect 25648 7936 25654 7948
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25648 7908 25881 7936
rect 25648 7896 25654 7908
rect 25869 7905 25881 7908
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 22465 7871 22523 7877
rect 21508 7840 22416 7868
rect 21508 7828 21514 7840
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 18892 7772 19625 7800
rect 19613 7769 19625 7772
rect 19659 7800 19671 7803
rect 19978 7800 19984 7812
rect 19659 7772 19984 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 20257 7803 20315 7809
rect 20257 7769 20269 7803
rect 20303 7800 20315 7803
rect 21266 7800 21272 7812
rect 20303 7772 21272 7800
rect 20303 7769 20315 7772
rect 20257 7763 20315 7769
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21545 7803 21603 7809
rect 21545 7769 21557 7803
rect 21591 7800 21603 7803
rect 22278 7800 22284 7812
rect 21591 7772 22284 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 22388 7800 22416 7840
rect 22465 7837 22477 7871
rect 22511 7837 22523 7871
rect 24670 7868 24676 7880
rect 24631 7840 24676 7868
rect 22465 7831 22523 7837
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 26896 7868 26924 7976
rect 30282 7964 30288 8016
rect 30340 8004 30346 8016
rect 32692 8004 32720 8044
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 33686 8032 33692 8084
rect 33744 8072 33750 8084
rect 34330 8072 34336 8084
rect 33744 8044 34336 8072
rect 33744 8032 33750 8044
rect 34330 8032 34336 8044
rect 34388 8032 34394 8084
rect 35066 8032 35072 8084
rect 35124 8072 35130 8084
rect 35124 8044 35894 8072
rect 35124 8032 35130 8044
rect 30340 7976 32720 8004
rect 30340 7964 30346 7976
rect 32766 7964 32772 8016
rect 32824 8004 32830 8016
rect 32824 7976 34100 8004
rect 32824 7964 32830 7976
rect 28261 7939 28319 7945
rect 28261 7905 28273 7939
rect 28307 7936 28319 7939
rect 28626 7936 28632 7948
rect 28307 7908 28632 7936
rect 28307 7905 28319 7908
rect 28261 7899 28319 7905
rect 28626 7896 28632 7908
rect 28684 7896 28690 7948
rect 28810 7896 28816 7948
rect 28868 7936 28874 7948
rect 28868 7908 29040 7936
rect 28868 7896 28874 7908
rect 25792 7840 26924 7868
rect 22388 7772 24348 7800
rect 17184 7704 18552 7732
rect 18693 7735 18751 7741
rect 17184 7692 17190 7704
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 21726 7732 21732 7744
rect 18739 7704 21732 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 21726 7692 21732 7704
rect 21784 7732 21790 7744
rect 24210 7732 24216 7744
rect 21784 7704 24216 7732
rect 21784 7692 21790 7704
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 24320 7732 24348 7772
rect 24578 7760 24584 7812
rect 24636 7800 24642 7812
rect 25792 7800 25820 7840
rect 26970 7828 26976 7880
rect 27028 7868 27034 7880
rect 29012 7877 29040 7908
rect 29086 7896 29092 7948
rect 29144 7936 29150 7948
rect 29144 7908 31340 7936
rect 29144 7896 29150 7908
rect 30024 7877 30052 7908
rect 28169 7871 28227 7877
rect 28169 7868 28181 7871
rect 27028 7840 28181 7868
rect 27028 7828 27034 7840
rect 28169 7837 28181 7840
rect 28215 7837 28227 7871
rect 28169 7831 28227 7837
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 30009 7871 30067 7877
rect 30009 7837 30021 7871
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 30098 7828 30104 7880
rect 30156 7868 30162 7880
rect 30282 7868 30288 7880
rect 30156 7840 30201 7868
rect 30243 7840 30288 7868
rect 30156 7828 30162 7840
rect 30282 7828 30288 7840
rect 30340 7828 30346 7880
rect 30377 7871 30435 7877
rect 30377 7837 30389 7871
rect 30423 7868 30435 7871
rect 31018 7868 31024 7880
rect 30423 7840 31024 7868
rect 30423 7837 30435 7840
rect 30377 7831 30435 7837
rect 31018 7828 31024 7840
rect 31076 7828 31082 7880
rect 24636 7772 25820 7800
rect 24636 7760 24642 7772
rect 25866 7760 25872 7812
rect 25924 7800 25930 7812
rect 26114 7803 26172 7809
rect 26114 7800 26126 7803
rect 25924 7772 26126 7800
rect 25924 7760 25930 7772
rect 26114 7769 26126 7772
rect 26160 7769 26172 7803
rect 31205 7803 31263 7809
rect 31205 7800 31217 7803
rect 26114 7763 26172 7769
rect 27080 7772 27476 7800
rect 25130 7732 25136 7744
rect 24320 7704 25136 7732
rect 25130 7692 25136 7704
rect 25188 7692 25194 7744
rect 25498 7692 25504 7744
rect 25556 7732 25562 7744
rect 27080 7732 27108 7772
rect 27246 7732 27252 7744
rect 25556 7704 27108 7732
rect 27207 7704 27252 7732
rect 25556 7692 25562 7704
rect 27246 7692 27252 7704
rect 27304 7692 27310 7744
rect 27448 7732 27476 7772
rect 30116 7772 31217 7800
rect 30116 7744 30144 7772
rect 30392 7744 30420 7772
rect 31205 7769 31217 7772
rect 31251 7769 31263 7803
rect 31312 7800 31340 7908
rect 32306 7896 32312 7948
rect 32364 7936 32370 7948
rect 34072 7945 34100 7976
rect 34238 7964 34244 8016
rect 34296 8004 34302 8016
rect 35250 8004 35256 8016
rect 34296 7976 35256 8004
rect 34296 7964 34302 7976
rect 35250 7964 35256 7976
rect 35308 7964 35314 8016
rect 35342 7964 35348 8016
rect 35400 8004 35406 8016
rect 35400 7976 35577 8004
rect 35400 7964 35406 7976
rect 32953 7939 33011 7945
rect 32953 7936 32965 7939
rect 32364 7908 32965 7936
rect 32364 7896 32370 7908
rect 32953 7905 32965 7908
rect 32999 7936 33011 7939
rect 34057 7939 34115 7945
rect 32999 7908 33999 7936
rect 32999 7905 33011 7908
rect 32953 7899 33011 7905
rect 33597 7871 33655 7877
rect 33597 7837 33609 7871
rect 33643 7837 33655 7871
rect 33597 7831 33655 7837
rect 33689 7871 33747 7877
rect 33689 7837 33701 7871
rect 33735 7837 33747 7871
rect 33870 7868 33876 7880
rect 33831 7840 33876 7868
rect 33689 7831 33747 7837
rect 33042 7800 33048 7812
rect 31312 7772 33048 7800
rect 31205 7763 31263 7769
rect 33042 7760 33048 7772
rect 33100 7760 33106 7812
rect 27982 7732 27988 7744
rect 27448 7704 27988 7732
rect 27982 7692 27988 7704
rect 28040 7692 28046 7744
rect 28077 7735 28135 7741
rect 28077 7701 28089 7735
rect 28123 7732 28135 7735
rect 28902 7732 28908 7744
rect 28123 7704 28908 7732
rect 28123 7701 28135 7704
rect 28077 7695 28135 7701
rect 28902 7692 28908 7704
rect 28960 7692 28966 7744
rect 29086 7732 29092 7744
rect 29047 7704 29092 7732
rect 29086 7692 29092 7704
rect 29144 7692 29150 7744
rect 30098 7692 30104 7744
rect 30156 7692 30162 7744
rect 30374 7692 30380 7744
rect 30432 7692 30438 7744
rect 30834 7692 30840 7744
rect 30892 7732 30898 7744
rect 32766 7732 32772 7744
rect 30892 7704 32772 7732
rect 30892 7692 30898 7704
rect 32766 7692 32772 7704
rect 32824 7692 32830 7744
rect 33612 7732 33640 7831
rect 33704 7800 33732 7831
rect 33870 7828 33876 7840
rect 33928 7828 33934 7880
rect 33971 7868 33999 7908
rect 34057 7905 34069 7939
rect 34103 7905 34115 7939
rect 34057 7899 34115 7905
rect 34422 7896 34428 7948
rect 34480 7936 34486 7948
rect 34480 7908 35480 7936
rect 34480 7896 34486 7908
rect 34698 7868 34704 7880
rect 33971 7840 34704 7868
rect 34698 7828 34704 7840
rect 34756 7828 34762 7880
rect 35066 7868 35072 7880
rect 35027 7840 35072 7868
rect 35066 7828 35072 7840
rect 35124 7828 35130 7880
rect 35452 7877 35480 7908
rect 35549 7877 35577 7976
rect 35866 7936 35894 8044
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36998 8072 37004 8084
rect 36136 8044 37004 8072
rect 36136 8032 36142 8044
rect 36998 8032 37004 8044
rect 37056 8032 37062 8084
rect 37274 8032 37280 8084
rect 37332 8072 37338 8084
rect 37550 8072 37556 8084
rect 37332 8044 37556 8072
rect 37332 8032 37338 8044
rect 37550 8032 37556 8044
rect 37608 8032 37614 8084
rect 38010 8032 38016 8084
rect 38068 8072 38074 8084
rect 39117 8075 39175 8081
rect 39117 8072 39129 8075
rect 38068 8044 39129 8072
rect 38068 8032 38074 8044
rect 39117 8041 39129 8044
rect 39163 8041 39175 8075
rect 40770 8072 40776 8084
rect 40731 8044 40776 8072
rect 39117 8035 39175 8041
rect 40770 8032 40776 8044
rect 40828 8032 40834 8084
rect 41782 8032 41788 8084
rect 41840 8072 41846 8084
rect 44910 8072 44916 8084
rect 41840 8044 44916 8072
rect 41840 8032 41846 8044
rect 36173 8007 36231 8013
rect 36173 7973 36185 8007
rect 36219 8004 36231 8007
rect 36906 8004 36912 8016
rect 36219 7976 36912 8004
rect 36219 7973 36231 7976
rect 36173 7967 36231 7973
rect 36906 7964 36912 7976
rect 36964 7964 36970 8016
rect 37366 8004 37372 8016
rect 37200 7976 37372 8004
rect 36633 7939 36691 7945
rect 35866 7908 36216 7936
rect 36188 7880 36216 7908
rect 36633 7905 36645 7939
rect 36679 7936 36691 7939
rect 36722 7936 36728 7948
rect 36679 7908 36728 7936
rect 36679 7905 36691 7908
rect 36633 7899 36691 7905
rect 36722 7896 36728 7908
rect 36780 7896 36786 7948
rect 36817 7939 36875 7945
rect 36817 7905 36829 7939
rect 36863 7936 36875 7939
rect 37200 7936 37228 7976
rect 37366 7964 37372 7976
rect 37424 7964 37430 8016
rect 37642 7964 37648 8016
rect 37700 8004 37706 8016
rect 37700 7976 40264 8004
rect 37700 7964 37706 7976
rect 39850 7936 39856 7948
rect 36863 7908 37228 7936
rect 37292 7908 39856 7936
rect 36863 7905 36875 7908
rect 36817 7899 36875 7905
rect 35217 7871 35275 7877
rect 35217 7837 35229 7871
rect 35263 7837 35275 7871
rect 35217 7831 35275 7837
rect 35437 7871 35495 7877
rect 35437 7837 35449 7871
rect 35483 7837 35495 7871
rect 35437 7831 35495 7837
rect 35534 7871 35592 7877
rect 35534 7837 35546 7871
rect 35580 7837 35592 7871
rect 35534 7831 35592 7837
rect 34146 7800 34152 7812
rect 33704 7772 34152 7800
rect 34146 7760 34152 7772
rect 34204 7760 34210 7812
rect 34514 7732 34520 7744
rect 33612 7704 34520 7732
rect 34514 7692 34520 7704
rect 34572 7692 34578 7744
rect 35232 7732 35260 7831
rect 36170 7828 36176 7880
rect 36228 7828 36234 7880
rect 37292 7868 37320 7908
rect 39850 7896 39856 7908
rect 39908 7896 39914 7948
rect 36280 7840 37320 7868
rect 37461 7871 37519 7877
rect 35342 7760 35348 7812
rect 35400 7800 35406 7812
rect 36280 7800 36308 7840
rect 37461 7837 37473 7871
rect 37507 7868 37519 7871
rect 37734 7868 37740 7880
rect 37507 7840 37740 7868
rect 37507 7837 37519 7840
rect 37461 7831 37519 7837
rect 37734 7828 37740 7840
rect 37792 7868 37798 7880
rect 38378 7868 38384 7880
rect 37792 7840 38384 7868
rect 37792 7828 37798 7840
rect 38378 7828 38384 7840
rect 38436 7828 38442 7880
rect 38470 7828 38476 7880
rect 38528 7868 38534 7880
rect 38565 7871 38623 7877
rect 38565 7868 38577 7871
rect 38528 7840 38577 7868
rect 38528 7828 38534 7840
rect 38565 7837 38577 7840
rect 38611 7837 38623 7871
rect 38746 7868 38752 7880
rect 38707 7840 38752 7868
rect 38565 7831 38623 7837
rect 38746 7828 38752 7840
rect 38804 7828 38810 7880
rect 38933 7871 38991 7877
rect 38933 7837 38945 7871
rect 38979 7868 38991 7871
rect 39114 7868 39120 7880
rect 38979 7840 39120 7868
rect 38979 7837 38991 7840
rect 38933 7831 38991 7837
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39390 7828 39396 7880
rect 39448 7868 39454 7880
rect 40025 7871 40083 7877
rect 39448 7840 39988 7868
rect 39448 7828 39454 7840
rect 35400 7772 35445 7800
rect 35544 7772 36308 7800
rect 36541 7803 36599 7809
rect 35400 7760 35406 7772
rect 35544 7732 35572 7772
rect 36541 7769 36553 7803
rect 36587 7800 36599 7803
rect 37274 7800 37280 7812
rect 36587 7772 37280 7800
rect 36587 7769 36599 7772
rect 36541 7763 36599 7769
rect 37274 7760 37280 7772
rect 37332 7760 37338 7812
rect 37366 7760 37372 7812
rect 37424 7800 37430 7812
rect 37829 7803 37887 7809
rect 37829 7800 37841 7803
rect 37424 7772 37841 7800
rect 37424 7760 37430 7772
rect 37829 7769 37841 7772
rect 37875 7769 37887 7803
rect 37829 7763 37887 7769
rect 38841 7803 38899 7809
rect 38841 7769 38853 7803
rect 38887 7800 38899 7803
rect 39758 7800 39764 7812
rect 38887 7772 39764 7800
rect 38887 7769 38899 7772
rect 38841 7763 38899 7769
rect 39758 7760 39764 7772
rect 39816 7760 39822 7812
rect 39960 7800 39988 7840
rect 40025 7837 40037 7871
rect 40071 7868 40083 7871
rect 40126 7868 40132 7880
rect 40071 7840 40132 7868
rect 40071 7837 40083 7840
rect 40025 7831 40083 7837
rect 40126 7828 40132 7840
rect 40184 7828 40190 7880
rect 40236 7877 40264 7976
rect 42242 7936 42248 7948
rect 42076 7908 42248 7936
rect 40221 7871 40279 7877
rect 40221 7837 40233 7871
rect 40267 7837 40279 7871
rect 40221 7831 40279 7837
rect 40681 7871 40739 7877
rect 40681 7837 40693 7871
rect 40727 7837 40739 7871
rect 40681 7831 40739 7837
rect 40696 7800 40724 7831
rect 41690 7828 41696 7880
rect 41748 7868 41754 7880
rect 42076 7877 42104 7908
rect 42242 7896 42248 7908
rect 42300 7896 42306 7948
rect 41923 7871 41981 7877
rect 41923 7868 41935 7871
rect 41748 7840 41935 7868
rect 41748 7828 41754 7840
rect 41923 7837 41935 7840
rect 41969 7837 41981 7871
rect 41923 7831 41981 7837
rect 42058 7871 42116 7877
rect 42058 7837 42070 7871
rect 42104 7837 42116 7871
rect 42058 7831 42116 7837
rect 42150 7828 42156 7880
rect 42208 7877 42214 7880
rect 42352 7877 42380 8044
rect 44910 8032 44916 8044
rect 44968 8032 44974 8084
rect 58250 8072 58256 8084
rect 58211 8044 58256 8072
rect 58250 8032 58256 8044
rect 58308 8032 58314 8084
rect 56137 8007 56195 8013
rect 56137 7973 56149 8007
rect 56183 7973 56195 8007
rect 56137 7967 56195 7973
rect 56152 7936 56180 7967
rect 56870 7936 56876 7948
rect 56152 7908 56640 7936
rect 56831 7908 56876 7936
rect 42208 7868 42216 7877
rect 42337 7871 42395 7877
rect 42208 7840 42253 7868
rect 42208 7831 42216 7840
rect 42337 7837 42349 7871
rect 42383 7837 42395 7871
rect 42337 7831 42395 7837
rect 42208 7828 42214 7831
rect 42702 7828 42708 7880
rect 42760 7868 42766 7880
rect 42797 7871 42855 7877
rect 42797 7868 42809 7871
rect 42760 7840 42809 7868
rect 42760 7828 42766 7840
rect 42797 7837 42809 7840
rect 42843 7868 42855 7871
rect 45462 7868 45468 7880
rect 42843 7840 45468 7868
rect 42843 7837 42855 7840
rect 42797 7831 42855 7837
rect 45462 7828 45468 7840
rect 45520 7828 45526 7880
rect 49694 7828 49700 7880
rect 49752 7868 49758 7880
rect 56413 7871 56471 7877
rect 56413 7868 56425 7871
rect 49752 7840 56425 7868
rect 49752 7828 49758 7840
rect 56413 7837 56425 7840
rect 56459 7837 56471 7871
rect 56612 7868 56640 7908
rect 56870 7896 56876 7908
rect 56928 7896 56934 7948
rect 57129 7871 57187 7877
rect 57129 7868 57141 7871
rect 56612 7840 57141 7868
rect 56413 7831 56471 7837
rect 57129 7837 57141 7840
rect 57175 7837 57187 7871
rect 57129 7831 57187 7837
rect 43042 7803 43100 7809
rect 43042 7800 43054 7803
rect 39960 7772 40724 7800
rect 42168 7772 43054 7800
rect 35232 7704 35572 7732
rect 35713 7735 35771 7741
rect 35713 7701 35725 7735
rect 35759 7732 35771 7735
rect 36998 7732 37004 7744
rect 35759 7704 37004 7732
rect 35759 7701 35771 7704
rect 35713 7695 35771 7701
rect 36998 7692 37004 7704
rect 37056 7692 37062 7744
rect 37550 7692 37556 7744
rect 37608 7732 37614 7744
rect 40129 7735 40187 7741
rect 40129 7732 40141 7735
rect 37608 7704 40141 7732
rect 37608 7692 37614 7704
rect 40129 7701 40141 7704
rect 40175 7701 40187 7735
rect 40129 7695 40187 7701
rect 41693 7735 41751 7741
rect 41693 7701 41705 7735
rect 41739 7732 41751 7735
rect 42168 7732 42196 7772
rect 43042 7769 43054 7772
rect 43088 7769 43100 7803
rect 43042 7763 43100 7769
rect 44266 7760 44272 7812
rect 44324 7800 44330 7812
rect 56134 7800 56140 7812
rect 44324 7772 56140 7800
rect 44324 7760 44330 7772
rect 56134 7760 56140 7772
rect 56192 7760 56198 7812
rect 56321 7803 56379 7809
rect 56321 7769 56333 7803
rect 56367 7800 56379 7803
rect 56594 7800 56600 7812
rect 56367 7772 56600 7800
rect 56367 7769 56379 7772
rect 56321 7763 56379 7769
rect 56594 7760 56600 7772
rect 56652 7760 56658 7812
rect 44174 7732 44180 7744
rect 41739 7704 42196 7732
rect 44135 7704 44180 7732
rect 41739 7701 41751 7704
rect 41693 7695 41751 7701
rect 44174 7692 44180 7704
rect 44232 7692 44238 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 18690 7528 18696 7540
rect 9692 7500 18696 7528
rect 8662 7460 8668 7472
rect 8623 7432 8668 7460
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 9692 7469 9720 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 20898 7528 20904 7540
rect 19392 7500 20904 7528
rect 19392 7488 19398 7500
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21542 7528 21548 7540
rect 21140 7500 21548 7528
rect 21140 7488 21146 7500
rect 21542 7488 21548 7500
rect 21600 7488 21606 7540
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22738 7528 22744 7540
rect 22336 7500 22744 7528
rect 22336 7488 22342 7500
rect 22738 7488 22744 7500
rect 22796 7528 22802 7540
rect 23106 7528 23112 7540
rect 22796 7500 23112 7528
rect 22796 7488 22802 7500
rect 23106 7488 23112 7500
rect 23164 7528 23170 7540
rect 23293 7531 23351 7537
rect 23293 7528 23305 7531
rect 23164 7500 23305 7528
rect 23164 7488 23170 7500
rect 23293 7497 23305 7500
rect 23339 7497 23351 7531
rect 25866 7528 25872 7540
rect 25827 7500 25872 7528
rect 23293 7491 23351 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 26510 7528 26516 7540
rect 26283 7500 26516 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 26510 7488 26516 7500
rect 26568 7488 26574 7540
rect 26694 7488 26700 7540
rect 26752 7528 26758 7540
rect 31110 7528 31116 7540
rect 26752 7500 30512 7528
rect 31071 7500 31116 7528
rect 26752 7488 26758 7500
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7429 9735 7463
rect 26329 7463 26387 7469
rect 26329 7460 26341 7463
rect 9677 7423 9735 7429
rect 12406 7432 26341 7460
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8251 7364 9352 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 7064 7296 7941 7324
rect 7064 7284 7070 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 8036 7256 8064 7355
rect 9324 7324 9352 7364
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 10318 7392 10324 7404
rect 9456 7364 9501 7392
rect 10279 7364 10324 7392
rect 9456 7352 9462 7364
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 12406 7392 12434 7432
rect 26329 7429 26341 7432
rect 26375 7460 26387 7463
rect 27246 7460 27252 7472
rect 26375 7432 27252 7460
rect 26375 7429 26387 7432
rect 26329 7423 26387 7429
rect 27246 7420 27252 7432
rect 27304 7420 27310 7472
rect 28629 7463 28687 7469
rect 28629 7429 28641 7463
rect 28675 7460 28687 7463
rect 30098 7460 30104 7472
rect 28675 7432 30104 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 30098 7420 30104 7432
rect 30156 7420 30162 7472
rect 30484 7460 30512 7500
rect 31110 7488 31116 7500
rect 31168 7488 31174 7540
rect 31297 7531 31355 7537
rect 31297 7497 31309 7531
rect 31343 7497 31355 7531
rect 32674 7528 32680 7540
rect 32635 7500 32680 7528
rect 31297 7491 31355 7497
rect 31312 7460 31340 7491
rect 32674 7488 32680 7500
rect 32732 7528 32738 7540
rect 33778 7528 33784 7540
rect 32732 7500 33784 7528
rect 32732 7488 32738 7500
rect 33778 7488 33784 7500
rect 33836 7488 33842 7540
rect 34057 7531 34115 7537
rect 34057 7497 34069 7531
rect 34103 7528 34115 7531
rect 35894 7528 35900 7540
rect 34103 7500 35900 7528
rect 34103 7497 34115 7500
rect 34057 7491 34115 7497
rect 35894 7488 35900 7500
rect 35952 7488 35958 7540
rect 36078 7488 36084 7540
rect 36136 7488 36142 7540
rect 36906 7488 36912 7540
rect 36964 7528 36970 7540
rect 41693 7531 41751 7537
rect 36964 7500 38792 7528
rect 36964 7488 36970 7500
rect 33134 7460 33140 7472
rect 30484 7432 31340 7460
rect 31496 7432 33140 7460
rect 10459 7364 12434 7392
rect 17037 7395 17095 7401
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17313 7395 17371 7401
rect 17083 7364 17264 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 9674 7324 9680 7336
rect 9324 7296 9680 7324
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 10134 7324 10140 7336
rect 10095 7296 10140 7324
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10502 7324 10508 7336
rect 10463 7296 10508 7324
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 17126 7324 17132 7336
rect 10652 7296 10697 7324
rect 17087 7296 17132 7324
rect 10652 7284 10658 7296
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 17236 7256 17264 7364
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17359 7364 17877 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 17865 7361 17877 7364
rect 17911 7392 17923 7395
rect 19334 7392 19340 7404
rect 17911 7364 19340 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7392 19763 7395
rect 19794 7392 19800 7404
rect 19751 7364 19800 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18141 7327 18199 7333
rect 18141 7324 18153 7327
rect 18104 7296 18153 7324
rect 18104 7284 18110 7296
rect 18141 7293 18153 7296
rect 18187 7324 18199 7327
rect 18966 7324 18972 7336
rect 18187 7296 18972 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19628 7324 19656 7355
rect 19794 7352 19800 7364
rect 19852 7392 19858 7404
rect 20254 7392 20260 7404
rect 19852 7364 20260 7392
rect 19852 7352 19858 7364
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 22002 7392 22008 7404
rect 20956 7364 21001 7392
rect 21284 7364 22008 7392
rect 20956 7352 20962 7364
rect 19199 7296 19334 7324
rect 19628 7296 19748 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 18322 7256 18328 7268
rect 8036 7228 12434 7256
rect 17236 7228 18328 7256
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8904 7160 9229 7188
rect 8904 7148 8910 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 12406 7188 12434 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 18598 7216 18604 7268
rect 18656 7256 18662 7268
rect 19058 7256 19064 7268
rect 18656 7228 19064 7256
rect 18656 7216 18662 7228
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 19306 7256 19334 7296
rect 19720 7256 19748 7296
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 19944 7296 20361 7324
rect 19944 7284 19950 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7324 20499 7327
rect 21284 7324 21312 7364
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7361 24731 7395
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 24673 7355 24731 7361
rect 24835 7364 27169 7392
rect 20487 7296 21312 7324
rect 20487 7293 20499 7296
rect 20441 7287 20499 7293
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 21416 7296 21461 7324
rect 21416 7284 21422 7296
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 24578 7324 24584 7336
rect 21600 7296 24584 7324
rect 21600 7284 21606 7296
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 20254 7256 20260 7268
rect 19306 7228 19656 7256
rect 19720 7228 20260 7256
rect 15470 7188 15476 7200
rect 12406 7160 15476 7188
rect 9217 7151 9275 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 17221 7191 17279 7197
rect 17221 7157 17233 7191
rect 17267 7188 17279 7191
rect 19518 7188 19524 7200
rect 17267 7160 19524 7188
rect 17267 7157 17279 7160
rect 17221 7151 17279 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19628 7188 19656 7228
rect 20254 7216 20260 7228
rect 20312 7216 20318 7268
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 21450 7256 21456 7268
rect 20772 7228 21456 7256
rect 20772 7216 20778 7228
rect 21450 7216 21456 7228
rect 21508 7256 21514 7268
rect 24688 7256 24716 7355
rect 21508 7228 24716 7256
rect 21508 7216 21514 7228
rect 22186 7188 22192 7200
rect 19628 7160 22192 7188
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 24210 7148 24216 7200
rect 24268 7188 24274 7200
rect 24835 7197 24863 7364
rect 27157 7361 27169 7364
rect 27203 7361 27215 7395
rect 31294 7395 31352 7401
rect 27157 7355 27215 7361
rect 27356 7364 27660 7392
rect 24946 7284 24952 7336
rect 25004 7324 25010 7336
rect 25041 7327 25099 7333
rect 25041 7324 25053 7327
rect 25004 7296 25053 7324
rect 25004 7284 25010 7296
rect 25041 7293 25053 7296
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 25409 7327 25467 7333
rect 25409 7293 25421 7327
rect 25455 7324 25467 7327
rect 25774 7324 25780 7336
rect 25455 7296 25780 7324
rect 25455 7293 25467 7296
rect 25409 7287 25467 7293
rect 25774 7284 25780 7296
rect 25832 7284 25838 7336
rect 26513 7327 26571 7333
rect 26513 7293 26525 7327
rect 26559 7324 26571 7327
rect 27356 7324 27384 7364
rect 27522 7324 27528 7336
rect 26559 7296 27384 7324
rect 27483 7296 27528 7324
rect 26559 7293 26571 7296
rect 26513 7287 26571 7293
rect 27522 7284 27528 7296
rect 27580 7284 27586 7336
rect 27632 7324 27660 7364
rect 31294 7361 31306 7395
rect 31340 7392 31352 7395
rect 31496 7392 31524 7432
rect 33134 7420 33140 7432
rect 33192 7420 33198 7472
rect 34698 7420 34704 7472
rect 34756 7460 34762 7472
rect 35434 7460 35440 7472
rect 34756 7432 35204 7460
rect 35395 7432 35440 7460
rect 34756 7420 34762 7432
rect 31340 7364 31524 7392
rect 31757 7395 31815 7401
rect 31340 7361 31352 7364
rect 31294 7355 31352 7361
rect 31757 7361 31769 7395
rect 31803 7392 31815 7395
rect 32030 7392 32036 7404
rect 31803 7364 32036 7392
rect 31803 7361 31815 7364
rect 31757 7355 31815 7361
rect 32030 7352 32036 7364
rect 32088 7352 32094 7404
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 35176 7401 35204 7432
rect 35434 7420 35440 7432
rect 35492 7420 35498 7472
rect 35069 7395 35127 7401
rect 35069 7392 35081 7395
rect 34296 7364 35081 7392
rect 34296 7352 34302 7364
rect 35069 7361 35081 7364
rect 35115 7361 35127 7395
rect 35069 7355 35127 7361
rect 35162 7395 35220 7401
rect 35162 7361 35174 7395
rect 35208 7361 35220 7395
rect 35162 7355 35220 7361
rect 35250 7352 35256 7404
rect 35308 7392 35314 7404
rect 35345 7395 35403 7401
rect 35345 7392 35357 7395
rect 35308 7364 35357 7392
rect 35308 7352 35314 7364
rect 35345 7361 35357 7364
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 35534 7395 35592 7401
rect 35534 7361 35546 7395
rect 35580 7392 35592 7395
rect 35580 7364 35756 7392
rect 35580 7361 35592 7364
rect 35534 7355 35592 7361
rect 28626 7324 28632 7336
rect 27632 7296 28632 7324
rect 28626 7284 28632 7296
rect 28684 7284 28690 7336
rect 32582 7284 32588 7336
rect 32640 7324 32646 7336
rect 32769 7327 32827 7333
rect 32769 7324 32781 7327
rect 32640 7296 32781 7324
rect 32640 7284 32646 7296
rect 32769 7293 32781 7296
rect 32815 7293 32827 7327
rect 32769 7287 32827 7293
rect 32861 7327 32919 7333
rect 32861 7293 32873 7327
rect 32907 7293 32919 7327
rect 32861 7287 32919 7293
rect 33873 7327 33931 7333
rect 33873 7293 33885 7327
rect 33919 7293 33931 7327
rect 34330 7324 34336 7336
rect 34291 7296 34336 7324
rect 33873 7287 33931 7293
rect 25222 7216 25228 7268
rect 25280 7256 25286 7268
rect 27433 7259 27491 7265
rect 27433 7256 27445 7259
rect 25280 7228 27445 7256
rect 25280 7216 25286 7228
rect 27433 7225 27445 7228
rect 27479 7225 27491 7259
rect 27433 7219 27491 7225
rect 27614 7216 27620 7268
rect 27672 7256 27678 7268
rect 29270 7256 29276 7268
rect 27672 7228 29276 7256
rect 27672 7216 27678 7228
rect 29270 7216 29276 7228
rect 29328 7216 29334 7268
rect 31018 7216 31024 7268
rect 31076 7256 31082 7268
rect 31076 7228 32444 7256
rect 31076 7216 31082 7228
rect 24835 7191 24896 7197
rect 24835 7188 24850 7191
rect 24268 7160 24850 7188
rect 24268 7148 24274 7160
rect 24838 7157 24850 7160
rect 24884 7157 24896 7191
rect 24838 7151 24896 7157
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25038 7188 25044 7200
rect 24995 7160 25044 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25038 7148 25044 7160
rect 25096 7188 25102 7200
rect 27295 7191 27353 7197
rect 27295 7188 27307 7191
rect 25096 7160 27307 7188
rect 25096 7148 25102 7160
rect 27295 7157 27307 7160
rect 27341 7157 27353 7191
rect 27295 7151 27353 7157
rect 27801 7191 27859 7197
rect 27801 7157 27813 7191
rect 27847 7188 27859 7191
rect 28258 7188 28264 7200
rect 27847 7160 28264 7188
rect 27847 7157 27859 7160
rect 27801 7151 27859 7157
rect 28258 7148 28264 7160
rect 28316 7188 28322 7200
rect 28810 7188 28816 7200
rect 28316 7160 28816 7188
rect 28316 7148 28322 7160
rect 28810 7148 28816 7160
rect 28868 7148 28874 7200
rect 29546 7148 29552 7200
rect 29604 7188 29610 7200
rect 29917 7191 29975 7197
rect 29917 7188 29929 7191
rect 29604 7160 29929 7188
rect 29604 7148 29610 7160
rect 29917 7157 29929 7160
rect 29963 7188 29975 7191
rect 30742 7188 30748 7200
rect 29963 7160 30748 7188
rect 29963 7157 29975 7160
rect 29917 7151 29975 7157
rect 30742 7148 30748 7160
rect 30800 7148 30806 7200
rect 31202 7148 31208 7200
rect 31260 7188 31266 7200
rect 31478 7188 31484 7200
rect 31260 7160 31484 7188
rect 31260 7148 31266 7160
rect 31478 7148 31484 7160
rect 31536 7188 31542 7200
rect 31665 7191 31723 7197
rect 31665 7188 31677 7191
rect 31536 7160 31677 7188
rect 31536 7148 31542 7160
rect 31665 7157 31677 7160
rect 31711 7157 31723 7191
rect 31665 7151 31723 7157
rect 31754 7148 31760 7200
rect 31812 7188 31818 7200
rect 32309 7191 32367 7197
rect 32309 7188 32321 7191
rect 31812 7160 32321 7188
rect 31812 7148 31818 7160
rect 32309 7157 32321 7160
rect 32355 7157 32367 7191
rect 32416 7188 32444 7228
rect 32674 7216 32680 7268
rect 32732 7256 32738 7268
rect 32876 7256 32904 7287
rect 32732 7228 32904 7256
rect 32732 7216 32738 7228
rect 33134 7216 33140 7268
rect 33192 7256 33198 7268
rect 33594 7256 33600 7268
rect 33192 7228 33600 7256
rect 33192 7216 33198 7228
rect 33594 7216 33600 7228
rect 33652 7216 33658 7268
rect 33888 7256 33916 7287
rect 34330 7284 34336 7296
rect 34388 7284 34394 7336
rect 34422 7284 34428 7336
rect 34480 7324 34486 7336
rect 35728 7324 35756 7364
rect 35802 7352 35808 7404
rect 35860 7392 35866 7404
rect 36096 7398 36124 7488
rect 36998 7420 37004 7472
rect 37056 7460 37062 7472
rect 37056 7432 37964 7460
rect 37056 7420 37062 7432
rect 36161 7401 36219 7407
rect 36161 7398 36173 7401
rect 35860 7364 36032 7392
rect 36096 7370 36173 7398
rect 35860 7352 35866 7364
rect 36004 7336 36032 7364
rect 36161 7367 36173 7370
rect 36207 7367 36219 7401
rect 36161 7361 36219 7367
rect 36449 7395 36507 7401
rect 36449 7361 36461 7395
rect 36495 7392 36507 7395
rect 37274 7392 37280 7404
rect 36495 7364 37280 7392
rect 36495 7361 36507 7364
rect 36449 7355 36507 7361
rect 37274 7352 37280 7364
rect 37332 7352 37338 7404
rect 37458 7392 37464 7404
rect 37419 7364 37464 7392
rect 37458 7352 37464 7364
rect 37516 7352 37522 7404
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7392 37703 7395
rect 37734 7392 37740 7404
rect 37691 7364 37740 7392
rect 37691 7361 37703 7364
rect 37645 7355 37703 7361
rect 37734 7352 37740 7364
rect 37792 7352 37798 7404
rect 37936 7401 37964 7432
rect 38028 7432 38654 7460
rect 37921 7395 37979 7401
rect 37921 7361 37933 7395
rect 37967 7361 37979 7395
rect 37921 7355 37979 7361
rect 34480 7296 34525 7324
rect 35728 7296 35940 7324
rect 34480 7284 34486 7296
rect 35713 7259 35771 7265
rect 35713 7256 35725 7259
rect 33888 7228 35725 7256
rect 35713 7225 35725 7228
rect 35759 7225 35771 7259
rect 35912 7256 35940 7296
rect 35986 7284 35992 7336
rect 36044 7324 36050 7336
rect 36633 7327 36691 7333
rect 36633 7324 36645 7327
rect 36044 7296 36645 7324
rect 36044 7284 36050 7296
rect 36633 7293 36645 7296
rect 36679 7293 36691 7327
rect 36633 7287 36691 7293
rect 37182 7284 37188 7336
rect 37240 7324 37246 7336
rect 37826 7324 37832 7336
rect 37240 7296 37832 7324
rect 37240 7284 37246 7296
rect 37826 7284 37832 7296
rect 37884 7284 37890 7336
rect 36078 7256 36084 7268
rect 35912 7228 36084 7256
rect 35713 7219 35771 7225
rect 36078 7216 36084 7228
rect 36136 7216 36142 7268
rect 36262 7256 36268 7268
rect 36223 7228 36268 7256
rect 36262 7216 36268 7228
rect 36320 7216 36326 7268
rect 36998 7216 37004 7268
rect 37056 7256 37062 7268
rect 37737 7259 37795 7265
rect 37737 7256 37749 7259
rect 37056 7228 37749 7256
rect 37056 7216 37062 7228
rect 37737 7225 37749 7228
rect 37783 7256 37795 7259
rect 38028 7256 38056 7432
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7392 38163 7395
rect 38194 7392 38200 7404
rect 38151 7364 38200 7392
rect 38151 7361 38163 7364
rect 38105 7355 38163 7361
rect 38194 7352 38200 7364
rect 38252 7352 38258 7404
rect 38626 7392 38654 7432
rect 38764 7401 38792 7500
rect 41693 7497 41705 7531
rect 41739 7528 41751 7531
rect 42610 7528 42616 7540
rect 41739 7500 42616 7528
rect 41739 7497 41751 7500
rect 41693 7491 41751 7497
rect 42610 7488 42616 7500
rect 42668 7488 42674 7540
rect 42705 7531 42763 7537
rect 42705 7497 42717 7531
rect 42751 7528 42763 7531
rect 43622 7528 43628 7540
rect 42751 7500 43628 7528
rect 42751 7497 42763 7500
rect 42705 7491 42763 7497
rect 43622 7488 43628 7500
rect 43680 7488 43686 7540
rect 44453 7531 44511 7537
rect 44453 7528 44465 7531
rect 43732 7500 44465 7528
rect 38933 7463 38991 7469
rect 38933 7429 38945 7463
rect 38979 7460 38991 7463
rect 39114 7460 39120 7472
rect 38979 7432 39120 7460
rect 38979 7429 38991 7432
rect 38933 7423 38991 7429
rect 39114 7420 39120 7432
rect 39172 7420 39178 7472
rect 42150 7420 42156 7472
rect 42208 7460 42214 7472
rect 43732 7460 43760 7500
rect 44453 7497 44465 7500
rect 44499 7497 44511 7531
rect 44453 7491 44511 7497
rect 55214 7488 55220 7540
rect 55272 7528 55278 7540
rect 55398 7528 55404 7540
rect 55272 7500 55404 7528
rect 55272 7488 55278 7500
rect 55398 7488 55404 7500
rect 55456 7488 55462 7540
rect 57238 7488 57244 7540
rect 57296 7528 57302 7540
rect 57296 7500 58204 7528
rect 57296 7488 57302 7500
rect 42208 7432 43760 7460
rect 42208 7420 42214 7432
rect 43898 7420 43904 7472
rect 43956 7420 43962 7472
rect 44174 7420 44180 7472
rect 44232 7460 44238 7472
rect 51074 7460 51080 7472
rect 44232 7432 51080 7460
rect 44232 7420 44238 7432
rect 38749 7395 38807 7401
rect 38626 7364 38700 7392
rect 38286 7284 38292 7336
rect 38344 7324 38350 7336
rect 38565 7327 38623 7333
rect 38565 7324 38577 7327
rect 38344 7296 38577 7324
rect 38344 7284 38350 7296
rect 38565 7293 38577 7296
rect 38611 7293 38623 7327
rect 38672 7324 38700 7364
rect 38749 7361 38761 7395
rect 38795 7361 38807 7395
rect 40126 7392 40132 7404
rect 38948 7382 40132 7392
rect 38749 7355 38807 7361
rect 38856 7364 40132 7382
rect 38856 7354 38976 7364
rect 38856 7324 38884 7354
rect 40126 7352 40132 7364
rect 40184 7352 40190 7404
rect 41598 7392 41604 7404
rect 41559 7364 41604 7392
rect 41598 7352 41604 7364
rect 41656 7352 41662 7404
rect 41782 7352 41788 7404
rect 41840 7392 41846 7404
rect 42613 7395 42671 7401
rect 41840 7364 41885 7392
rect 41840 7352 41846 7364
rect 42613 7361 42625 7395
rect 42659 7361 42671 7395
rect 42613 7355 42671 7361
rect 41969 7327 42027 7333
rect 41969 7324 41981 7327
rect 38672 7296 38884 7324
rect 38948 7296 41981 7324
rect 38565 7287 38623 7293
rect 37783 7228 38056 7256
rect 37783 7225 37795 7228
rect 37737 7219 37795 7225
rect 38378 7216 38384 7268
rect 38436 7256 38442 7268
rect 38948 7256 38976 7296
rect 41969 7293 41981 7296
rect 42015 7293 42027 7327
rect 41969 7287 42027 7293
rect 38436 7228 38976 7256
rect 38436 7216 38442 7228
rect 40402 7216 40408 7268
rect 40460 7256 40466 7268
rect 41417 7259 41475 7265
rect 41417 7256 41429 7259
rect 40460 7228 41429 7256
rect 40460 7216 40466 7228
rect 41417 7225 41429 7228
rect 41463 7256 41475 7259
rect 42058 7256 42064 7268
rect 41463 7228 42064 7256
rect 41463 7225 41475 7228
rect 41417 7219 41475 7225
rect 42058 7216 42064 7228
rect 42116 7216 42122 7268
rect 42628 7256 42656 7355
rect 42702 7352 42708 7404
rect 42760 7392 42766 7404
rect 42797 7395 42855 7401
rect 42797 7392 42809 7395
rect 42760 7364 42809 7392
rect 42760 7352 42766 7364
rect 42797 7361 42809 7364
rect 42843 7392 42855 7395
rect 42886 7392 42892 7404
rect 42843 7364 42892 7392
rect 42843 7361 42855 7364
rect 42797 7355 42855 7361
rect 42886 7352 42892 7364
rect 42944 7352 42950 7404
rect 43349 7395 43407 7401
rect 43349 7361 43361 7395
rect 43395 7392 43407 7395
rect 43916 7392 43944 7420
rect 44652 7401 44680 7432
rect 51074 7420 51080 7432
rect 51132 7420 51138 7472
rect 56134 7420 56140 7472
rect 56192 7460 56198 7472
rect 56321 7463 56379 7469
rect 56321 7460 56333 7463
rect 56192 7432 56333 7460
rect 56192 7420 56198 7432
rect 56321 7429 56333 7432
rect 56367 7429 56379 7463
rect 56321 7423 56379 7429
rect 56505 7463 56563 7469
rect 56505 7429 56517 7463
rect 56551 7460 56563 7463
rect 56551 7432 57008 7460
rect 56551 7429 56563 7432
rect 56505 7423 56563 7429
rect 43395 7364 43944 7392
rect 44637 7395 44695 7401
rect 43395 7361 43407 7364
rect 43349 7355 43407 7361
rect 44637 7361 44649 7395
rect 44683 7361 44695 7395
rect 44818 7392 44824 7404
rect 44779 7364 44824 7392
rect 44637 7355 44695 7361
rect 44818 7352 44824 7364
rect 44876 7352 44882 7404
rect 44913 7395 44971 7401
rect 44913 7361 44925 7395
rect 44959 7361 44971 7395
rect 44913 7355 44971 7361
rect 56597 7395 56655 7401
rect 56597 7361 56609 7395
rect 56643 7361 56655 7395
rect 56597 7355 56655 7361
rect 43254 7284 43260 7336
rect 43312 7324 43318 7336
rect 43625 7327 43683 7333
rect 43625 7324 43637 7327
rect 43312 7296 43637 7324
rect 43312 7284 43318 7296
rect 43625 7293 43637 7296
rect 43671 7293 43683 7327
rect 43625 7287 43683 7293
rect 42794 7256 42800 7268
rect 42628 7228 42800 7256
rect 42794 7216 42800 7228
rect 42852 7256 42858 7268
rect 44928 7256 44956 7355
rect 53926 7284 53932 7336
rect 53984 7324 53990 7336
rect 56612 7324 56640 7355
rect 53984 7296 56640 7324
rect 53984 7284 53990 7296
rect 42852 7228 44956 7256
rect 56980 7256 57008 7432
rect 57057 7395 57115 7401
rect 57057 7361 57069 7395
rect 57103 7392 57115 7395
rect 58069 7398 58127 7401
rect 58176 7398 58204 7500
rect 58069 7395 58204 7398
rect 57103 7364 57974 7392
rect 57103 7361 57115 7364
rect 57057 7355 57115 7361
rect 57330 7324 57336 7336
rect 57291 7296 57336 7324
rect 57330 7284 57336 7296
rect 57388 7284 57394 7336
rect 57946 7324 57974 7364
rect 58069 7361 58081 7395
rect 58115 7370 58204 7395
rect 58115 7361 58127 7370
rect 58069 7355 58127 7361
rect 58250 7352 58256 7404
rect 58308 7392 58314 7404
rect 58308 7364 58388 7392
rect 58308 7352 58314 7364
rect 58360 7324 58388 7364
rect 57946 7296 58388 7324
rect 58161 7259 58219 7265
rect 58161 7256 58173 7259
rect 56980 7228 58173 7256
rect 42852 7216 42858 7228
rect 58161 7225 58173 7228
rect 58207 7225 58219 7259
rect 58161 7219 58219 7225
rect 39206 7188 39212 7200
rect 32416 7160 39212 7188
rect 32309 7151 32367 7157
rect 39206 7148 39212 7160
rect 39264 7148 39270 7200
rect 42886 7148 42892 7200
rect 42944 7188 42950 7200
rect 44818 7188 44824 7200
rect 42944 7160 44824 7188
rect 42944 7148 42950 7160
rect 44818 7148 44824 7160
rect 44876 7148 44882 7200
rect 56321 7191 56379 7197
rect 56321 7157 56333 7191
rect 56367 7188 56379 7191
rect 56778 7188 56784 7200
rect 56367 7160 56784 7188
rect 56367 7157 56379 7160
rect 56321 7151 56379 7157
rect 56778 7148 56784 7160
rect 56836 7148 56842 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10560 6956 10885 6984
rect 10560 6944 10566 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 17586 6984 17592 6996
rect 17547 6956 17592 6984
rect 10873 6947 10931 6953
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 14550 6876 14556 6928
rect 14608 6916 14614 6928
rect 18892 6916 18920 6947
rect 19288 6944 19294 6996
rect 19346 6984 19352 6996
rect 19426 6984 19432 6996
rect 19346 6956 19432 6984
rect 19346 6944 19352 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 22922 6984 22928 6996
rect 19576 6956 22928 6984
rect 19576 6944 19582 6956
rect 22922 6944 22928 6956
rect 22980 6984 22986 6996
rect 22980 6956 23244 6984
rect 22980 6944 22986 6956
rect 22094 6916 22100 6928
rect 14608 6888 18368 6916
rect 18892 6888 22100 6916
rect 14608 6876 14614 6888
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 2746 6820 9689 6848
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 2746 6780 2774 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 17218 6848 17224 6860
rect 9999 6820 17224 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17420 6820 17724 6848
rect 9858 6780 9864 6792
rect 1627 6752 2774 6780
rect 9819 6752 9864 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 10060 6712 10088 6743
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10689 6783 10747 6789
rect 10192 6752 10237 6780
rect 10192 6740 10198 6752
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11330 6780 11336 6792
rect 10735 6752 11336 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11330 6740 11336 6752
rect 11388 6780 11394 6792
rect 11698 6780 11704 6792
rect 11388 6752 11704 6780
rect 11388 6740 11394 6752
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 16301 6783 16359 6789
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 16390 6780 16396 6792
rect 16347 6752 16396 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 17420 6789 17448 6820
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6749 17463 6783
rect 17586 6780 17592 6792
rect 17547 6752 17592 6780
rect 17405 6743 17463 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 17696 6780 17724 6820
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18230 6848 18236 6860
rect 18104 6820 18236 6848
rect 18104 6808 18110 6820
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18340 6848 18368 6888
rect 22094 6876 22100 6888
rect 22152 6876 22158 6928
rect 18598 6848 18604 6860
rect 18340 6820 18604 6848
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 21729 6851 21787 6857
rect 21729 6848 21741 6851
rect 18748 6820 21741 6848
rect 18748 6808 18754 6820
rect 21729 6817 21741 6820
rect 21775 6848 21787 6851
rect 22830 6848 22836 6860
rect 21775 6820 22836 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 23216 6848 23244 6956
rect 24210 6944 24216 6996
rect 24268 6984 24274 6996
rect 24581 6987 24639 6993
rect 24581 6984 24593 6987
rect 24268 6956 24593 6984
rect 24268 6944 24274 6956
rect 24581 6953 24593 6956
rect 24627 6984 24639 6987
rect 25222 6984 25228 6996
rect 24627 6956 25228 6984
rect 24627 6953 24639 6956
rect 24581 6947 24639 6953
rect 25222 6944 25228 6956
rect 25280 6944 25286 6996
rect 29546 6984 29552 6996
rect 27448 6956 29552 6984
rect 23750 6876 23756 6928
rect 23808 6916 23814 6928
rect 24946 6916 24952 6928
rect 23808 6888 24952 6916
rect 23808 6876 23814 6888
rect 24946 6876 24952 6888
rect 25004 6916 25010 6928
rect 25004 6888 25176 6916
rect 25004 6876 25010 6888
rect 23216 6820 25084 6848
rect 18138 6780 18144 6792
rect 17696 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 19794 6780 19800 6792
rect 18555 6752 19800 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 19794 6740 19800 6752
rect 19852 6780 19858 6792
rect 20070 6780 20076 6792
rect 19852 6752 20076 6780
rect 19852 6740 19858 6752
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 10502 6712 10508 6724
rect 10060 6684 10508 6712
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 18718 6715 18776 6721
rect 18718 6712 18730 6715
rect 13504 6684 18730 6712
rect 13504 6672 13510 6684
rect 18718 6681 18730 6684
rect 18764 6712 18776 6715
rect 18966 6712 18972 6724
rect 18764 6684 18972 6712
rect 18764 6681 18776 6684
rect 18718 6675 18776 6681
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 20180 6712 20208 6743
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 20312 6752 20453 6780
rect 20312 6740 20318 6752
rect 20441 6749 20453 6752
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 20809 6783 20867 6789
rect 20809 6780 20821 6783
rect 20680 6752 20821 6780
rect 20680 6740 20686 6752
rect 20809 6749 20821 6752
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 21082 6740 21088 6792
rect 21140 6780 21146 6792
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 21140 6752 21189 6780
rect 21140 6740 21146 6752
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6780 22063 6783
rect 22186 6780 22192 6792
rect 22051 6752 22192 6780
rect 22051 6749 22063 6752
rect 22005 6743 22063 6749
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 22298 6789 22304 6792
rect 22281 6783 22304 6789
rect 22281 6749 22293 6783
rect 22281 6743 22304 6749
rect 22298 6740 22304 6743
rect 22356 6740 22362 6792
rect 22462 6780 22468 6792
rect 22423 6752 22468 6780
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6780 22799 6783
rect 22787 6752 23060 6780
rect 22787 6749 22799 6752
rect 22741 6743 22799 6749
rect 21266 6712 21272 6724
rect 19668 6684 21272 6712
rect 19668 6672 19674 6684
rect 21266 6672 21272 6684
rect 21324 6672 21330 6724
rect 23032 6712 23060 6752
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23661 6783 23719 6789
rect 23661 6780 23673 6783
rect 23164 6752 23673 6780
rect 23164 6740 23170 6752
rect 23661 6749 23673 6752
rect 23707 6780 23719 6783
rect 23750 6780 23756 6792
rect 23707 6752 23756 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 23934 6780 23940 6792
rect 23895 6752 23940 6780
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 24118 6780 24124 6792
rect 24075 6752 24124 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24765 6783 24823 6789
rect 24765 6749 24777 6783
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 23382 6712 23388 6724
rect 23032 6684 23388 6712
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 23952 6712 23980 6740
rect 23676 6684 23980 6712
rect 24780 6712 24808 6743
rect 24854 6740 24860 6792
rect 24912 6780 24918 6792
rect 25056 6789 25084 6820
rect 25148 6789 25176 6888
rect 25590 6848 25596 6860
rect 25551 6820 25596 6848
rect 25590 6808 25596 6820
rect 25648 6808 25654 6860
rect 25041 6783 25099 6789
rect 24912 6752 24957 6780
rect 24912 6740 24918 6752
rect 25041 6749 25053 6783
rect 25087 6749 25099 6783
rect 25041 6743 25099 6749
rect 25133 6783 25191 6789
rect 25133 6749 25145 6783
rect 25179 6749 25191 6783
rect 25133 6743 25191 6749
rect 27062 6740 27068 6792
rect 27120 6780 27126 6792
rect 27448 6789 27476 6956
rect 29546 6944 29552 6956
rect 29604 6944 29610 6996
rect 30282 6944 30288 6996
rect 30340 6984 30346 6996
rect 33318 6984 33324 6996
rect 30340 6956 33324 6984
rect 30340 6944 30346 6956
rect 33134 6916 33140 6928
rect 32324 6888 33140 6916
rect 29454 6808 29460 6860
rect 29512 6848 29518 6860
rect 30190 6848 30196 6860
rect 29512 6820 30196 6848
rect 29512 6808 29518 6820
rect 30190 6808 30196 6820
rect 30248 6848 30254 6860
rect 30377 6851 30435 6857
rect 30377 6848 30389 6851
rect 30248 6820 30389 6848
rect 30248 6808 30254 6820
rect 30377 6817 30389 6820
rect 30423 6817 30435 6851
rect 30377 6811 30435 6817
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 32324 6848 32352 6888
rect 33134 6876 33140 6888
rect 33192 6876 33198 6928
rect 30524 6820 30569 6848
rect 30852 6820 32352 6848
rect 32401 6851 32459 6857
rect 30524 6808 30530 6820
rect 27433 6783 27491 6789
rect 27433 6780 27445 6783
rect 27120 6752 27445 6780
rect 27120 6740 27126 6752
rect 27433 6749 27445 6752
rect 27479 6749 27491 6783
rect 27433 6743 27491 6749
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 29270 6780 29276 6792
rect 27580 6752 29276 6780
rect 27580 6740 27586 6752
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 30852 6780 30880 6820
rect 32401 6817 32413 6851
rect 32447 6848 32459 6851
rect 32766 6848 32772 6860
rect 32447 6820 32772 6848
rect 32447 6817 32459 6820
rect 32401 6811 32459 6817
rect 32766 6808 32772 6820
rect 32824 6808 32830 6860
rect 33244 6848 33272 6956
rect 33318 6944 33324 6956
rect 33376 6944 33382 6996
rect 34146 6944 34152 6996
rect 34204 6984 34210 6996
rect 35250 6984 35256 6996
rect 34204 6956 35256 6984
rect 34204 6944 34210 6956
rect 35250 6944 35256 6956
rect 35308 6984 35314 6996
rect 35710 6984 35716 6996
rect 35308 6956 35716 6984
rect 35308 6944 35314 6956
rect 35710 6944 35716 6956
rect 35768 6944 35774 6996
rect 35986 6984 35992 6996
rect 35866 6956 35992 6984
rect 33594 6876 33600 6928
rect 33652 6916 33658 6928
rect 34882 6916 34888 6928
rect 33652 6888 34888 6916
rect 33652 6876 33658 6888
rect 34882 6876 34888 6888
rect 34940 6876 34946 6928
rect 35866 6916 35894 6956
rect 35986 6944 35992 6956
rect 36044 6944 36050 6996
rect 36078 6944 36084 6996
rect 36136 6984 36142 6996
rect 38289 6987 38347 6993
rect 36136 6956 38240 6984
rect 36136 6944 36142 6956
rect 35268 6888 35894 6916
rect 36449 6919 36507 6925
rect 33686 6848 33692 6860
rect 32876 6820 33272 6848
rect 33428 6820 33692 6848
rect 31110 6780 31116 6792
rect 29932 6752 30880 6780
rect 31071 6752 31116 6780
rect 25682 6712 25688 6724
rect 24780 6684 25688 6712
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 17494 6644 17500 6656
rect 14884 6616 17500 6644
rect 14884 6604 14890 6616
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 23014 6644 23020 6656
rect 20404 6616 23020 6644
rect 20404 6604 20410 6616
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23109 6647 23167 6653
rect 23109 6613 23121 6647
rect 23155 6644 23167 6647
rect 23676 6644 23704 6684
rect 25682 6672 25688 6684
rect 25740 6672 25746 6724
rect 25860 6715 25918 6721
rect 25860 6681 25872 6715
rect 25906 6712 25918 6715
rect 26050 6712 26056 6724
rect 25906 6684 26056 6712
rect 25906 6681 25918 6684
rect 25860 6675 25918 6681
rect 26050 6672 26056 6684
rect 26108 6672 26114 6724
rect 27700 6715 27758 6721
rect 27700 6681 27712 6715
rect 27746 6712 27758 6715
rect 27982 6712 27988 6724
rect 27746 6684 27988 6712
rect 27746 6681 27758 6684
rect 27700 6675 27758 6681
rect 27982 6672 27988 6684
rect 28040 6672 28046 6724
rect 28718 6712 28724 6724
rect 28092 6684 28724 6712
rect 23155 6616 23704 6644
rect 23155 6613 23167 6616
rect 23109 6607 23167 6613
rect 23750 6604 23756 6656
rect 23808 6644 23814 6656
rect 26970 6644 26976 6656
rect 23808 6616 26976 6644
rect 23808 6604 23814 6616
rect 26970 6604 26976 6616
rect 27028 6604 27034 6656
rect 27338 6604 27344 6656
rect 27396 6644 27402 6656
rect 27522 6644 27528 6656
rect 27396 6616 27528 6644
rect 27396 6604 27402 6616
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 27890 6604 27896 6656
rect 27948 6644 27954 6656
rect 28092 6644 28120 6684
rect 28718 6672 28724 6684
rect 28776 6672 28782 6724
rect 28810 6644 28816 6656
rect 27948 6616 28120 6644
rect 28771 6616 28816 6644
rect 27948 6604 27954 6616
rect 28810 6604 28816 6616
rect 28868 6604 28874 6656
rect 29932 6653 29960 6752
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 31202 6740 31208 6792
rect 31260 6780 31266 6792
rect 31481 6783 31539 6789
rect 31481 6780 31493 6783
rect 31260 6752 31493 6780
rect 31260 6740 31266 6752
rect 31481 6749 31493 6752
rect 31527 6749 31539 6783
rect 31481 6743 31539 6749
rect 32585 6783 32643 6789
rect 32585 6749 32597 6783
rect 32631 6749 32643 6783
rect 32585 6743 32643 6749
rect 31018 6672 31024 6724
rect 31076 6712 31082 6724
rect 31297 6715 31355 6721
rect 31297 6712 31309 6715
rect 31076 6684 31309 6712
rect 31076 6672 31082 6684
rect 31297 6681 31309 6684
rect 31343 6681 31355 6715
rect 31297 6675 31355 6681
rect 31389 6715 31447 6721
rect 31389 6681 31401 6715
rect 31435 6712 31447 6715
rect 31570 6712 31576 6724
rect 31435 6684 31576 6712
rect 31435 6681 31447 6684
rect 31389 6675 31447 6681
rect 31570 6672 31576 6684
rect 31628 6672 31634 6724
rect 32600 6712 32628 6743
rect 32674 6740 32680 6792
rect 32732 6780 32738 6792
rect 32876 6789 32904 6820
rect 32861 6783 32919 6789
rect 32732 6752 32777 6780
rect 32732 6740 32738 6752
rect 32861 6749 32873 6783
rect 32907 6749 32919 6783
rect 32861 6743 32919 6749
rect 32953 6783 33011 6789
rect 32953 6749 32965 6783
rect 32999 6780 33011 6783
rect 33134 6780 33140 6792
rect 32999 6752 33140 6780
rect 32999 6749 33011 6752
rect 32953 6743 33011 6749
rect 33134 6740 33140 6752
rect 33192 6740 33198 6792
rect 33428 6789 33456 6820
rect 33686 6808 33692 6820
rect 33744 6848 33750 6860
rect 34238 6848 34244 6860
rect 33744 6820 34244 6848
rect 33744 6808 33750 6820
rect 34238 6808 34244 6820
rect 34296 6808 34302 6860
rect 34790 6848 34796 6860
rect 34348 6820 34796 6848
rect 33413 6783 33471 6789
rect 33413 6749 33425 6783
rect 33459 6749 33471 6783
rect 33413 6743 33471 6749
rect 33561 6783 33619 6789
rect 33561 6749 33573 6783
rect 33607 6780 33619 6783
rect 33778 6780 33784 6792
rect 33607 6749 33640 6780
rect 33739 6752 33784 6780
rect 33561 6743 33640 6749
rect 33042 6712 33048 6724
rect 32600 6684 33048 6712
rect 33042 6672 33048 6684
rect 33100 6672 33106 6724
rect 33612 6712 33640 6743
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 33962 6789 33968 6792
rect 33919 6783 33968 6789
rect 33919 6749 33931 6783
rect 33965 6749 33968 6783
rect 33919 6743 33968 6749
rect 33962 6740 33968 6743
rect 34020 6740 34026 6792
rect 33428 6684 33640 6712
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6613 29975 6647
rect 29917 6607 29975 6613
rect 30285 6647 30343 6653
rect 30285 6613 30297 6647
rect 30331 6644 30343 6647
rect 30374 6644 30380 6656
rect 30331 6616 30380 6644
rect 30331 6613 30343 6616
rect 30285 6607 30343 6613
rect 30374 6604 30380 6616
rect 30432 6644 30438 6656
rect 31478 6644 31484 6656
rect 30432 6616 31484 6644
rect 30432 6604 30438 6616
rect 31478 6604 31484 6616
rect 31536 6604 31542 6656
rect 31662 6644 31668 6656
rect 31623 6616 31668 6644
rect 31662 6604 31668 6616
rect 31720 6604 31726 6656
rect 32214 6604 32220 6656
rect 32272 6644 32278 6656
rect 33226 6644 33232 6656
rect 32272 6616 33232 6644
rect 32272 6604 32278 6616
rect 33226 6604 33232 6616
rect 33284 6644 33290 6656
rect 33428 6644 33456 6684
rect 33686 6672 33692 6724
rect 33744 6712 33750 6724
rect 34348 6712 34376 6820
rect 34790 6808 34796 6820
rect 34848 6808 34854 6860
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 33744 6684 34376 6712
rect 34440 6752 34897 6780
rect 33744 6672 33750 6684
rect 33284 6616 33456 6644
rect 34057 6647 34115 6653
rect 33284 6604 33290 6616
rect 34057 6613 34069 6647
rect 34103 6644 34115 6647
rect 34440 6644 34468 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 34606 6672 34612 6724
rect 34664 6712 34670 6724
rect 35268 6712 35296 6888
rect 36449 6885 36461 6919
rect 36495 6916 36507 6919
rect 36906 6916 36912 6928
rect 36495 6888 36912 6916
rect 36495 6885 36507 6888
rect 36449 6879 36507 6885
rect 36906 6876 36912 6888
rect 36964 6916 36970 6928
rect 37826 6916 37832 6928
rect 36964 6888 37832 6916
rect 36964 6876 36970 6888
rect 37826 6876 37832 6888
rect 37884 6876 37890 6928
rect 38212 6916 38240 6956
rect 38289 6953 38301 6987
rect 38335 6984 38347 6987
rect 38378 6984 38384 6996
rect 38335 6956 38384 6984
rect 38335 6953 38347 6956
rect 38289 6947 38347 6953
rect 38378 6944 38384 6956
rect 38436 6944 38442 6996
rect 42794 6984 42800 6996
rect 42755 6956 42800 6984
rect 42794 6944 42800 6956
rect 42852 6944 42858 6996
rect 58250 6984 58256 6996
rect 58211 6956 58256 6984
rect 58250 6944 58256 6956
rect 58308 6944 58314 6996
rect 38212 6888 38654 6916
rect 35462 6851 35520 6857
rect 35462 6817 35474 6851
rect 35508 6848 35520 6851
rect 35618 6848 35624 6860
rect 35508 6820 35624 6848
rect 35508 6817 35520 6820
rect 35462 6811 35520 6817
rect 35618 6808 35624 6820
rect 35676 6808 35682 6860
rect 35912 6820 37412 6848
rect 35342 6740 35348 6792
rect 35400 6789 35406 6792
rect 35400 6783 35421 6789
rect 35409 6749 35421 6783
rect 35400 6743 35421 6749
rect 35400 6740 35406 6743
rect 35710 6740 35716 6792
rect 35768 6780 35774 6792
rect 35912 6780 35940 6820
rect 35768 6752 35940 6780
rect 35768 6740 35774 6752
rect 36078 6740 36084 6792
rect 36136 6780 36142 6792
rect 36173 6783 36231 6789
rect 36173 6780 36185 6783
rect 36136 6752 36185 6780
rect 36136 6740 36142 6752
rect 36173 6749 36185 6752
rect 36219 6749 36231 6783
rect 36173 6743 36231 6749
rect 36354 6740 36360 6792
rect 36412 6780 36418 6792
rect 36998 6780 37004 6792
rect 36412 6752 37004 6780
rect 36412 6740 36418 6752
rect 36998 6740 37004 6752
rect 37056 6740 37062 6792
rect 37384 6789 37412 6820
rect 37642 6808 37648 6860
rect 37700 6848 37706 6860
rect 37921 6851 37979 6857
rect 37921 6848 37933 6851
rect 37700 6820 37933 6848
rect 37700 6808 37706 6820
rect 37921 6817 37933 6820
rect 37967 6848 37979 6851
rect 38286 6848 38292 6860
rect 37967 6820 38292 6848
rect 37967 6817 37979 6820
rect 37921 6811 37979 6817
rect 38286 6808 38292 6820
rect 38344 6808 38350 6860
rect 38626 6848 38654 6888
rect 41598 6876 41604 6928
rect 41656 6916 41662 6928
rect 47670 6916 47676 6928
rect 41656 6888 47676 6916
rect 41656 6876 41662 6888
rect 40129 6851 40187 6857
rect 40129 6848 40141 6851
rect 38626 6820 40141 6848
rect 40129 6817 40141 6820
rect 40175 6817 40187 6851
rect 42058 6848 42064 6860
rect 40129 6811 40187 6817
rect 41156 6820 41920 6848
rect 42019 6820 42064 6848
rect 37185 6783 37243 6789
rect 37185 6749 37197 6783
rect 37231 6749 37243 6783
rect 37185 6743 37243 6749
rect 37369 6783 37427 6789
rect 37369 6749 37381 6783
rect 37415 6749 37427 6783
rect 38105 6783 38163 6789
rect 37369 6743 37427 6749
rect 37461 6761 37519 6767
rect 34664 6684 35296 6712
rect 34664 6672 34670 6684
rect 35986 6672 35992 6724
rect 36044 6712 36050 6724
rect 37200 6712 37228 6743
rect 37461 6727 37473 6761
rect 37507 6727 37519 6761
rect 38105 6749 38117 6783
rect 38151 6749 38163 6783
rect 38105 6743 38163 6749
rect 37461 6721 37519 6727
rect 36044 6684 37228 6712
rect 36044 6672 36050 6684
rect 34103 6616 34468 6644
rect 35069 6647 35127 6653
rect 34103 6613 34115 6616
rect 34057 6607 34115 6613
rect 35069 6613 35081 6647
rect 35115 6644 35127 6647
rect 36078 6644 36084 6656
rect 35115 6616 36084 6644
rect 35115 6613 35127 6616
rect 35069 6607 35127 6613
rect 36078 6604 36084 6616
rect 36136 6604 36142 6656
rect 36262 6604 36268 6656
rect 36320 6644 36326 6656
rect 36538 6644 36544 6656
rect 36320 6616 36544 6644
rect 36320 6604 36326 6616
rect 36538 6604 36544 6616
rect 36596 6604 36602 6656
rect 36998 6644 37004 6656
rect 36959 6616 37004 6644
rect 36998 6604 37004 6616
rect 37056 6604 37062 6656
rect 37476 6644 37504 6721
rect 37826 6672 37832 6724
rect 37884 6712 37890 6724
rect 38121 6712 38149 6743
rect 38470 6740 38476 6792
rect 38528 6780 38534 6792
rect 40034 6780 40040 6792
rect 38528 6752 40040 6780
rect 38528 6740 38534 6752
rect 40034 6740 40040 6752
rect 40092 6740 40098 6792
rect 37884 6684 38149 6712
rect 37884 6672 37890 6684
rect 38194 6672 38200 6724
rect 38252 6712 38258 6724
rect 40144 6712 40172 6811
rect 40586 6740 40592 6792
rect 40644 6780 40650 6792
rect 40862 6780 40868 6792
rect 40644 6752 40868 6780
rect 40644 6740 40650 6752
rect 40862 6740 40868 6752
rect 40920 6780 40926 6792
rect 41156 6789 41184 6820
rect 40957 6783 41015 6789
rect 40957 6780 40969 6783
rect 40920 6752 40969 6780
rect 40920 6740 40926 6752
rect 40957 6749 40969 6752
rect 41003 6749 41015 6783
rect 40957 6743 41015 6749
rect 41141 6783 41199 6789
rect 41141 6749 41153 6783
rect 41187 6749 41199 6783
rect 41785 6783 41843 6789
rect 41785 6780 41797 6783
rect 41141 6743 41199 6749
rect 41248 6752 41797 6780
rect 41248 6712 41276 6752
rect 41785 6749 41797 6752
rect 41831 6749 41843 6783
rect 41785 6743 41843 6749
rect 38252 6684 39252 6712
rect 40144 6684 41276 6712
rect 41325 6715 41383 6721
rect 38252 6672 38258 6684
rect 37918 6644 37924 6656
rect 37476 6616 37924 6644
rect 37918 6604 37924 6616
rect 37976 6604 37982 6656
rect 39224 6644 39252 6684
rect 41325 6681 41337 6715
rect 41371 6712 41383 6715
rect 41690 6712 41696 6724
rect 41371 6684 41696 6712
rect 41371 6681 41383 6684
rect 41325 6675 41383 6681
rect 41690 6672 41696 6684
rect 41748 6672 41754 6724
rect 41892 6712 41920 6820
rect 42058 6808 42064 6820
rect 42116 6808 42122 6860
rect 43057 6848 43085 6888
rect 47670 6876 47676 6888
rect 47728 6876 47734 6928
rect 43993 6851 44051 6857
rect 43993 6848 44005 6851
rect 42996 6820 43085 6848
rect 43456 6820 44005 6848
rect 42996 6789 43024 6820
rect 43456 6792 43484 6820
rect 43993 6817 44005 6820
rect 44039 6817 44051 6851
rect 56870 6848 56876 6860
rect 56831 6820 56876 6848
rect 43993 6811 44051 6817
rect 56870 6808 56876 6820
rect 56928 6808 56934 6860
rect 42973 6783 43031 6789
rect 42973 6749 42985 6783
rect 43019 6749 43031 6783
rect 43105 6783 43163 6789
rect 43105 6780 43117 6783
rect 42973 6743 43031 6749
rect 43088 6749 43117 6780
rect 43151 6749 43163 6783
rect 43254 6780 43260 6792
rect 43215 6752 43260 6780
rect 43088 6743 43163 6749
rect 43088 6712 43116 6743
rect 43254 6740 43260 6752
rect 43312 6740 43318 6792
rect 43349 6783 43407 6789
rect 43349 6749 43361 6783
rect 43395 6780 43407 6783
rect 43438 6780 43444 6792
rect 43395 6752 43444 6780
rect 43395 6749 43407 6752
rect 43349 6743 43407 6749
rect 43438 6740 43444 6752
rect 43496 6740 43502 6792
rect 43806 6780 43812 6792
rect 43767 6752 43812 6780
rect 43806 6740 43812 6752
rect 43864 6740 43870 6792
rect 56778 6740 56784 6792
rect 56836 6780 56842 6792
rect 57129 6783 57187 6789
rect 57129 6780 57141 6783
rect 56836 6752 57141 6780
rect 56836 6740 56842 6752
rect 57129 6749 57141 6752
rect 57175 6749 57187 6783
rect 57129 6743 57187 6749
rect 45278 6712 45284 6724
rect 41892 6684 45284 6712
rect 45278 6672 45284 6684
rect 45336 6672 45342 6724
rect 56042 6712 56048 6724
rect 51046 6684 56048 6712
rect 51046 6644 51074 6684
rect 56042 6672 56048 6684
rect 56100 6672 56106 6724
rect 39224 6616 51074 6644
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10594 6440 10600 6452
rect 10183 6412 10600 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 15344 6412 17325 6440
rect 15344 6400 15350 6412
rect 17313 6409 17325 6412
rect 17359 6409 17371 6443
rect 17313 6403 17371 6409
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 19334 6440 19340 6452
rect 18104 6412 19340 6440
rect 18104 6400 18110 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 21082 6440 21088 6452
rect 20036 6412 21088 6440
rect 20036 6400 20042 6412
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 21177 6443 21235 6449
rect 21177 6409 21189 6443
rect 21223 6440 21235 6443
rect 22646 6440 22652 6452
rect 21223 6412 22652 6440
rect 21223 6409 21235 6412
rect 21177 6403 21235 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 22830 6400 22836 6452
rect 22888 6440 22894 6452
rect 23290 6440 23296 6452
rect 22888 6412 23296 6440
rect 22888 6400 22894 6412
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 26786 6400 26792 6452
rect 26844 6440 26850 6452
rect 27525 6443 27583 6449
rect 27525 6440 27537 6443
rect 26844 6412 27537 6440
rect 26844 6400 26850 6412
rect 27525 6409 27537 6412
rect 27571 6409 27583 6443
rect 27982 6440 27988 6452
rect 27943 6412 27988 6440
rect 27525 6403 27583 6409
rect 27982 6400 27988 6412
rect 28040 6400 28046 6452
rect 28353 6443 28411 6449
rect 28353 6409 28365 6443
rect 28399 6440 28411 6443
rect 29454 6440 29460 6452
rect 28399 6412 29460 6440
rect 28399 6409 28411 6412
rect 28353 6403 28411 6409
rect 29454 6400 29460 6412
rect 29512 6400 29518 6452
rect 36170 6440 36176 6452
rect 29564 6412 36176 6440
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 20530 6372 20536 6384
rect 9732 6344 9777 6372
rect 12406 6344 20536 6372
rect 9732 6332 9738 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 9582 6304 9588 6316
rect 1627 6276 9588 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11606 6304 11612 6316
rect 10919 6276 11612 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11756 6276 11801 6304
rect 11756 6264 11762 6276
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 12406 6236 12434 6344
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 21726 6332 21732 6384
rect 21784 6332 21790 6384
rect 22094 6332 22100 6384
rect 22152 6372 22158 6384
rect 28445 6375 28503 6381
rect 28445 6372 28457 6375
rect 22152 6344 28457 6372
rect 22152 6332 22158 6344
rect 28445 6341 28457 6344
rect 28491 6372 28503 6375
rect 28810 6372 28816 6384
rect 28491 6344 28816 6372
rect 28491 6341 28503 6344
rect 28445 6335 28503 6341
rect 28810 6332 28816 6344
rect 28868 6332 28874 6384
rect 29178 6332 29184 6384
rect 29236 6372 29242 6384
rect 29273 6375 29331 6381
rect 29273 6372 29285 6375
rect 29236 6344 29285 6372
rect 29236 6332 29242 6344
rect 29273 6341 29285 6344
rect 29319 6341 29331 6375
rect 29273 6335 29331 6341
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 15896 6276 16865 6304
rect 15896 6264 15902 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18748 6276 18889 6304
rect 18748 6264 18754 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19978 6304 19984 6316
rect 19300 6276 19984 6304
rect 19300 6264 19306 6276
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20254 6304 20260 6316
rect 20128 6276 20260 6304
rect 20128 6264 20134 6276
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20714 6304 20720 6316
rect 20675 6276 20720 6304
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21324 6276 21373 6304
rect 21324 6264 21330 6276
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21744 6304 21772 6332
rect 22002 6304 22008 6316
rect 21744 6276 22008 6304
rect 21361 6267 21419 6273
rect 22002 6264 22008 6276
rect 22060 6264 22066 6316
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 8996 6208 12434 6236
rect 8996 6196 9002 6208
rect 18966 6196 18972 6248
rect 19024 6236 19030 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 19024 6208 19165 6236
rect 19024 6196 19030 6208
rect 19153 6205 19165 6208
rect 19199 6236 19211 6239
rect 19886 6236 19892 6248
rect 19199 6208 19892 6236
rect 19199 6205 19211 6208
rect 19153 6199 19211 6205
rect 19886 6196 19892 6208
rect 19944 6236 19950 6248
rect 20732 6236 20760 6264
rect 19944 6208 20760 6236
rect 19944 6196 19950 6208
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 21910 6236 21916 6248
rect 21784 6208 21916 6236
rect 21784 6196 21790 6208
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22296 6236 22324 6267
rect 22462 6264 22468 6316
rect 22520 6304 22526 6316
rect 22741 6307 22799 6313
rect 22741 6304 22753 6307
rect 22520 6276 22753 6304
rect 22520 6264 22526 6276
rect 22741 6273 22753 6276
rect 22787 6273 22799 6307
rect 23198 6304 23204 6316
rect 23159 6276 23204 6304
rect 22741 6267 22799 6273
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 24946 6304 24952 6316
rect 23348 6276 24952 6304
rect 23348 6264 23354 6276
rect 24946 6264 24952 6276
rect 25004 6264 25010 6316
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6304 25559 6307
rect 27341 6307 27399 6313
rect 25547 6276 27292 6304
rect 25547 6273 25559 6276
rect 25501 6267 25559 6273
rect 24210 6236 24216 6248
rect 22296 6208 24216 6236
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 25777 6239 25835 6245
rect 25777 6205 25789 6239
rect 25823 6205 25835 6239
rect 27154 6236 27160 6248
rect 27115 6208 27160 6236
rect 25777 6199 25835 6205
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 5132 6140 9965 6168
rect 5132 6128 5138 6140
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 11054 6168 11060 6180
rect 11015 6140 11060 6168
rect 9953 6131 10011 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 17126 6168 17132 6180
rect 17087 6140 17132 6168
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 22097 6171 22155 6177
rect 17828 6140 22048 6168
rect 17828 6128 17834 6140
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 10376 6072 11897 6100
rect 10376 6060 10382 6072
rect 11885 6069 11897 6072
rect 11931 6069 11943 6103
rect 16298 6100 16304 6112
rect 16259 6072 16304 6100
rect 11885 6063 11943 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6100 18475 6103
rect 21910 6100 21916 6112
rect 18463 6072 21916 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 21910 6060 21916 6072
rect 21968 6060 21974 6112
rect 22020 6100 22048 6140
rect 22097 6137 22109 6171
rect 22143 6168 22155 6171
rect 22186 6168 22192 6180
rect 22143 6140 22192 6168
rect 22143 6137 22155 6140
rect 22097 6131 22155 6137
rect 22186 6128 22192 6140
rect 22244 6168 22250 6180
rect 25038 6168 25044 6180
rect 22244 6140 25044 6168
rect 22244 6128 22250 6140
rect 25038 6128 25044 6140
rect 25096 6128 25102 6180
rect 25498 6128 25504 6180
rect 25556 6168 25562 6180
rect 25792 6168 25820 6199
rect 27154 6196 27160 6208
rect 27212 6196 27218 6248
rect 27264 6236 27292 6276
rect 27341 6273 27353 6307
rect 27387 6304 27399 6307
rect 27522 6304 27528 6316
rect 27387 6276 27528 6304
rect 27387 6273 27399 6276
rect 27341 6267 27399 6273
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 29362 6304 29368 6316
rect 28460 6276 29368 6304
rect 28460 6236 28488 6276
rect 29362 6264 29368 6276
rect 29420 6264 29426 6316
rect 29564 6313 29592 6412
rect 36170 6400 36176 6412
rect 36228 6400 36234 6452
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 36596 6412 37688 6440
rect 36596 6400 36602 6412
rect 31662 6372 31668 6384
rect 29840 6344 31668 6372
rect 29457 6307 29515 6313
rect 29457 6273 29469 6307
rect 29503 6273 29515 6307
rect 29457 6267 29515 6273
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6273 29607 6307
rect 29730 6304 29736 6316
rect 29691 6276 29736 6304
rect 29549 6267 29607 6273
rect 28626 6236 28632 6248
rect 27264 6208 28488 6236
rect 28587 6208 28632 6236
rect 28626 6196 28632 6208
rect 28684 6196 28690 6248
rect 29472 6236 29500 6267
rect 29730 6264 29736 6276
rect 29788 6264 29794 6316
rect 29840 6313 29868 6344
rect 31662 6332 31668 6344
rect 31720 6332 31726 6384
rect 32490 6332 32496 6384
rect 32548 6372 32554 6384
rect 34238 6372 34244 6384
rect 32548 6344 33548 6372
rect 34151 6344 34244 6372
rect 32548 6332 32554 6344
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6273 29883 6307
rect 30282 6304 30288 6316
rect 30243 6276 30288 6304
rect 29825 6267 29883 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 31389 6307 31447 6313
rect 31389 6304 31401 6307
rect 30392 6276 31401 6304
rect 29914 6236 29920 6248
rect 29472 6208 29920 6236
rect 29914 6196 29920 6208
rect 29972 6196 29978 6248
rect 25556 6140 25820 6168
rect 25556 6128 25562 6140
rect 26602 6128 26608 6180
rect 26660 6168 26666 6180
rect 30392 6168 30420 6276
rect 31389 6273 31401 6276
rect 31435 6273 31447 6307
rect 32306 6304 32312 6316
rect 32267 6276 32312 6304
rect 31389 6267 31447 6273
rect 32306 6264 32312 6276
rect 32364 6264 32370 6316
rect 32576 6307 32634 6313
rect 32576 6273 32588 6307
rect 32622 6304 32634 6307
rect 33520 6304 33548 6344
rect 34238 6332 34244 6344
rect 34296 6372 34302 6384
rect 34790 6372 34796 6384
rect 34296 6344 34796 6372
rect 34296 6332 34302 6344
rect 34790 6332 34796 6344
rect 34848 6332 34854 6384
rect 35250 6372 35256 6384
rect 35211 6344 35256 6372
rect 35250 6332 35256 6344
rect 35308 6332 35314 6384
rect 35345 6375 35403 6381
rect 35345 6341 35357 6375
rect 35391 6372 35403 6375
rect 36262 6372 36268 6384
rect 35391 6344 36268 6372
rect 35391 6341 35403 6344
rect 35345 6335 35403 6341
rect 36262 6332 36268 6344
rect 36320 6332 36326 6384
rect 34425 6307 34483 6313
rect 34425 6304 34437 6307
rect 32622 6276 33456 6304
rect 33520 6276 34437 6304
rect 32622 6273 32634 6276
rect 32576 6267 32634 6273
rect 30561 6239 30619 6245
rect 30561 6205 30573 6239
rect 30607 6236 30619 6239
rect 33428 6236 33456 6276
rect 34425 6273 34437 6276
rect 34471 6273 34483 6307
rect 34425 6267 34483 6273
rect 34514 6264 34520 6316
rect 34572 6304 34578 6316
rect 35158 6313 35164 6316
rect 34977 6307 35035 6313
rect 34572 6276 34617 6304
rect 34572 6264 34578 6276
rect 34977 6273 34989 6307
rect 35023 6273 35035 6307
rect 34977 6267 35035 6273
rect 35115 6307 35164 6313
rect 35115 6273 35127 6307
rect 35161 6273 35164 6307
rect 35115 6267 35164 6273
rect 34146 6236 34152 6248
rect 30607 6208 31984 6236
rect 33428 6208 34152 6236
rect 30607 6205 30619 6208
rect 30561 6199 30619 6205
rect 26660 6140 30420 6168
rect 26660 6128 26666 6140
rect 22278 6100 22284 6112
rect 22020 6072 22284 6100
rect 22278 6060 22284 6072
rect 22336 6060 22342 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 28994 6100 29000 6112
rect 23808 6072 29000 6100
rect 23808 6060 23814 6072
rect 28994 6060 29000 6072
rect 29052 6060 29058 6112
rect 29178 6060 29184 6112
rect 29236 6100 29242 6112
rect 30576 6100 30604 6199
rect 30837 6171 30895 6177
rect 30837 6137 30849 6171
rect 30883 6168 30895 6171
rect 30883 6140 31616 6168
rect 30883 6137 30895 6140
rect 30837 6131 30895 6137
rect 29236 6072 30604 6100
rect 30653 6103 30711 6109
rect 29236 6060 29242 6072
rect 30653 6069 30665 6103
rect 30699 6100 30711 6103
rect 31110 6100 31116 6112
rect 30699 6072 31116 6100
rect 30699 6069 30711 6072
rect 30653 6063 30711 6069
rect 31110 6060 31116 6072
rect 31168 6060 31174 6112
rect 31478 6100 31484 6112
rect 31439 6072 31484 6100
rect 31478 6060 31484 6072
rect 31536 6060 31542 6112
rect 31588 6100 31616 6140
rect 31846 6100 31852 6112
rect 31588 6072 31852 6100
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 31956 6100 31984 6208
rect 34146 6196 34152 6208
rect 34204 6196 34210 6248
rect 34532 6236 34560 6264
rect 34348 6208 34560 6236
rect 33594 6128 33600 6180
rect 33652 6168 33658 6180
rect 33689 6171 33747 6177
rect 33689 6168 33701 6171
rect 33652 6140 33701 6168
rect 33652 6128 33658 6140
rect 33689 6137 33701 6140
rect 33735 6137 33747 6171
rect 33689 6131 33747 6137
rect 34054 6128 34060 6180
rect 34112 6168 34118 6180
rect 34241 6171 34299 6177
rect 34241 6168 34253 6171
rect 34112 6140 34253 6168
rect 34112 6128 34118 6140
rect 34241 6137 34253 6140
rect 34287 6137 34299 6171
rect 34241 6131 34299 6137
rect 34348 6100 34376 6208
rect 34606 6196 34612 6248
rect 34664 6236 34670 6248
rect 34992 6236 35020 6267
rect 35158 6264 35164 6267
rect 35216 6264 35222 6316
rect 35526 6313 35532 6316
rect 35483 6307 35532 6313
rect 35483 6273 35495 6307
rect 35529 6273 35532 6307
rect 35483 6267 35532 6273
rect 35526 6264 35532 6267
rect 35584 6264 35590 6316
rect 35802 6264 35808 6316
rect 35860 6304 35866 6316
rect 36354 6304 36360 6316
rect 35860 6276 36360 6304
rect 35860 6264 35866 6276
rect 36354 6264 36360 6276
rect 36412 6264 36418 6316
rect 36541 6307 36599 6313
rect 36541 6273 36553 6307
rect 36587 6304 36599 6307
rect 36998 6304 37004 6316
rect 36587 6276 37004 6304
rect 36587 6273 36599 6276
rect 36541 6267 36599 6273
rect 36998 6264 37004 6276
rect 37056 6264 37062 6316
rect 37090 6264 37096 6316
rect 37148 6304 37154 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37148 6276 37473 6304
rect 37148 6264 37154 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37660 6304 37688 6412
rect 38194 6400 38200 6452
rect 38252 6440 38258 6452
rect 38252 6412 38424 6440
rect 38252 6400 38258 6412
rect 37728 6375 37786 6381
rect 37728 6341 37740 6375
rect 37774 6372 37786 6375
rect 38286 6372 38292 6384
rect 37774 6344 38292 6372
rect 37774 6341 37786 6344
rect 37728 6335 37786 6341
rect 38286 6332 38292 6344
rect 38344 6332 38350 6384
rect 38396 6372 38424 6412
rect 39022 6400 39028 6452
rect 39080 6440 39086 6452
rect 39485 6443 39543 6449
rect 39485 6440 39497 6443
rect 39080 6412 39497 6440
rect 39080 6400 39086 6412
rect 39485 6409 39497 6412
rect 39531 6409 39543 6443
rect 39485 6403 39543 6409
rect 40034 6400 40040 6452
rect 40092 6440 40098 6452
rect 43254 6440 43260 6452
rect 40092 6412 43260 6440
rect 40092 6400 40098 6412
rect 43254 6400 43260 6412
rect 43312 6400 43318 6452
rect 56134 6440 56140 6452
rect 55784 6412 56140 6440
rect 43272 6372 43300 6400
rect 44085 6375 44143 6381
rect 38396 6344 39344 6372
rect 43272 6344 43668 6372
rect 39316 6313 39344 6344
rect 39301 6307 39359 6313
rect 37660 6276 38654 6304
rect 37461 6267 37519 6273
rect 34664 6208 35020 6236
rect 34664 6196 34670 6208
rect 35618 6196 35624 6248
rect 35676 6196 35682 6248
rect 36081 6239 36139 6245
rect 36081 6236 36093 6239
rect 35912 6208 36093 6236
rect 34422 6128 34428 6180
rect 34480 6168 34486 6180
rect 35636 6168 35664 6196
rect 35912 6168 35940 6208
rect 36081 6205 36093 6208
rect 36127 6236 36139 6239
rect 37182 6236 37188 6248
rect 36127 6208 37188 6236
rect 36127 6205 36139 6208
rect 36081 6199 36139 6205
rect 37182 6196 37188 6208
rect 37240 6196 37246 6248
rect 38626 6236 38654 6276
rect 39301 6273 39313 6307
rect 39347 6273 39359 6307
rect 39301 6267 39359 6273
rect 41782 6264 41788 6316
rect 41840 6304 41846 6316
rect 43640 6313 43668 6344
rect 44085 6341 44097 6375
rect 44131 6372 44143 6375
rect 45094 6372 45100 6384
rect 44131 6344 45100 6372
rect 44131 6341 44143 6344
rect 44085 6335 44143 6341
rect 45094 6332 45100 6344
rect 45152 6332 45158 6384
rect 55784 6381 55812 6412
rect 56134 6400 56140 6412
rect 56192 6400 56198 6452
rect 55769 6375 55827 6381
rect 55769 6341 55781 6375
rect 55815 6341 55827 6375
rect 55769 6335 55827 6341
rect 55953 6375 56011 6381
rect 55953 6341 55965 6375
rect 55999 6372 56011 6375
rect 57238 6372 57244 6384
rect 55999 6344 57244 6372
rect 55999 6341 56011 6344
rect 55953 6335 56011 6341
rect 57238 6332 57244 6344
rect 57296 6332 57302 6384
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 41840 6276 42901 6304
rect 41840 6264 41846 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 42889 6267 42947 6273
rect 43533 6307 43591 6313
rect 43533 6273 43545 6307
rect 43579 6273 43591 6307
rect 43533 6267 43591 6273
rect 43625 6307 43683 6313
rect 43625 6273 43637 6307
rect 43671 6273 43683 6307
rect 43625 6267 43683 6273
rect 43548 6236 43576 6267
rect 56042 6264 56048 6316
rect 56100 6304 56106 6316
rect 56597 6307 56655 6313
rect 56100 6276 56145 6304
rect 56100 6264 56106 6276
rect 56597 6273 56609 6307
rect 56643 6304 56655 6307
rect 56686 6304 56692 6316
rect 56643 6276 56692 6304
rect 56643 6273 56655 6276
rect 56597 6267 56655 6273
rect 56686 6264 56692 6276
rect 56744 6264 56750 6316
rect 58066 6304 58072 6316
rect 58027 6276 58072 6304
rect 58066 6264 58072 6276
rect 58124 6264 58130 6316
rect 45002 6236 45008 6248
rect 38626 6208 43484 6236
rect 43548 6208 45008 6236
rect 34480 6140 35940 6168
rect 34480 6128 34486 6140
rect 35986 6128 35992 6180
rect 36044 6168 36050 6180
rect 36357 6171 36415 6177
rect 36357 6168 36369 6171
rect 36044 6140 36369 6168
rect 36044 6128 36050 6140
rect 36357 6137 36369 6140
rect 36403 6137 36415 6171
rect 41690 6168 41696 6180
rect 36357 6131 36415 6137
rect 38396 6140 41696 6168
rect 31956 6072 34376 6100
rect 34698 6060 34704 6112
rect 34756 6100 34762 6112
rect 35621 6103 35679 6109
rect 35621 6100 35633 6103
rect 34756 6072 35633 6100
rect 34756 6060 34762 6072
rect 35621 6069 35633 6072
rect 35667 6069 35679 6103
rect 35621 6063 35679 6069
rect 36170 6060 36176 6112
rect 36228 6100 36234 6112
rect 38396 6100 38424 6140
rect 41690 6128 41696 6140
rect 41748 6128 41754 6180
rect 43456 6168 43484 6208
rect 45002 6196 45008 6208
rect 45060 6196 45066 6248
rect 56134 6196 56140 6248
rect 56192 6236 56198 6248
rect 56873 6239 56931 6245
rect 56873 6236 56885 6239
rect 56192 6208 56885 6236
rect 56192 6196 56198 6208
rect 56873 6205 56885 6208
rect 56919 6205 56931 6239
rect 56873 6199 56931 6205
rect 48590 6168 48596 6180
rect 43456 6140 48596 6168
rect 48590 6128 48596 6140
rect 48648 6128 48654 6180
rect 55214 6128 55220 6180
rect 55272 6168 55278 6180
rect 58253 6171 58311 6177
rect 58253 6168 58265 6171
rect 55272 6140 58265 6168
rect 55272 6128 55278 6140
rect 58253 6137 58265 6140
rect 58299 6137 58311 6171
rect 58253 6131 58311 6137
rect 36228 6072 38424 6100
rect 36228 6060 36234 6072
rect 38470 6060 38476 6112
rect 38528 6100 38534 6112
rect 38841 6103 38899 6109
rect 38841 6100 38853 6103
rect 38528 6072 38853 6100
rect 38528 6060 38534 6072
rect 38841 6069 38853 6072
rect 38887 6069 38899 6103
rect 55766 6100 55772 6112
rect 55727 6072 55772 6100
rect 38841 6063 38899 6069
rect 55766 6060 55772 6072
rect 55824 6060 55830 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 13265 5899 13323 5905
rect 13265 5896 13277 5899
rect 11020 5868 13277 5896
rect 11020 5856 11026 5868
rect 13265 5865 13277 5868
rect 13311 5865 13323 5899
rect 13265 5859 13323 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 18966 5896 18972 5908
rect 16540 5868 18972 5896
rect 16540 5856 16546 5868
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20990 5896 20996 5908
rect 20312 5868 20996 5896
rect 20312 5856 20318 5868
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 23566 5856 23572 5908
rect 23624 5896 23630 5908
rect 24581 5899 24639 5905
rect 24581 5896 24593 5899
rect 23624 5868 24593 5896
rect 23624 5856 23630 5868
rect 24581 5865 24593 5868
rect 24627 5865 24639 5899
rect 25590 5896 25596 5908
rect 24581 5859 24639 5865
rect 25240 5868 25596 5896
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 17126 5828 17132 5840
rect 5592 5800 17132 5828
rect 5592 5788 5598 5800
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 23198 5828 23204 5840
rect 19996 5800 23204 5828
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 16114 5760 16120 5772
rect 10919 5732 16120 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 17310 5760 17316 5772
rect 16316 5732 17316 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 9214 5692 9220 5704
rect 1627 5664 9220 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 16316 5692 16344 5732
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19334 5760 19340 5772
rect 18748 5732 19340 5760
rect 18748 5720 18754 5732
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 19886 5760 19892 5772
rect 19847 5732 19892 5760
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 19996 5769 20024 5800
rect 23198 5788 23204 5800
rect 23256 5788 23262 5840
rect 23842 5788 23848 5840
rect 23900 5828 23906 5840
rect 24029 5831 24087 5837
rect 24029 5828 24041 5831
rect 23900 5800 24041 5828
rect 23900 5788 23906 5800
rect 24029 5797 24041 5800
rect 24075 5797 24087 5831
rect 24029 5791 24087 5797
rect 19981 5763 20039 5769
rect 19981 5729 19993 5763
rect 20027 5729 20039 5763
rect 20901 5763 20959 5769
rect 19981 5723 20039 5729
rect 20088 5732 20484 5760
rect 14783 5664 16344 5692
rect 16393 5695 16451 5701
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16482 5692 16488 5704
rect 16439 5664 16488 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 16850 5652 16856 5704
rect 16908 5692 16914 5704
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 16908 5664 17049 5692
rect 16908 5652 16914 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17586 5692 17592 5704
rect 17543 5664 17592 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18414 5692 18420 5704
rect 18375 5664 18420 5692
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 20088 5692 20116 5732
rect 18840 5664 20116 5692
rect 18840 5652 18846 5664
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 20312 5664 20361 5692
rect 20312 5652 20318 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20456 5692 20484 5732
rect 20901 5729 20913 5763
rect 20947 5760 20959 5763
rect 21082 5760 21088 5772
rect 20947 5732 21088 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 22830 5760 22836 5772
rect 22791 5732 22836 5760
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 25130 5720 25136 5772
rect 25188 5760 25194 5772
rect 25240 5769 25268 5868
rect 25590 5856 25596 5868
rect 25648 5896 25654 5908
rect 27062 5896 27068 5908
rect 25648 5868 27068 5896
rect 25648 5856 25654 5868
rect 27062 5856 27068 5868
rect 27120 5896 27126 5908
rect 27120 5868 27200 5896
rect 27120 5856 27126 5868
rect 26602 5828 26608 5840
rect 26563 5800 26608 5828
rect 26602 5788 26608 5800
rect 26660 5788 26666 5840
rect 27172 5769 27200 5868
rect 27338 5856 27344 5908
rect 27396 5896 27402 5908
rect 30285 5899 30343 5905
rect 27396 5868 29500 5896
rect 27396 5856 27402 5868
rect 29362 5828 29368 5840
rect 28368 5800 29368 5828
rect 25225 5763 25283 5769
rect 25225 5760 25237 5763
rect 25188 5732 25237 5760
rect 25188 5720 25194 5732
rect 25225 5729 25237 5732
rect 25271 5729 25283 5763
rect 25225 5723 25283 5729
rect 27157 5763 27215 5769
rect 27157 5729 27169 5763
rect 27203 5729 27215 5763
rect 27157 5723 27215 5729
rect 21818 5692 21824 5704
rect 20456 5664 21496 5692
rect 21779 5664 21824 5692
rect 20349 5655 20407 5661
rect 1854 5624 1860 5636
rect 1815 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 10502 5584 10508 5636
rect 10560 5624 10566 5636
rect 10689 5627 10747 5633
rect 10689 5624 10701 5627
rect 10560 5596 10701 5624
rect 10560 5584 10566 5596
rect 10689 5593 10701 5596
rect 10735 5593 10747 5627
rect 10689 5587 10747 5593
rect 11609 5627 11667 5633
rect 11609 5593 11621 5627
rect 11655 5624 11667 5627
rect 11655 5596 12020 5624
rect 11655 5593 11667 5596
rect 11609 5587 11667 5593
rect 11698 5556 11704 5568
rect 11659 5528 11704 5556
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 11992 5556 12020 5596
rect 12250 5584 12256 5636
rect 12308 5624 12314 5636
rect 12345 5627 12403 5633
rect 12345 5624 12357 5627
rect 12308 5596 12357 5624
rect 12308 5584 12314 5596
rect 12345 5593 12357 5596
rect 12391 5593 12403 5627
rect 12526 5624 12532 5636
rect 12487 5596 12532 5624
rect 12345 5587 12403 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 13136 5596 13185 5624
rect 13136 5584 13142 5596
rect 13173 5593 13185 5596
rect 13219 5593 13231 5627
rect 13173 5587 13231 5593
rect 14642 5584 14648 5636
rect 14700 5624 14706 5636
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 14700 5596 15025 5624
rect 14700 5584 14706 5596
rect 15013 5593 15025 5596
rect 15059 5593 15071 5627
rect 17770 5624 17776 5636
rect 17731 5596 17776 5624
rect 15013 5587 15071 5593
rect 17770 5584 17776 5596
rect 17828 5584 17834 5636
rect 18693 5627 18751 5633
rect 18693 5593 18705 5627
rect 18739 5593 18751 5627
rect 18693 5587 18751 5593
rect 12618 5556 12624 5568
rect 11992 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 18708 5556 18736 5587
rect 19978 5584 19984 5636
rect 20036 5624 20042 5636
rect 20441 5627 20499 5633
rect 20036 5596 20392 5624
rect 20036 5584 20042 5596
rect 20254 5556 20260 5568
rect 18708 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20364 5556 20392 5596
rect 20441 5593 20453 5627
rect 20487 5624 20499 5627
rect 21266 5624 21272 5636
rect 20487 5596 21272 5624
rect 20487 5593 20499 5596
rect 20441 5587 20499 5593
rect 21266 5584 21272 5596
rect 21324 5584 21330 5636
rect 21468 5624 21496 5664
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 22066 5664 23673 5692
rect 22066 5624 22094 5664
rect 23661 5661 23673 5664
rect 23707 5692 23719 5695
rect 24302 5692 24308 5704
rect 23707 5664 24308 5692
rect 23707 5661 23719 5664
rect 23661 5655 23719 5661
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24394 5652 24400 5704
rect 24452 5692 24458 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 24452 5664 24593 5692
rect 24452 5652 24458 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24728 5664 24777 5692
rect 24728 5652 24734 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 28368 5692 28396 5800
rect 29362 5788 29368 5800
rect 29420 5788 29426 5840
rect 29472 5828 29500 5868
rect 30285 5865 30297 5899
rect 30331 5896 30343 5899
rect 37642 5896 37648 5908
rect 30331 5868 36216 5896
rect 30331 5865 30343 5868
rect 30285 5859 30343 5865
rect 31478 5828 31484 5840
rect 29472 5800 31484 5828
rect 31478 5788 31484 5800
rect 31536 5788 31542 5840
rect 32033 5831 32091 5837
rect 31772 5800 31984 5828
rect 28442 5720 28448 5772
rect 28500 5760 28506 5772
rect 28500 5732 29316 5760
rect 28500 5720 28506 5732
rect 28994 5692 29000 5704
rect 24765 5655 24823 5661
rect 27356 5664 28396 5692
rect 28955 5664 29000 5692
rect 21468 5596 22094 5624
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 23845 5627 23903 5633
rect 23845 5624 23857 5627
rect 23532 5596 23857 5624
rect 23532 5584 23538 5596
rect 23845 5593 23857 5596
rect 23891 5593 23903 5627
rect 23845 5587 23903 5593
rect 24854 5584 24860 5636
rect 24912 5624 24918 5636
rect 25470 5627 25528 5633
rect 25470 5624 25482 5627
rect 24912 5596 25482 5624
rect 24912 5584 24918 5596
rect 25470 5593 25482 5596
rect 25516 5593 25528 5627
rect 25470 5587 25528 5593
rect 25590 5584 25596 5636
rect 25648 5624 25654 5636
rect 27356 5624 27384 5664
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 29178 5692 29184 5704
rect 29139 5664 29184 5692
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 29288 5692 29316 5732
rect 29730 5720 29736 5772
rect 29788 5760 29794 5772
rect 30466 5760 30472 5772
rect 29788 5732 30472 5760
rect 29788 5720 29794 5732
rect 30466 5720 30472 5732
rect 30524 5760 30530 5772
rect 30929 5763 30987 5769
rect 30929 5760 30941 5763
rect 30524 5732 30941 5760
rect 30524 5720 30530 5732
rect 30929 5729 30941 5732
rect 30975 5760 30987 5763
rect 31772 5760 31800 5800
rect 30975 5732 31800 5760
rect 31956 5760 31984 5800
rect 32033 5797 32045 5831
rect 32079 5828 32091 5831
rect 33226 5828 33232 5840
rect 32079 5800 33232 5828
rect 32079 5797 32091 5800
rect 32033 5791 32091 5797
rect 33226 5788 33232 5800
rect 33284 5788 33290 5840
rect 33318 5788 33324 5840
rect 33376 5828 33382 5840
rect 33505 5831 33563 5837
rect 33505 5828 33517 5831
rect 33376 5800 33517 5828
rect 33376 5788 33382 5800
rect 33505 5797 33517 5800
rect 33551 5797 33563 5831
rect 33505 5791 33563 5797
rect 34974 5788 34980 5840
rect 35032 5828 35038 5840
rect 35618 5828 35624 5840
rect 35032 5800 35624 5828
rect 35032 5788 35038 5800
rect 35618 5788 35624 5800
rect 35676 5788 35682 5840
rect 32677 5763 32735 5769
rect 32677 5760 32689 5763
rect 31956 5732 32689 5760
rect 30975 5729 30987 5732
rect 30929 5723 30987 5729
rect 32677 5729 32689 5732
rect 32723 5760 32735 5763
rect 35526 5760 35532 5772
rect 32723 5732 35532 5760
rect 32723 5729 32735 5732
rect 32677 5723 32735 5729
rect 35526 5720 35532 5732
rect 35584 5720 35590 5772
rect 35894 5720 35900 5772
rect 35952 5760 35958 5772
rect 35989 5763 36047 5769
rect 35989 5760 36001 5763
rect 35952 5732 36001 5760
rect 35952 5720 35958 5732
rect 35989 5729 36001 5732
rect 36035 5729 36047 5763
rect 35989 5723 36047 5729
rect 29288 5664 30880 5692
rect 25648 5596 27384 5624
rect 27424 5627 27482 5633
rect 25648 5584 25654 5596
rect 27424 5593 27436 5627
rect 27470 5624 27482 5627
rect 27706 5624 27712 5636
rect 27470 5596 27712 5624
rect 27470 5593 27482 5596
rect 27424 5587 27482 5593
rect 27706 5584 27712 5596
rect 27764 5584 27770 5636
rect 27798 5584 27804 5636
rect 27856 5624 27862 5636
rect 28074 5624 28080 5636
rect 27856 5596 28080 5624
rect 27856 5584 27862 5596
rect 28074 5584 28080 5596
rect 28132 5624 28138 5636
rect 30745 5627 30803 5633
rect 30745 5624 30757 5627
rect 28132 5596 30757 5624
rect 28132 5584 28138 5596
rect 30745 5593 30757 5596
rect 30791 5593 30803 5627
rect 30852 5624 30880 5664
rect 31018 5652 31024 5704
rect 31076 5692 31082 5704
rect 33229 5695 33287 5701
rect 33229 5692 33241 5695
rect 31076 5664 33241 5692
rect 31076 5652 31082 5664
rect 33229 5661 33241 5664
rect 33275 5661 33287 5695
rect 33229 5655 33287 5661
rect 33410 5652 33416 5704
rect 33468 5692 33474 5704
rect 34974 5692 34980 5704
rect 33468 5664 34980 5692
rect 33468 5652 33474 5664
rect 34974 5652 34980 5664
rect 35032 5652 35038 5704
rect 36188 5701 36216 5868
rect 36832 5868 37648 5896
rect 36832 5769 36860 5868
rect 37642 5856 37648 5868
rect 37700 5856 37706 5908
rect 37737 5899 37795 5905
rect 37737 5865 37749 5899
rect 37783 5896 37795 5899
rect 37826 5896 37832 5908
rect 37783 5868 37832 5896
rect 37783 5865 37795 5868
rect 37737 5859 37795 5865
rect 37826 5856 37832 5868
rect 37884 5856 37890 5908
rect 38746 5856 38752 5908
rect 38804 5896 38810 5908
rect 39114 5896 39120 5908
rect 38804 5868 39120 5896
rect 38804 5856 38810 5868
rect 39114 5856 39120 5868
rect 39172 5856 39178 5908
rect 41690 5896 41696 5908
rect 41651 5868 41696 5896
rect 41690 5856 41696 5868
rect 41748 5856 41754 5908
rect 43714 5856 43720 5908
rect 43772 5896 43778 5908
rect 44545 5899 44603 5905
rect 44545 5896 44557 5899
rect 43772 5868 44557 5896
rect 43772 5856 43778 5868
rect 44545 5865 44557 5868
rect 44591 5865 44603 5899
rect 45278 5896 45284 5908
rect 45239 5868 45284 5896
rect 44545 5859 44603 5865
rect 45278 5856 45284 5868
rect 45336 5856 45342 5908
rect 53926 5828 53932 5840
rect 36924 5800 53932 5828
rect 36817 5763 36875 5769
rect 36817 5729 36829 5763
rect 36863 5729 36875 5763
rect 36817 5723 36875 5729
rect 35069 5695 35127 5701
rect 35069 5661 35081 5695
rect 35115 5692 35127 5695
rect 36173 5695 36231 5701
rect 35115 5664 35940 5692
rect 35115 5661 35127 5664
rect 35069 5655 35127 5661
rect 31662 5624 31668 5636
rect 30852 5596 31668 5624
rect 30745 5587 30803 5593
rect 31662 5584 31668 5596
rect 31720 5584 31726 5636
rect 31846 5584 31852 5636
rect 31904 5624 31910 5636
rect 34149 5627 34207 5633
rect 34149 5624 34161 5627
rect 31904 5596 34161 5624
rect 31904 5584 31910 5596
rect 34149 5593 34161 5596
rect 34195 5593 34207 5627
rect 34149 5587 34207 5593
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 35345 5627 35403 5633
rect 35345 5624 35357 5627
rect 34572 5596 35357 5624
rect 34572 5584 34578 5596
rect 35345 5593 35357 5596
rect 35391 5593 35403 5627
rect 35912 5624 35940 5664
rect 36173 5661 36185 5695
rect 36219 5661 36231 5695
rect 36173 5655 36231 5661
rect 36262 5652 36268 5704
rect 36320 5692 36326 5704
rect 36924 5692 36952 5800
rect 53926 5788 53932 5800
rect 53984 5788 53990 5840
rect 37090 5760 37096 5772
rect 37016 5732 37096 5760
rect 37016 5701 37044 5732
rect 37090 5720 37096 5732
rect 37148 5720 37154 5772
rect 37366 5720 37372 5772
rect 37424 5760 37430 5772
rect 38197 5763 38255 5769
rect 38197 5760 38209 5763
rect 37424 5732 38209 5760
rect 37424 5720 37430 5732
rect 38197 5729 38209 5732
rect 38243 5729 38255 5763
rect 38197 5723 38255 5729
rect 38378 5720 38384 5772
rect 38436 5760 38442 5772
rect 43165 5763 43223 5769
rect 43165 5760 43177 5763
rect 38436 5732 43177 5760
rect 38436 5720 38442 5732
rect 43165 5729 43177 5732
rect 43211 5729 43223 5763
rect 43714 5760 43720 5772
rect 43165 5723 43223 5729
rect 43272 5732 43720 5760
rect 36320 5664 36952 5692
rect 37001 5695 37059 5701
rect 36320 5652 36326 5664
rect 37001 5661 37013 5695
rect 37047 5661 37059 5695
rect 40402 5692 40408 5704
rect 37001 5655 37059 5661
rect 37108 5664 40408 5692
rect 37108 5624 37136 5664
rect 40402 5652 40408 5664
rect 40460 5652 40466 5704
rect 40862 5652 40868 5704
rect 40920 5692 40926 5704
rect 42429 5695 42487 5701
rect 42429 5692 42441 5695
rect 40920 5664 42441 5692
rect 40920 5652 40926 5664
rect 42429 5661 42441 5664
rect 42475 5661 42487 5695
rect 42429 5655 42487 5661
rect 42705 5695 42763 5701
rect 42705 5661 42717 5695
rect 42751 5692 42763 5695
rect 42794 5692 42800 5704
rect 42751 5664 42800 5692
rect 42751 5661 42763 5664
rect 42705 5655 42763 5661
rect 38470 5624 38476 5636
rect 35912 5596 37136 5624
rect 38120 5596 38476 5624
rect 35345 5587 35403 5593
rect 20898 5556 20904 5568
rect 20364 5528 20904 5556
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 26142 5556 26148 5568
rect 22152 5528 26148 5556
rect 22152 5516 22158 5528
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 28166 5516 28172 5568
rect 28224 5556 28230 5568
rect 28537 5559 28595 5565
rect 28537 5556 28549 5559
rect 28224 5528 28549 5556
rect 28224 5516 28230 5528
rect 28537 5525 28549 5528
rect 28583 5525 28595 5559
rect 28537 5519 28595 5525
rect 28718 5516 28724 5568
rect 28776 5556 28782 5568
rect 29089 5559 29147 5565
rect 29089 5556 29101 5559
rect 28776 5528 29101 5556
rect 28776 5516 28782 5528
rect 29089 5525 29101 5528
rect 29135 5525 29147 5559
rect 30650 5556 30656 5568
rect 30611 5528 30656 5556
rect 29089 5519 29147 5525
rect 30650 5516 30656 5528
rect 30708 5516 30714 5568
rect 31478 5516 31484 5568
rect 31536 5556 31542 5568
rect 32214 5556 32220 5568
rect 31536 5528 32220 5556
rect 31536 5516 31542 5528
rect 32214 5516 32220 5528
rect 32272 5516 32278 5568
rect 32398 5556 32404 5568
rect 32359 5528 32404 5556
rect 32398 5516 32404 5528
rect 32456 5516 32462 5568
rect 32493 5559 32551 5565
rect 32493 5525 32505 5559
rect 32539 5556 32551 5559
rect 32582 5556 32588 5568
rect 32539 5528 32588 5556
rect 32539 5525 32551 5528
rect 32493 5519 32551 5525
rect 32582 5516 32588 5528
rect 32640 5516 32646 5568
rect 33410 5516 33416 5568
rect 33468 5556 33474 5568
rect 33689 5559 33747 5565
rect 33689 5556 33701 5559
rect 33468 5528 33701 5556
rect 33468 5516 33474 5528
rect 33689 5525 33701 5528
rect 33735 5525 33747 5559
rect 33689 5519 33747 5525
rect 34606 5516 34612 5568
rect 34664 5556 34670 5568
rect 36357 5559 36415 5565
rect 36357 5556 36369 5559
rect 34664 5528 36369 5556
rect 34664 5516 34670 5528
rect 36357 5525 36369 5528
rect 36403 5525 36415 5559
rect 37182 5556 37188 5568
rect 37143 5528 37188 5556
rect 36357 5519 36415 5525
rect 37182 5516 37188 5528
rect 37240 5516 37246 5568
rect 37826 5516 37832 5568
rect 37884 5556 37890 5568
rect 38120 5565 38148 5596
rect 38470 5584 38476 5596
rect 38528 5584 38534 5636
rect 38930 5584 38936 5636
rect 38988 5624 38994 5636
rect 39025 5627 39083 5633
rect 39025 5624 39037 5627
rect 38988 5596 39037 5624
rect 38988 5584 38994 5596
rect 39025 5593 39037 5596
rect 39071 5593 39083 5627
rect 41598 5624 41604 5636
rect 41559 5596 41604 5624
rect 39025 5587 39083 5593
rect 41598 5584 41604 5596
rect 41656 5584 41662 5636
rect 38105 5559 38163 5565
rect 38105 5556 38117 5559
rect 37884 5528 38117 5556
rect 37884 5516 37890 5528
rect 38105 5525 38117 5528
rect 38151 5525 38163 5559
rect 38105 5519 38163 5525
rect 38194 5516 38200 5568
rect 38252 5556 38258 5568
rect 39117 5559 39175 5565
rect 39117 5556 39129 5559
rect 38252 5528 39129 5556
rect 38252 5516 38258 5528
rect 39117 5525 39129 5528
rect 39163 5525 39175 5559
rect 42444 5556 42472 5655
rect 42794 5652 42800 5664
rect 42852 5652 42858 5704
rect 42886 5652 42892 5704
rect 42944 5692 42950 5704
rect 43272 5692 43300 5732
rect 43714 5720 43720 5732
rect 43772 5720 43778 5772
rect 56870 5760 56876 5772
rect 56831 5732 56876 5760
rect 56870 5720 56876 5732
rect 56928 5720 56934 5772
rect 45189 5695 45247 5701
rect 45189 5692 45201 5695
rect 42944 5664 43300 5692
rect 43640 5664 45201 5692
rect 42944 5652 42950 5664
rect 42613 5627 42671 5633
rect 42613 5593 42625 5627
rect 42659 5624 42671 5627
rect 43640 5624 43668 5664
rect 45189 5661 45201 5664
rect 45235 5692 45247 5695
rect 45235 5664 51074 5692
rect 45235 5661 45247 5664
rect 45189 5655 45247 5661
rect 42659 5596 43668 5624
rect 42659 5593 42671 5596
rect 42613 5587 42671 5593
rect 43714 5584 43720 5636
rect 43772 5624 43778 5636
rect 43772 5596 43817 5624
rect 43772 5584 43778 5596
rect 44358 5584 44364 5636
rect 44416 5624 44422 5636
rect 44453 5627 44511 5633
rect 44453 5624 44465 5627
rect 44416 5596 44465 5624
rect 44416 5584 44422 5596
rect 44453 5593 44465 5596
rect 44499 5593 44511 5627
rect 51046 5624 51074 5664
rect 55766 5652 55772 5704
rect 55824 5692 55830 5704
rect 57129 5695 57187 5701
rect 57129 5692 57141 5695
rect 55824 5664 57141 5692
rect 55824 5652 55830 5664
rect 57129 5661 57141 5664
rect 57175 5661 57187 5695
rect 57129 5655 57187 5661
rect 58342 5624 58348 5636
rect 51046 5596 58348 5624
rect 44453 5587 44511 5593
rect 58342 5584 58348 5596
rect 58400 5584 58406 5636
rect 43438 5556 43444 5568
rect 42444 5528 43444 5556
rect 39117 5519 39175 5525
rect 43438 5516 43444 5528
rect 43496 5516 43502 5568
rect 43806 5556 43812 5568
rect 43767 5528 43812 5556
rect 43806 5516 43812 5528
rect 43864 5516 43870 5568
rect 57330 5516 57336 5568
rect 57388 5556 57394 5568
rect 58253 5559 58311 5565
rect 58253 5556 58265 5559
rect 57388 5528 58265 5556
rect 57388 5516 57394 5528
rect 58253 5525 58265 5528
rect 58299 5525 58311 5559
rect 58253 5519 58311 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 9582 5352 9588 5364
rect 9543 5324 9588 5352
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 9858 5352 9864 5364
rect 9771 5324 9864 5352
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 8386 5216 8392 5228
rect 1627 5188 8392 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8628 5188 8769 5216
rect 8628 5176 8634 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9784 5225 9812 5324
rect 9858 5312 9864 5324
rect 9916 5352 9922 5364
rect 23750 5352 23756 5364
rect 9916 5324 23756 5352
rect 9916 5312 9922 5324
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 23937 5355 23995 5361
rect 23937 5321 23949 5355
rect 23983 5352 23995 5355
rect 24854 5352 24860 5364
rect 23983 5324 24860 5352
rect 23983 5321 23995 5324
rect 23937 5315 23995 5321
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 27706 5352 27712 5364
rect 27667 5324 27712 5352
rect 27706 5312 27712 5324
rect 27764 5312 27770 5364
rect 28074 5352 28080 5364
rect 28035 5324 28080 5352
rect 28074 5312 28080 5324
rect 28132 5312 28138 5364
rect 28997 5355 29055 5361
rect 28997 5321 29009 5355
rect 29043 5352 29055 5355
rect 31478 5352 31484 5364
rect 29043 5324 31484 5352
rect 29043 5321 29055 5324
rect 28997 5315 29055 5321
rect 31478 5312 31484 5324
rect 31536 5312 31542 5364
rect 31680 5324 34468 5352
rect 10594 5284 10600 5296
rect 9876 5256 10600 5284
rect 9876 5225 9904 5256
rect 10594 5244 10600 5256
rect 10652 5244 10658 5296
rect 11149 5287 11207 5293
rect 11149 5253 11161 5287
rect 11195 5284 11207 5287
rect 11238 5284 11244 5296
rect 11195 5256 11244 5284
rect 11195 5253 11207 5256
rect 11149 5247 11207 5253
rect 11238 5244 11244 5256
rect 11296 5244 11302 5296
rect 11974 5244 11980 5296
rect 12032 5284 12038 5296
rect 15838 5284 15844 5296
rect 12032 5256 14044 5284
rect 15799 5256 15844 5284
rect 12032 5244 12038 5256
rect 9769 5219 9827 5225
rect 9088 5188 9674 5216
rect 9088 5176 9094 5188
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 9646 5080 9674 5188
rect 9769 5185 9781 5219
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 9861 5179 9919 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10836 5188 10977 5216
rect 10836 5176 10842 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11848 5188 11897 5216
rect 11848 5176 11854 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 13814 5216 13820 5228
rect 13403 5188 13820 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5148 10011 5151
rect 10318 5148 10324 5160
rect 9999 5120 10324 5148
rect 9999 5117 10011 5120
rect 9953 5111 10011 5117
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12360 5148 12388 5179
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 14016 5225 14044 5256
rect 15838 5244 15844 5256
rect 15896 5284 15902 5296
rect 18509 5287 18567 5293
rect 18509 5284 18521 5287
rect 15896 5256 18521 5284
rect 15896 5244 15902 5256
rect 18509 5253 18521 5256
rect 18555 5253 18567 5287
rect 18509 5247 18567 5253
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 24026 5284 24032 5296
rect 19392 5256 24032 5284
rect 19392 5244 19398 5256
rect 24026 5244 24032 5256
rect 24084 5244 24090 5296
rect 24946 5244 24952 5296
rect 25004 5284 25010 5296
rect 25378 5287 25436 5293
rect 25378 5284 25390 5287
rect 25004 5256 25390 5284
rect 25004 5244 25010 5256
rect 25378 5253 25390 5256
rect 25424 5253 25436 5287
rect 25378 5247 25436 5253
rect 28718 5244 28724 5296
rect 28776 5284 28782 5296
rect 28776 5256 30144 5284
rect 28776 5244 28782 5256
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 16942 5216 16948 5228
rect 14148 5188 16252 5216
rect 16903 5188 16948 5216
rect 14148 5176 14154 5188
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 11388 5120 14749 5148
rect 11388 5108 11394 5120
rect 10042 5080 10048 5092
rect 7616 5052 8984 5080
rect 9646 5052 10048 5080
rect 7616 5040 7622 5052
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8536 4984 8861 5012
rect 8536 4972 8542 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 8956 5012 8984 5052
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 12621 5083 12679 5089
rect 12621 5080 12633 5083
rect 11480 5052 12633 5080
rect 11480 5040 11486 5052
rect 12621 5049 12633 5052
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 12158 5012 12164 5024
rect 8956 4984 12164 5012
rect 8849 4975 8907 4981
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12805 5015 12863 5021
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 13354 5012 13360 5024
rect 12851 4984 13360 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13464 5012 13492 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 13541 5083 13599 5089
rect 13541 5049 13553 5083
rect 13587 5080 13599 5083
rect 15013 5083 15071 5089
rect 15013 5080 15025 5083
rect 13587 5052 15025 5080
rect 13587 5049 13599 5052
rect 13541 5043 13599 5049
rect 15013 5049 15025 5052
rect 15059 5049 15071 5083
rect 16114 5080 16120 5092
rect 16075 5052 16120 5080
rect 15013 5043 15071 5049
rect 16114 5040 16120 5052
rect 16172 5040 16178 5092
rect 16224 5080 16252 5188
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 17083 5188 17601 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17589 5185 17601 5188
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 19242 5216 19248 5228
rect 17911 5188 19248 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 19426 5216 19432 5228
rect 19387 5188 19432 5216
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5216 19763 5219
rect 19978 5216 19984 5228
rect 19751 5188 19984 5216
rect 19751 5185 19763 5188
rect 19705 5179 19763 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20622 5216 20628 5228
rect 20487 5188 20628 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 20622 5176 20628 5188
rect 20680 5216 20686 5228
rect 21818 5216 21824 5228
rect 20680 5188 21824 5216
rect 20680 5176 20686 5188
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22462 5216 22468 5228
rect 22235 5188 22468 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22830 5216 22836 5228
rect 22791 5188 22836 5216
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 24305 5219 24363 5225
rect 24305 5216 24317 5219
rect 23952 5188 24317 5216
rect 16301 5151 16359 5157
rect 16301 5117 16313 5151
rect 16347 5148 16359 5151
rect 16758 5148 16764 5160
rect 16347 5120 16764 5148
rect 16347 5117 16359 5120
rect 16301 5111 16359 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 18966 5148 18972 5160
rect 18927 5120 18972 5148
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 20806 5148 20812 5160
rect 19116 5120 20812 5148
rect 19116 5108 19122 5120
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 18785 5083 18843 5089
rect 18785 5080 18797 5083
rect 16224 5052 18797 5080
rect 18785 5049 18797 5052
rect 18831 5049 18843 5083
rect 19150 5080 19156 5092
rect 18785 5043 18843 5049
rect 18892 5052 19156 5080
rect 14185 5015 14243 5021
rect 14185 5012 14197 5015
rect 13464 4984 14197 5012
rect 14185 4981 14197 4984
rect 14231 4981 14243 5015
rect 14185 4975 14243 4981
rect 15197 5015 15255 5021
rect 15197 4981 15209 5015
rect 15243 5012 15255 5015
rect 18892 5012 18920 5052
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 19242 5040 19248 5092
rect 19300 5080 19306 5092
rect 20254 5080 20260 5092
rect 19300 5052 20260 5080
rect 19300 5040 19306 5052
rect 20254 5040 20260 5052
rect 20312 5040 20318 5092
rect 20824 5080 20852 5108
rect 23952 5080 23980 5188
rect 24305 5185 24317 5188
rect 24351 5216 24363 5219
rect 24486 5216 24492 5228
rect 24351 5188 24492 5216
rect 24351 5185 24363 5188
rect 24305 5179 24363 5185
rect 24486 5176 24492 5188
rect 24544 5176 24550 5228
rect 25130 5216 25136 5228
rect 25091 5188 25136 5216
rect 25130 5176 25136 5188
rect 25188 5176 25194 5228
rect 28258 5176 28264 5228
rect 28316 5216 28322 5228
rect 28902 5216 28908 5228
rect 28316 5188 28908 5216
rect 28316 5176 28322 5188
rect 28902 5176 28908 5188
rect 28960 5176 28966 5228
rect 29089 5219 29147 5225
rect 29089 5185 29101 5219
rect 29135 5216 29147 5219
rect 29178 5216 29184 5228
rect 29135 5188 29184 5216
rect 29135 5185 29147 5188
rect 29089 5179 29147 5185
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 29546 5216 29552 5228
rect 29507 5188 29552 5216
rect 29546 5176 29552 5188
rect 29604 5176 29610 5228
rect 29822 5225 29828 5228
rect 29816 5179 29828 5225
rect 29880 5216 29886 5228
rect 30116 5216 30144 5256
rect 30190 5244 30196 5296
rect 30248 5284 30254 5296
rect 31018 5284 31024 5296
rect 30248 5256 31024 5284
rect 30248 5244 30254 5256
rect 31018 5244 31024 5256
rect 31076 5244 31082 5296
rect 31680 5284 31708 5324
rect 34440 5293 34468 5324
rect 35342 5312 35348 5364
rect 35400 5352 35406 5364
rect 36078 5352 36084 5364
rect 35400 5324 36084 5352
rect 35400 5312 35406 5324
rect 36078 5312 36084 5324
rect 36136 5312 36142 5364
rect 36446 5312 36452 5364
rect 36504 5352 36510 5364
rect 38470 5352 38476 5364
rect 36504 5324 38476 5352
rect 36504 5312 36510 5324
rect 38470 5312 38476 5324
rect 38528 5312 38534 5364
rect 38562 5312 38568 5364
rect 38620 5352 38626 5364
rect 40589 5355 40647 5361
rect 40589 5352 40601 5355
rect 38620 5324 40601 5352
rect 38620 5312 38626 5324
rect 40589 5321 40601 5324
rect 40635 5321 40647 5355
rect 40589 5315 40647 5321
rect 40770 5312 40776 5364
rect 40828 5352 40834 5364
rect 43346 5352 43352 5364
rect 40828 5324 43352 5352
rect 40828 5312 40834 5324
rect 43346 5312 43352 5324
rect 43404 5312 43410 5364
rect 43530 5352 43536 5364
rect 43491 5324 43536 5352
rect 43530 5312 43536 5324
rect 43588 5312 43594 5364
rect 45002 5352 45008 5364
rect 44963 5324 45008 5352
rect 45002 5312 45008 5324
rect 45060 5352 45066 5364
rect 45370 5352 45376 5364
rect 45060 5324 45376 5352
rect 45060 5312 45066 5324
rect 45370 5312 45376 5324
rect 45428 5312 45434 5364
rect 57238 5352 57244 5364
rect 57199 5324 57244 5352
rect 57238 5312 57244 5324
rect 57296 5312 57302 5364
rect 34425 5287 34483 5293
rect 31128 5256 31708 5284
rect 32324 5256 34192 5284
rect 31128 5216 31156 5256
rect 29880 5188 29916 5216
rect 30116 5188 31156 5216
rect 31573 5219 31631 5225
rect 29822 5176 29828 5179
rect 29880 5176 29886 5188
rect 31573 5185 31585 5219
rect 31619 5216 31631 5219
rect 31754 5216 31760 5228
rect 31619 5188 31760 5216
rect 31619 5185 31631 5188
rect 31573 5179 31631 5185
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 32324 5225 32352 5256
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31904 5188 32321 5216
rect 31904 5176 31910 5188
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 33505 5219 33563 5225
rect 33505 5216 33517 5219
rect 32309 5179 32367 5185
rect 33428 5188 33517 5216
rect 24394 5148 24400 5160
rect 24355 5120 24400 5148
rect 24394 5108 24400 5120
rect 24452 5108 24458 5160
rect 24581 5151 24639 5157
rect 24581 5117 24593 5151
rect 24627 5148 24639 5151
rect 24670 5148 24676 5160
rect 24627 5120 24676 5148
rect 24627 5117 24639 5120
rect 24581 5111 24639 5117
rect 24670 5108 24676 5120
rect 24728 5108 24734 5160
rect 28166 5148 28172 5160
rect 28127 5120 28172 5148
rect 28166 5108 28172 5120
rect 28224 5108 28230 5160
rect 28353 5151 28411 5157
rect 28353 5117 28365 5151
rect 28399 5148 28411 5151
rect 28626 5148 28632 5160
rect 28399 5120 28632 5148
rect 28399 5117 28411 5120
rect 28353 5111 28411 5117
rect 20824 5052 23980 5080
rect 27890 5040 27896 5092
rect 27948 5080 27954 5092
rect 28368 5080 28396 5111
rect 28626 5108 28632 5120
rect 28684 5148 28690 5160
rect 29454 5148 29460 5160
rect 28684 5120 29460 5148
rect 28684 5108 28690 5120
rect 29454 5108 29460 5120
rect 29512 5108 29518 5160
rect 31386 5148 31392 5160
rect 31347 5120 31392 5148
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 31938 5108 31944 5160
rect 31996 5148 32002 5160
rect 32401 5151 32459 5157
rect 32401 5148 32413 5151
rect 31996 5120 32413 5148
rect 31996 5108 32002 5120
rect 32401 5117 32413 5120
rect 32447 5117 32459 5151
rect 32401 5111 32459 5117
rect 33428 5148 33456 5188
rect 33505 5185 33517 5188
rect 33551 5185 33563 5219
rect 33505 5179 33563 5185
rect 33689 5219 33747 5225
rect 33689 5185 33701 5219
rect 33735 5216 33747 5219
rect 33778 5216 33784 5228
rect 33735 5188 33784 5216
rect 33735 5185 33747 5188
rect 33689 5179 33747 5185
rect 33778 5176 33784 5188
rect 33836 5176 33842 5228
rect 34164 5225 34192 5256
rect 34425 5253 34437 5287
rect 34471 5253 34483 5287
rect 36357 5287 36415 5293
rect 36357 5284 36369 5287
rect 34425 5247 34483 5253
rect 34532 5256 36369 5284
rect 34149 5219 34207 5225
rect 34149 5185 34161 5219
rect 34195 5185 34207 5219
rect 34149 5179 34207 5185
rect 34238 5176 34244 5228
rect 34296 5216 34302 5228
rect 34532 5216 34560 5256
rect 36357 5253 36369 5256
rect 36403 5253 36415 5287
rect 36357 5247 36415 5253
rect 37553 5287 37611 5293
rect 37553 5253 37565 5287
rect 37599 5284 37611 5287
rect 38654 5284 38660 5296
rect 37599 5256 38660 5284
rect 37599 5253 37611 5256
rect 37553 5247 37611 5253
rect 38654 5244 38660 5256
rect 38712 5284 38718 5296
rect 39025 5287 39083 5293
rect 39025 5284 39037 5287
rect 38712 5256 39037 5284
rect 38712 5244 38718 5256
rect 39025 5253 39037 5256
rect 39071 5253 39083 5287
rect 39945 5287 40003 5293
rect 39945 5284 39957 5287
rect 39025 5247 39083 5253
rect 39132 5256 39957 5284
rect 35066 5216 35072 5228
rect 34296 5188 34560 5216
rect 35027 5188 35072 5216
rect 34296 5176 34302 5188
rect 35066 5176 35072 5188
rect 35124 5176 35130 5228
rect 35802 5216 35808 5228
rect 35232 5188 35808 5216
rect 34054 5148 34060 5160
rect 33428 5120 34060 5148
rect 27948 5052 28396 5080
rect 27948 5040 27954 5052
rect 30558 5040 30564 5092
rect 30616 5080 30622 5092
rect 31110 5080 31116 5092
rect 30616 5052 31116 5080
rect 30616 5040 30622 5052
rect 31110 5040 31116 5052
rect 31168 5040 31174 5092
rect 31478 5040 31484 5092
rect 31536 5080 31542 5092
rect 31757 5083 31815 5089
rect 31757 5080 31769 5083
rect 31536 5052 31769 5080
rect 31536 5040 31542 5052
rect 31757 5049 31769 5052
rect 31803 5049 31815 5083
rect 31757 5043 31815 5049
rect 32030 5040 32036 5092
rect 32088 5080 32094 5092
rect 33428 5080 33456 5120
rect 34054 5108 34060 5120
rect 34112 5148 34118 5160
rect 35232 5148 35260 5188
rect 35802 5176 35808 5188
rect 35860 5176 35866 5228
rect 36170 5216 36176 5228
rect 36131 5188 36176 5216
rect 36170 5176 36176 5188
rect 36228 5176 36234 5228
rect 38286 5216 38292 5228
rect 38247 5188 38292 5216
rect 38286 5176 38292 5188
rect 38344 5176 38350 5228
rect 38562 5176 38568 5228
rect 38620 5216 38626 5228
rect 39132 5216 39160 5256
rect 39945 5253 39957 5256
rect 39991 5253 40003 5287
rect 39945 5247 40003 5253
rect 40310 5244 40316 5296
rect 40368 5284 40374 5296
rect 41233 5287 41291 5293
rect 41233 5284 41245 5287
rect 40368 5256 41245 5284
rect 40368 5244 40374 5256
rect 41233 5253 41245 5256
rect 41279 5253 41291 5287
rect 41233 5247 41291 5253
rect 41417 5287 41475 5293
rect 41417 5253 41429 5287
rect 41463 5284 41475 5287
rect 41506 5284 41512 5296
rect 41463 5256 41512 5284
rect 41463 5253 41475 5256
rect 41417 5247 41475 5253
rect 41506 5244 41512 5256
rect 41564 5244 41570 5296
rect 43548 5256 51074 5284
rect 43548 5228 43576 5256
rect 38620 5188 39160 5216
rect 38620 5176 38626 5188
rect 39574 5176 39580 5228
rect 39632 5216 39638 5228
rect 39761 5219 39819 5225
rect 39761 5216 39773 5219
rect 39632 5188 39773 5216
rect 39632 5176 39638 5188
rect 39761 5185 39773 5188
rect 39807 5185 39819 5219
rect 40494 5216 40500 5228
rect 40455 5188 40500 5216
rect 39761 5179 39819 5185
rect 40494 5176 40500 5188
rect 40552 5176 40558 5228
rect 41690 5176 41696 5228
rect 41748 5216 41754 5228
rect 42705 5219 42763 5225
rect 42705 5216 42717 5219
rect 41748 5188 42717 5216
rect 41748 5176 41754 5188
rect 42705 5185 42717 5188
rect 42751 5185 42763 5219
rect 42705 5179 42763 5185
rect 43349 5219 43407 5225
rect 43349 5185 43361 5219
rect 43395 5185 43407 5219
rect 43349 5179 43407 5185
rect 35342 5148 35348 5160
rect 34112 5120 35260 5148
rect 35303 5120 35348 5148
rect 34112 5108 34118 5120
rect 35342 5108 35348 5120
rect 35400 5108 35406 5160
rect 35894 5108 35900 5160
rect 35952 5148 35958 5160
rect 35989 5151 36047 5157
rect 35989 5148 36001 5151
rect 35952 5120 36001 5148
rect 35952 5108 35958 5120
rect 35989 5117 36001 5120
rect 36035 5117 36047 5151
rect 35989 5111 36047 5117
rect 37366 5108 37372 5160
rect 37424 5148 37430 5160
rect 38473 5151 38531 5157
rect 38473 5148 38485 5151
rect 37424 5120 38485 5148
rect 37424 5108 37430 5120
rect 38473 5117 38485 5120
rect 38519 5117 38531 5151
rect 38473 5111 38531 5117
rect 40126 5108 40132 5160
rect 40184 5148 40190 5160
rect 43364 5148 43392 5179
rect 43530 5176 43536 5228
rect 43588 5176 43594 5228
rect 44818 5216 44824 5228
rect 44731 5188 44824 5216
rect 44818 5176 44824 5188
rect 44876 5216 44882 5228
rect 45278 5216 45284 5228
rect 44876 5188 45284 5216
rect 44876 5176 44882 5188
rect 45278 5176 45284 5188
rect 45336 5176 45342 5228
rect 45646 5216 45652 5228
rect 45607 5188 45652 5216
rect 45646 5176 45652 5188
rect 45704 5176 45710 5228
rect 45738 5176 45744 5228
rect 45796 5216 45802 5228
rect 46569 5219 46627 5225
rect 46569 5216 46581 5219
rect 45796 5188 46581 5216
rect 45796 5176 45802 5188
rect 46569 5185 46581 5188
rect 46615 5185 46627 5219
rect 51046 5216 51074 5256
rect 53190 5216 53196 5228
rect 51046 5188 53196 5216
rect 46569 5179 46627 5185
rect 53190 5176 53196 5188
rect 53248 5176 53254 5228
rect 57146 5216 57152 5228
rect 57107 5188 57152 5216
rect 57146 5176 57152 5188
rect 57204 5176 57210 5228
rect 57330 5216 57336 5228
rect 57291 5188 57336 5216
rect 57330 5176 57336 5188
rect 57388 5176 57394 5228
rect 58066 5216 58072 5228
rect 58027 5188 58072 5216
rect 58066 5176 58072 5188
rect 58124 5176 58130 5228
rect 40184 5120 43392 5148
rect 44637 5151 44695 5157
rect 40184 5108 40190 5120
rect 44637 5117 44649 5151
rect 44683 5148 44695 5151
rect 44910 5148 44916 5160
rect 44683 5120 44916 5148
rect 44683 5117 44695 5120
rect 44637 5111 44695 5117
rect 44910 5108 44916 5120
rect 44968 5108 44974 5160
rect 45002 5108 45008 5160
rect 45060 5148 45066 5160
rect 46753 5151 46811 5157
rect 46753 5148 46765 5151
rect 45060 5120 46765 5148
rect 45060 5108 45066 5120
rect 46753 5117 46765 5120
rect 46799 5117 46811 5151
rect 46753 5111 46811 5117
rect 32088 5052 33456 5080
rect 32088 5040 32094 5052
rect 33502 5040 33508 5092
rect 33560 5080 33566 5092
rect 33560 5052 33605 5080
rect 33560 5040 33566 5052
rect 35066 5040 35072 5092
rect 35124 5080 35130 5092
rect 38746 5080 38752 5092
rect 35124 5052 38752 5080
rect 35124 5040 35130 5052
rect 38746 5040 38752 5052
rect 38804 5040 38810 5092
rect 39390 5040 39396 5092
rect 39448 5080 39454 5092
rect 58253 5083 58311 5089
rect 58253 5080 58265 5083
rect 39448 5052 58265 5080
rect 39448 5040 39454 5052
rect 58253 5049 58265 5052
rect 58299 5049 58311 5083
rect 58253 5043 58311 5049
rect 15243 4984 18920 5012
rect 15243 4981 15255 4984
rect 15197 4975 15255 4981
rect 19058 4972 19064 5024
rect 19116 5012 19122 5024
rect 21358 5012 21364 5024
rect 19116 4984 21364 5012
rect 19116 4972 19122 4984
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 24026 4972 24032 5024
rect 24084 5012 24090 5024
rect 25866 5012 25872 5024
rect 24084 4984 25872 5012
rect 24084 4972 24090 4984
rect 25866 4972 25872 4984
rect 25924 5012 25930 5024
rect 26513 5015 26571 5021
rect 26513 5012 26525 5015
rect 25924 4984 26525 5012
rect 25924 4972 25930 4984
rect 26513 4981 26525 4984
rect 26559 4981 26571 5015
rect 26513 4975 26571 4981
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 30190 5012 30196 5024
rect 27580 4984 30196 5012
rect 27580 4972 27586 4984
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 30282 4972 30288 5024
rect 30340 5012 30346 5024
rect 30929 5015 30987 5021
rect 30929 5012 30941 5015
rect 30340 4984 30941 5012
rect 30340 4972 30346 4984
rect 30929 4981 30941 4984
rect 30975 4981 30987 5015
rect 32398 5012 32404 5024
rect 32359 4984 32404 5012
rect 30929 4975 30987 4981
rect 32398 4972 32404 4984
rect 32456 4972 32462 5024
rect 32674 5012 32680 5024
rect 32635 4984 32680 5012
rect 32674 4972 32680 4984
rect 32732 4972 32738 5024
rect 33229 5015 33287 5021
rect 33229 4981 33241 5015
rect 33275 5012 33287 5015
rect 34422 5012 34428 5024
rect 33275 4984 34428 5012
rect 33275 4981 33287 4984
rect 33229 4975 33287 4981
rect 34422 4972 34428 4984
rect 34480 4972 34486 5024
rect 34790 4972 34796 5024
rect 34848 5012 34854 5024
rect 36538 5012 36544 5024
rect 34848 4984 36544 5012
rect 34848 4972 34854 4984
rect 36538 4972 36544 4984
rect 36596 4972 36602 5024
rect 36630 4972 36636 5024
rect 36688 5012 36694 5024
rect 37645 5015 37703 5021
rect 37645 5012 37657 5015
rect 36688 4984 37657 5012
rect 36688 4972 36694 4984
rect 37645 4981 37657 4984
rect 37691 4981 37703 5015
rect 37645 4975 37703 4981
rect 38470 4972 38476 5024
rect 38528 5012 38534 5024
rect 39117 5015 39175 5021
rect 39117 5012 39129 5015
rect 38528 4984 39129 5012
rect 38528 4972 38534 4984
rect 39117 4981 39129 4984
rect 39163 4981 39175 5015
rect 39117 4975 39175 4981
rect 39206 4972 39212 5024
rect 39264 5012 39270 5024
rect 40586 5012 40592 5024
rect 39264 4984 40592 5012
rect 39264 4972 39270 4984
rect 40586 4972 40592 4984
rect 40644 4972 40650 5024
rect 42702 4972 42708 5024
rect 42760 5012 42766 5024
rect 42797 5015 42855 5021
rect 42797 5012 42809 5015
rect 42760 4984 42809 5012
rect 42760 4972 42766 4984
rect 42797 4981 42809 4984
rect 42843 4981 42855 5015
rect 42797 4975 42855 4981
rect 43990 4972 43996 5024
rect 44048 5012 44054 5024
rect 45741 5015 45799 5021
rect 45741 5012 45753 5015
rect 44048 4984 45753 5012
rect 44048 4972 44054 4984
rect 45741 4981 45753 4984
rect 45787 4981 45799 5015
rect 45741 4975 45799 4981
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 9214 4808 9220 4820
rect 9175 4780 9220 4808
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 9398 4768 9404 4820
rect 9456 4768 9462 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9640 4780 10088 4808
rect 9640 4768 9646 4780
rect 7006 4740 7012 4752
rect 6967 4712 7012 4740
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 8573 4743 8631 4749
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 8662 4740 8668 4752
rect 8619 4712 8668 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 9416 4613 9444 4768
rect 10060 4740 10088 4780
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10192 4780 10701 4808
rect 10192 4768 10198 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 13633 4811 13691 4817
rect 12400 4780 13584 4808
rect 12400 4768 12406 4780
rect 10505 4743 10563 4749
rect 10505 4740 10517 4743
rect 10060 4712 10517 4740
rect 10505 4709 10517 4712
rect 10551 4709 10563 4743
rect 11698 4740 11704 4752
rect 11659 4712 11704 4740
rect 10505 4703 10563 4709
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 11793 4743 11851 4749
rect 11793 4709 11805 4743
rect 11839 4740 11851 4743
rect 12066 4740 12072 4752
rect 11839 4712 12072 4740
rect 11839 4709 11851 4712
rect 11793 4703 11851 4709
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 12526 4740 12532 4752
rect 12487 4712 12532 4740
rect 12526 4700 12532 4712
rect 12584 4700 12590 4752
rect 12894 4700 12900 4752
rect 12952 4740 12958 4752
rect 13449 4743 13507 4749
rect 13449 4740 13461 4743
rect 12952 4712 13461 4740
rect 12952 4700 12958 4712
rect 13449 4709 13461 4712
rect 13495 4709 13507 4743
rect 13556 4740 13584 4780
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13679 4780 19380 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 15013 4743 15071 4749
rect 15013 4740 15025 4743
rect 13556 4712 15025 4740
rect 13449 4703 13507 4709
rect 15013 4709 15025 4712
rect 15059 4709 15071 4743
rect 15013 4703 15071 4709
rect 15197 4743 15255 4749
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 19352 4740 19380 4780
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 26513 4811 26571 4817
rect 26513 4808 26525 4811
rect 19484 4780 26525 4808
rect 19484 4768 19490 4780
rect 26513 4777 26525 4780
rect 26559 4777 26571 4811
rect 26513 4771 26571 4777
rect 28074 4768 28080 4820
rect 28132 4808 28138 4820
rect 28537 4811 28595 4817
rect 28537 4808 28549 4811
rect 28132 4780 28549 4808
rect 28132 4768 28138 4780
rect 28537 4777 28549 4780
rect 28583 4808 28595 4811
rect 29822 4808 29828 4820
rect 28583 4780 28672 4808
rect 29783 4780 29828 4808
rect 28583 4777 28595 4780
rect 28537 4771 28595 4777
rect 28644 4752 28672 4780
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 30650 4768 30656 4820
rect 30708 4808 30714 4820
rect 32401 4811 32459 4817
rect 32401 4808 32413 4811
rect 30708 4780 32413 4808
rect 30708 4768 30714 4780
rect 32401 4777 32413 4780
rect 32447 4808 32459 4811
rect 33778 4808 33784 4820
rect 32447 4780 33784 4808
rect 32447 4777 32459 4780
rect 32401 4771 32459 4777
rect 33778 4768 33784 4780
rect 33836 4768 33842 4820
rect 34977 4811 35035 4817
rect 34977 4777 34989 4811
rect 35023 4808 35035 4811
rect 37090 4808 37096 4820
rect 35023 4780 37096 4808
rect 35023 4777 35035 4780
rect 34977 4771 35035 4777
rect 37090 4768 37096 4780
rect 37148 4768 37154 4820
rect 37829 4811 37887 4817
rect 37829 4777 37841 4811
rect 37875 4808 37887 4811
rect 37918 4808 37924 4820
rect 37875 4780 37924 4808
rect 37875 4777 37887 4780
rect 37829 4771 37887 4777
rect 37918 4768 37924 4780
rect 37976 4768 37982 4820
rect 40218 4768 40224 4820
rect 40276 4808 40282 4820
rect 40957 4811 41015 4817
rect 40957 4808 40969 4811
rect 40276 4780 40969 4808
rect 40276 4768 40282 4780
rect 40957 4777 40969 4780
rect 41003 4777 41015 4811
rect 42981 4811 43039 4817
rect 42981 4808 42993 4811
rect 40957 4771 41015 4777
rect 41386 4780 42993 4808
rect 20990 4740 20996 4752
rect 15243 4712 19288 4740
rect 19352 4712 20996 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 9640 4644 9685 4672
rect 9640 4632 9646 4644
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 9824 4644 10241 4672
rect 9824 4632 9830 4644
rect 10229 4641 10241 4644
rect 10275 4672 10287 4675
rect 10318 4672 10324 4684
rect 10275 4644 10324 4672
rect 10275 4641 10287 4644
rect 10229 4635 10287 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11330 4632 11336 4644
rect 11388 4672 11394 4684
rect 12158 4672 12164 4684
rect 11388 4644 12164 4672
rect 11388 4632 11394 4644
rect 12158 4632 12164 4644
rect 12216 4672 12222 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 12216 4644 12265 4672
rect 12216 4632 12222 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 19058 4672 19064 4684
rect 12253 4635 12311 4641
rect 18340 4644 19064 4672
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9493 4567 9551 4573
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 6825 4539 6883 4545
rect 6825 4536 6837 4539
rect 6696 4508 6837 4536
rect 6696 4496 6702 4508
rect 6825 4505 6837 4508
rect 6871 4505 6883 4539
rect 6825 4499 6883 4505
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8018 4536 8024 4548
rect 7699 4508 8024 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8018 4496 8024 4508
rect 8076 4496 8082 4548
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 8662 4536 8668 4548
rect 8435 4508 8668 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 9306 4496 9312 4548
rect 9364 4536 9370 4548
rect 9508 4536 9536 4567
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 15654 4604 15660 4616
rect 15615 4576 15660 4604
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 16574 4604 16580 4616
rect 16535 4576 16580 4604
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 18340 4604 18368 4644
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 19260 4672 19288 4712
rect 20990 4700 20996 4712
rect 21048 4700 21054 4752
rect 22002 4700 22008 4752
rect 22060 4740 22066 4752
rect 22097 4743 22155 4749
rect 22097 4740 22109 4743
rect 22060 4712 22109 4740
rect 22060 4700 22066 4712
rect 22097 4709 22109 4712
rect 22143 4709 22155 4743
rect 23474 4740 23480 4752
rect 22097 4703 22155 4709
rect 22204 4712 23480 4740
rect 21082 4672 21088 4684
rect 19260 4644 21088 4672
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 22204 4672 22232 4712
rect 23474 4700 23480 4712
rect 23532 4700 23538 4752
rect 28626 4700 28632 4752
rect 28684 4700 28690 4752
rect 36078 4700 36084 4752
rect 36136 4740 36142 4752
rect 38841 4743 38899 4749
rect 38841 4740 38853 4743
rect 36136 4712 38853 4740
rect 36136 4700 36142 4712
rect 38841 4709 38853 4712
rect 38887 4709 38899 4743
rect 38841 4703 38899 4709
rect 39298 4700 39304 4752
rect 39356 4740 39362 4752
rect 40313 4743 40371 4749
rect 40313 4740 40325 4743
rect 39356 4712 40325 4740
rect 39356 4700 39362 4712
rect 40313 4709 40325 4712
rect 40359 4709 40371 4743
rect 40313 4703 40371 4709
rect 40586 4700 40592 4752
rect 40644 4740 40650 4752
rect 41386 4740 41414 4780
rect 42981 4777 42993 4780
rect 43027 4777 43039 4811
rect 42981 4771 43039 4777
rect 44266 4768 44272 4820
rect 44324 4808 44330 4820
rect 45738 4808 45744 4820
rect 44324 4780 45744 4808
rect 44324 4768 44330 4780
rect 45738 4768 45744 4780
rect 45796 4768 45802 4820
rect 48222 4808 48228 4820
rect 45848 4780 48228 4808
rect 40644 4712 41414 4740
rect 40644 4700 40650 4712
rect 41506 4700 41512 4752
rect 41564 4740 41570 4752
rect 44085 4743 44143 4749
rect 44085 4740 44097 4743
rect 41564 4712 44097 4740
rect 41564 4700 41570 4712
rect 44085 4709 44097 4712
rect 44131 4709 44143 4743
rect 44085 4703 44143 4709
rect 44910 4700 44916 4752
rect 44968 4740 44974 4752
rect 45848 4740 45876 4780
rect 48222 4768 48228 4780
rect 48280 4768 48286 4820
rect 54202 4808 54208 4820
rect 54163 4780 54208 4808
rect 54202 4768 54208 4780
rect 54260 4768 54266 4820
rect 56686 4768 56692 4820
rect 56744 4808 56750 4820
rect 57333 4811 57391 4817
rect 57333 4808 57345 4811
rect 56744 4780 57345 4808
rect 56744 4768 56750 4780
rect 57333 4777 57345 4780
rect 57379 4777 57391 4811
rect 57333 4771 57391 4777
rect 44968 4712 45876 4740
rect 44968 4700 44974 4712
rect 21508 4644 22048 4672
rect 21508 4632 21514 4644
rect 17696 4576 18368 4604
rect 18417 4607 18475 4613
rect 9364 4508 9536 4536
rect 9364 4496 9370 4508
rect 12158 4496 12164 4548
rect 12216 4536 12222 4548
rect 13173 4539 13231 4545
rect 13173 4536 13185 4539
rect 12216 4508 13185 4536
rect 12216 4496 12222 4508
rect 13173 4505 13185 4508
rect 13219 4505 13231 4539
rect 13173 4499 13231 4505
rect 13538 4496 13544 4548
rect 13596 4536 13602 4548
rect 14737 4539 14795 4545
rect 14737 4536 14749 4539
rect 13596 4508 14749 4536
rect 13596 4496 13602 4508
rect 14737 4505 14749 4508
rect 14783 4536 14795 4539
rect 15838 4536 15844 4548
rect 14783 4508 15844 4536
rect 14783 4505 14795 4508
rect 14737 4499 14795 4505
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 15933 4539 15991 4545
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16758 4536 16764 4548
rect 15979 4508 16764 4536
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 16853 4539 16911 4545
rect 16853 4505 16865 4539
rect 16899 4536 16911 4539
rect 17218 4536 17224 4548
rect 16899 4508 17224 4536
rect 16899 4505 16911 4508
rect 16853 4499 16911 4505
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 9122 4468 9128 4480
rect 7791 4440 9128 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9490 4428 9496 4480
rect 9548 4468 9554 4480
rect 12342 4468 12348 4480
rect 9548 4440 12348 4468
rect 9548 4428 9554 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12713 4471 12771 4477
rect 12713 4437 12725 4471
rect 12759 4468 12771 4471
rect 17696 4468 17724 4576
rect 18417 4573 18429 4607
rect 18463 4604 18475 4607
rect 18506 4604 18512 4616
rect 18463 4576 18512 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19521 4607 19579 4613
rect 18616 4576 19334 4604
rect 17773 4539 17831 4545
rect 17773 4505 17785 4539
rect 17819 4536 17831 4539
rect 18616 4536 18644 4576
rect 17819 4508 18644 4536
rect 18693 4539 18751 4545
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 18693 4505 18705 4539
rect 18739 4505 18751 4539
rect 19306 4536 19334 4576
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 19610 4604 19616 4616
rect 19567 4576 19616 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 20714 4604 20720 4616
rect 19730 4576 20720 4604
rect 19730 4536 19758 4576
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 22020 4613 22048 4644
rect 22112 4644 22232 4672
rect 22112 4616 22140 4644
rect 22554 4632 22560 4684
rect 22612 4672 22618 4684
rect 22741 4675 22799 4681
rect 22741 4672 22753 4675
rect 22612 4644 22753 4672
rect 22612 4632 22618 4644
rect 22741 4641 22753 4644
rect 22787 4672 22799 4675
rect 23750 4672 23756 4684
rect 22787 4644 23756 4672
rect 22787 4641 22799 4644
rect 22741 4635 22799 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 23934 4672 23940 4684
rect 23895 4644 23940 4672
rect 23934 4632 23940 4644
rect 23992 4672 23998 4684
rect 24854 4672 24860 4684
rect 23992 4644 24860 4672
rect 23992 4632 23998 4644
rect 24854 4632 24860 4644
rect 24912 4632 24918 4684
rect 25130 4672 25136 4684
rect 25091 4644 25136 4672
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 27433 4675 27491 4681
rect 27433 4641 27445 4675
rect 27479 4641 27491 4675
rect 27433 4635 27491 4641
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20864 4576 20913 4604
rect 20864 4564 20870 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22244 4576 22293 4604
rect 22244 4564 22250 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 24762 4564 24768 4616
rect 24820 4604 24826 4616
rect 27341 4607 27399 4613
rect 27341 4604 27353 4607
rect 24820 4576 27353 4604
rect 24820 4564 24826 4576
rect 27341 4573 27353 4576
rect 27387 4573 27399 4607
rect 27448 4604 27476 4635
rect 27522 4632 27528 4684
rect 27580 4672 27586 4684
rect 27580 4644 27625 4672
rect 27580 4632 27586 4644
rect 28948 4632 28954 4684
rect 29006 4672 29012 4684
rect 30282 4672 30288 4684
rect 29006 4644 30288 4672
rect 29006 4632 29012 4644
rect 30282 4632 30288 4644
rect 30340 4632 30346 4684
rect 30466 4672 30472 4684
rect 30427 4644 30472 4672
rect 30466 4632 30472 4644
rect 30524 4632 30530 4684
rect 34606 4672 34612 4684
rect 32784 4644 34612 4672
rect 27982 4604 27988 4616
rect 27448 4576 27988 4604
rect 27341 4567 27399 4573
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 28350 4564 28356 4616
rect 28408 4604 28414 4616
rect 28445 4607 28503 4613
rect 28445 4604 28457 4607
rect 28408 4576 28457 4604
rect 28408 4564 28414 4576
rect 28445 4573 28457 4576
rect 28491 4573 28503 4607
rect 28445 4567 28503 4573
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 29178 4604 29184 4616
rect 28859 4576 29184 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 19306 4508 19758 4536
rect 19797 4539 19855 4545
rect 18693 4499 18751 4505
rect 19797 4505 19809 4539
rect 19843 4536 19855 4539
rect 20622 4536 20628 4548
rect 19843 4508 20628 4536
rect 19843 4505 19855 4508
rect 19797 4499 19855 4505
rect 12759 4440 17724 4468
rect 18708 4468 18736 4499
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 23661 4539 23719 4545
rect 23661 4505 23673 4539
rect 23707 4536 23719 4539
rect 24486 4536 24492 4548
rect 23707 4508 24492 4536
rect 23707 4505 23719 4508
rect 23661 4499 23719 4505
rect 24486 4496 24492 4508
rect 24544 4496 24550 4548
rect 24578 4496 24584 4548
rect 24636 4536 24642 4548
rect 25378 4539 25436 4545
rect 25378 4536 25390 4539
rect 24636 4508 25390 4536
rect 24636 4496 24642 4508
rect 25378 4505 25390 4508
rect 25424 4505 25436 4539
rect 27798 4536 27804 4548
rect 25378 4499 25436 4505
rect 26804 4508 27804 4536
rect 22646 4468 22652 4480
rect 18708 4440 22652 4468
rect 12759 4437 12771 4440
rect 12713 4431 12771 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 23566 4468 23572 4480
rect 23339 4440 23572 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4468 23811 4471
rect 26804 4468 26832 4508
rect 27798 4496 27804 4508
rect 27856 4496 27862 4548
rect 28460 4536 28488 4567
rect 29178 4564 29184 4576
rect 29236 4564 29242 4616
rect 30098 4564 30104 4616
rect 30156 4604 30162 4616
rect 30193 4607 30251 4613
rect 30193 4604 30205 4607
rect 30156 4576 30205 4604
rect 30156 4564 30162 4576
rect 30193 4573 30205 4576
rect 30239 4573 30251 4607
rect 30193 4567 30251 4573
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4604 31079 4607
rect 32306 4604 32312 4616
rect 31067 4576 32312 4604
rect 31067 4573 31079 4576
rect 31021 4567 31079 4573
rect 32306 4564 32312 4576
rect 32364 4564 32370 4616
rect 30834 4536 30840 4548
rect 28460 4508 30840 4536
rect 30834 4496 30840 4508
rect 30892 4496 30898 4548
rect 31288 4539 31346 4545
rect 31288 4505 31300 4539
rect 31334 4536 31346 4539
rect 32784 4536 32812 4644
rect 34606 4632 34612 4644
rect 34664 4632 34670 4684
rect 35526 4672 35532 4684
rect 35487 4644 35532 4672
rect 35526 4632 35532 4644
rect 35584 4632 35590 4684
rect 38286 4672 38292 4684
rect 36004 4644 38292 4672
rect 33594 4604 33600 4616
rect 33555 4576 33600 4604
rect 33594 4564 33600 4576
rect 33652 4564 33658 4616
rect 34057 4607 34115 4613
rect 34057 4573 34069 4607
rect 34103 4604 34115 4607
rect 36004 4604 36032 4644
rect 38286 4632 38292 4644
rect 38344 4632 38350 4684
rect 39942 4672 39948 4684
rect 38396 4644 39948 4672
rect 36170 4604 36176 4616
rect 34103 4576 36032 4604
rect 36131 4576 36176 4604
rect 34103 4573 34115 4576
rect 34057 4567 34115 4573
rect 32950 4536 32956 4548
rect 31334 4508 32812 4536
rect 32911 4508 32956 4536
rect 31334 4505 31346 4508
rect 31288 4499 31346 4505
rect 32950 4496 32956 4508
rect 33008 4496 33014 4548
rect 33134 4536 33140 4548
rect 33095 4508 33140 4536
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 26970 4468 26976 4480
rect 23799 4440 26832 4468
rect 26931 4440 26976 4468
rect 23799 4437 23811 4440
rect 23753 4431 23811 4437
rect 26970 4428 26976 4440
rect 27028 4428 27034 4480
rect 28994 4428 29000 4480
rect 29052 4468 29058 4480
rect 29052 4440 29097 4468
rect 29052 4428 29058 4440
rect 29178 4428 29184 4480
rect 29236 4468 29242 4480
rect 34072 4468 34100 4567
rect 36170 4564 36176 4576
rect 36228 4564 36234 4616
rect 36538 4564 36544 4616
rect 36596 4604 36602 4616
rect 37185 4607 37243 4613
rect 37185 4604 37197 4607
rect 36596 4576 37197 4604
rect 36596 4564 36602 4576
rect 37185 4573 37197 4576
rect 37231 4573 37243 4607
rect 37185 4567 37243 4573
rect 34333 4539 34391 4545
rect 34333 4505 34345 4539
rect 34379 4536 34391 4539
rect 34422 4536 34428 4548
rect 34379 4508 34428 4536
rect 34379 4505 34391 4508
rect 34333 4499 34391 4505
rect 34422 4496 34428 4508
rect 34480 4496 34486 4548
rect 36449 4539 36507 4545
rect 36449 4536 36461 4539
rect 35360 4508 36461 4536
rect 29236 4440 34100 4468
rect 29236 4428 29242 4440
rect 34238 4428 34244 4480
rect 34296 4468 34302 4480
rect 35360 4477 35388 4508
rect 36449 4505 36461 4508
rect 36495 4536 36507 4539
rect 36998 4536 37004 4548
rect 36495 4508 37004 4536
rect 36495 4505 36507 4508
rect 36449 4499 36507 4505
rect 36998 4496 37004 4508
rect 37056 4496 37062 4548
rect 37200 4536 37228 4567
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 37608 4576 38025 4604
rect 37608 4564 37614 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 38105 4607 38163 4613
rect 38105 4573 38117 4607
rect 38151 4604 38163 4607
rect 38396 4604 38424 4644
rect 39942 4632 39948 4644
rect 40000 4632 40006 4684
rect 40034 4632 40040 4684
rect 40092 4672 40098 4684
rect 43254 4672 43260 4684
rect 40092 4644 41414 4672
rect 40092 4632 40098 4644
rect 38151 4576 38424 4604
rect 38151 4573 38163 4576
rect 38105 4567 38163 4573
rect 38562 4564 38568 4616
rect 38620 4604 38626 4616
rect 40773 4607 40831 4613
rect 40773 4604 40785 4607
rect 38620 4576 40785 4604
rect 38620 4564 38626 4576
rect 40773 4573 40785 4576
rect 40819 4573 40831 4607
rect 41386 4604 41414 4644
rect 42500 4644 43260 4672
rect 41601 4607 41659 4613
rect 41601 4604 41613 4607
rect 41386 4576 41613 4604
rect 40773 4567 40831 4573
rect 41601 4573 41613 4576
rect 41647 4573 41659 4607
rect 42334 4604 42340 4616
rect 42295 4576 42340 4604
rect 41601 4567 41659 4573
rect 42334 4564 42340 4576
rect 42392 4564 42398 4616
rect 42500 4613 42528 4644
rect 43254 4632 43260 4644
rect 43312 4632 43318 4684
rect 43990 4672 43996 4684
rect 43824 4644 43996 4672
rect 42485 4607 42543 4613
rect 42485 4573 42497 4607
rect 42531 4573 42543 4607
rect 42485 4567 42543 4573
rect 42794 4564 42800 4616
rect 42852 4613 42858 4616
rect 42852 4604 42860 4613
rect 43530 4604 43536 4616
rect 42852 4576 42897 4604
rect 43491 4576 43536 4604
rect 42852 4567 42860 4576
rect 42852 4564 42858 4567
rect 43530 4564 43536 4576
rect 43588 4564 43594 4616
rect 43824 4613 43852 4644
rect 43990 4632 43996 4644
rect 44048 4632 44054 4684
rect 45462 4632 45468 4684
rect 45520 4672 45526 4684
rect 46109 4675 46167 4681
rect 46109 4672 46121 4675
rect 45520 4644 46121 4672
rect 45520 4632 45526 4644
rect 46109 4641 46121 4644
rect 46155 4641 46167 4675
rect 58158 4672 58164 4684
rect 58119 4644 58164 4672
rect 46109 4635 46167 4641
rect 58158 4632 58164 4644
rect 58216 4632 58222 4684
rect 43809 4607 43867 4613
rect 43809 4573 43821 4607
rect 43855 4573 43867 4607
rect 43809 4567 43867 4573
rect 43901 4607 43959 4613
rect 43901 4573 43913 4607
rect 43947 4573 43959 4607
rect 43901 4567 43959 4573
rect 37829 4539 37887 4545
rect 37829 4536 37841 4539
rect 37200 4508 37841 4536
rect 37829 4505 37841 4508
rect 37875 4505 37887 4539
rect 37829 4499 37887 4505
rect 35345 4471 35403 4477
rect 35345 4468 35357 4471
rect 34296 4440 35357 4468
rect 34296 4428 34302 4440
rect 35345 4437 35357 4440
rect 35391 4437 35403 4471
rect 35345 4431 35403 4437
rect 35437 4471 35495 4477
rect 35437 4437 35449 4471
rect 35483 4468 35495 4471
rect 35894 4468 35900 4480
rect 35483 4440 35900 4468
rect 35483 4437 35495 4440
rect 35437 4431 35495 4437
rect 35894 4428 35900 4440
rect 35952 4428 35958 4480
rect 35986 4428 35992 4480
rect 36044 4468 36050 4480
rect 37277 4471 37335 4477
rect 37277 4468 37289 4471
rect 36044 4440 37289 4468
rect 36044 4428 36050 4440
rect 37277 4437 37289 4440
rect 37323 4437 37335 4471
rect 37844 4468 37872 4499
rect 37918 4496 37924 4548
rect 37976 4536 37982 4548
rect 38657 4539 38715 4545
rect 38657 4536 38669 4539
rect 37976 4508 38669 4536
rect 37976 4496 37982 4508
rect 38657 4505 38669 4508
rect 38703 4505 38715 4539
rect 38657 4499 38715 4505
rect 38930 4496 38936 4548
rect 38988 4536 38994 4548
rect 40129 4539 40187 4545
rect 40129 4536 40141 4539
rect 38988 4508 40141 4536
rect 38988 4496 38994 4508
rect 40129 4505 40141 4508
rect 40175 4505 40187 4539
rect 40129 4499 40187 4505
rect 41322 4496 41328 4548
rect 41380 4536 41386 4548
rect 42613 4539 42671 4545
rect 42613 4536 42625 4539
rect 41380 4508 42625 4536
rect 41380 4496 41386 4508
rect 42613 4505 42625 4508
rect 42659 4505 42671 4539
rect 42613 4499 42671 4505
rect 42705 4539 42763 4545
rect 42705 4505 42717 4539
rect 42751 4536 42763 4539
rect 43162 4536 43168 4548
rect 42751 4508 43168 4536
rect 42751 4505 42763 4508
rect 42705 4499 42763 4505
rect 40862 4468 40868 4480
rect 37844 4440 40868 4468
rect 37277 4431 37335 4437
rect 40862 4428 40868 4440
rect 40920 4428 40926 4480
rect 41046 4428 41052 4480
rect 41104 4468 41110 4480
rect 41693 4471 41751 4477
rect 41693 4468 41705 4471
rect 41104 4440 41705 4468
rect 41104 4428 41110 4440
rect 41693 4437 41705 4440
rect 41739 4437 41751 4471
rect 42628 4468 42656 4499
rect 43162 4496 43168 4508
rect 43220 4496 43226 4548
rect 43714 4536 43720 4548
rect 43675 4508 43720 4536
rect 43714 4496 43720 4508
rect 43772 4496 43778 4548
rect 43916 4536 43944 4567
rect 45554 4564 45560 4616
rect 45612 4604 45618 4616
rect 51994 4604 52000 4616
rect 45612 4576 52000 4604
rect 45612 4564 45618 4576
rect 51994 4564 52000 4576
rect 52052 4564 52058 4616
rect 57330 4564 57336 4616
rect 57388 4604 57394 4616
rect 57885 4607 57943 4613
rect 57885 4604 57897 4607
rect 57388 4576 57897 4604
rect 57388 4564 57394 4576
rect 57885 4573 57897 4576
rect 57931 4573 57943 4607
rect 57885 4567 57943 4573
rect 45281 4539 45339 4545
rect 45281 4536 45293 4539
rect 43829 4508 43944 4536
rect 44192 4508 45293 4536
rect 43254 4468 43260 4480
rect 42628 4440 43260 4468
rect 41693 4431 41751 4437
rect 43254 4428 43260 4440
rect 43312 4468 43318 4480
rect 43829 4468 43857 4508
rect 43312 4440 43857 4468
rect 43312 4428 43318 4440
rect 43898 4428 43904 4480
rect 43956 4468 43962 4480
rect 44192 4468 44220 4508
rect 45281 4505 45293 4508
rect 45327 4505 45339 4539
rect 45281 4499 45339 4505
rect 45462 4496 45468 4548
rect 45520 4536 45526 4548
rect 46354 4539 46412 4545
rect 46354 4536 46366 4539
rect 45520 4508 46366 4536
rect 45520 4496 45526 4508
rect 46354 4505 46366 4508
rect 46400 4505 46412 4539
rect 46354 4499 46412 4505
rect 53926 4496 53932 4548
rect 53984 4536 53990 4548
rect 54113 4539 54171 4545
rect 54113 4536 54125 4539
rect 53984 4508 54125 4536
rect 53984 4496 53990 4508
rect 54113 4505 54125 4508
rect 54159 4505 54171 4539
rect 57238 4536 57244 4548
rect 57199 4508 57244 4536
rect 54113 4499 54171 4505
rect 57238 4496 57244 4508
rect 57296 4496 57302 4548
rect 43956 4440 44220 4468
rect 43956 4428 43962 4440
rect 44542 4428 44548 4480
rect 44600 4468 44606 4480
rect 45373 4471 45431 4477
rect 45373 4468 45385 4471
rect 44600 4440 45385 4468
rect 44600 4428 44606 4440
rect 45373 4437 45385 4440
rect 45419 4437 45431 4471
rect 45373 4431 45431 4437
rect 47489 4471 47547 4477
rect 47489 4437 47501 4471
rect 47535 4468 47547 4471
rect 48406 4468 48412 4480
rect 47535 4440 48412 4468
rect 47535 4437 47547 4440
rect 47489 4431 47547 4437
rect 48406 4428 48412 4440
rect 48464 4428 48470 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 5626 4264 5632 4276
rect 2884 4236 5632 4264
rect 2884 4205 2912 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 12894 4264 12900 4276
rect 7064 4236 12900 4264
rect 7064 4224 7070 4236
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4233 13323 4267
rect 13265 4227 13323 4233
rect 14108 4236 17080 4264
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4165 2927 4199
rect 2869 4159 2927 4165
rect 3605 4199 3663 4205
rect 3605 4165 3617 4199
rect 3651 4196 3663 4199
rect 4341 4199 4399 4205
rect 3651 4168 4292 4196
rect 3651 4165 3663 4168
rect 3605 4159 3663 4165
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 3142 4128 3148 4140
rect 1627 4100 3148 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3789 4131 3847 4137
rect 3789 4128 3801 4131
rect 3752 4100 3801 4128
rect 3752 4088 3758 4100
rect 3789 4097 3801 4100
rect 3835 4097 3847 4131
rect 4264 4128 4292 4168
rect 4341 4165 4353 4199
rect 4387 4196 4399 4199
rect 4614 4196 4620 4208
rect 4387 4168 4620 4196
rect 4387 4165 4399 4168
rect 4341 4159 4399 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 5813 4199 5871 4205
rect 4724 4168 5764 4196
rect 4724 4128 4752 4168
rect 4264 4100 4752 4128
rect 5736 4128 5764 4168
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6362 4196 6368 4208
rect 5859 4168 6368 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 7101 4199 7159 4205
rect 7101 4165 7113 4199
rect 7147 4196 7159 4199
rect 7742 4196 7748 4208
rect 7147 4168 7748 4196
rect 7147 4165 7159 4168
rect 7101 4159 7159 4165
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 8110 4196 8116 4208
rect 7984 4168 8116 4196
rect 7984 4156 7990 4168
rect 8110 4156 8116 4168
rect 8168 4196 8174 4208
rect 8168 4168 9076 4196
rect 8168 4156 8174 4168
rect 6914 4128 6920 4140
rect 5736 4100 6920 4128
rect 3789 4091 3847 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 8846 4128 8852 4140
rect 7668 4100 8156 4128
rect 8807 4100 8852 4128
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 7668 4060 7696 4100
rect 2924 4032 7696 4060
rect 7745 4063 7803 4069
rect 2924 4020 2930 4032
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 7926 4060 7932 4072
rect 7791 4032 7932 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 3053 3995 3111 4001
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 5350 3992 5356 4004
rect 3099 3964 5356 3992
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6454 3992 6460 4004
rect 6043 3964 6460 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 6604 3964 8033 3992
rect 6604 3952 6610 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 5534 3924 5540 3936
rect 4479 3896 5540 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8128 3924 8156 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9048 4137 9076 4168
rect 11974 4156 11980 4208
rect 12032 4196 12038 4208
rect 13280 4196 13308 4227
rect 13538 4196 13544 4208
rect 12032 4168 13308 4196
rect 13372 4168 13544 4196
rect 12032 4156 12038 4168
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9582 4128 9588 4140
rect 9079 4100 9588 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4128 10379 4131
rect 12158 4128 12164 4140
rect 10367 4100 12164 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 13173 4131 13231 4137
rect 12728 4100 13124 4128
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8444 4032 8677 4060
rect 8444 4020 8450 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9125 4063 9183 4069
rect 8996 4032 9041 4060
rect 8996 4020 9002 4032
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4060 12679 4063
rect 12728 4060 12756 4100
rect 12667 4032 12756 4060
rect 13096 4060 13124 4100
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13372 4128 13400 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 13998 4128 14004 4140
rect 13219 4100 13400 4128
rect 13959 4100 14004 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14108 4060 14136 4236
rect 15930 4156 15936 4208
rect 15988 4196 15994 4208
rect 16117 4199 16175 4205
rect 16117 4196 16129 4199
rect 15988 4168 16129 4196
rect 15988 4156 15994 4168
rect 16117 4165 16129 4168
rect 16163 4165 16175 4199
rect 16942 4196 16948 4208
rect 16903 4168 16948 4196
rect 16117 4159 16175 4165
rect 16942 4156 16948 4168
rect 17000 4156 17006 4208
rect 17052 4196 17080 4236
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 18322 4264 18328 4276
rect 17276 4236 18328 4264
rect 17276 4224 17282 4236
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19392 4236 19620 4264
rect 19392 4224 19398 4236
rect 19242 4196 19248 4208
rect 17052 4168 19248 4196
rect 19242 4156 19248 4168
rect 19300 4156 19306 4208
rect 19592 4196 19620 4236
rect 19702 4224 19708 4276
rect 19760 4264 19766 4276
rect 20346 4264 20352 4276
rect 19760 4236 19805 4264
rect 19996 4236 20352 4264
rect 19760 4224 19766 4236
rect 19996 4205 20024 4236
rect 20346 4224 20352 4236
rect 20404 4224 20410 4276
rect 20717 4267 20775 4273
rect 20717 4233 20729 4267
rect 20763 4233 20775 4267
rect 20717 4227 20775 4233
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 20898 4264 20904 4276
rect 20855 4236 20904 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 19815 4199 19873 4205
rect 19815 4196 19827 4199
rect 19592 4168 19827 4196
rect 19815 4165 19827 4168
rect 19861 4165 19873 4199
rect 19815 4159 19873 4165
rect 19981 4199 20039 4205
rect 19981 4165 19993 4199
rect 20027 4165 20039 4199
rect 19981 4159 20039 4165
rect 20438 4156 20444 4208
rect 20496 4196 20502 4208
rect 20732 4196 20760 4227
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 22094 4264 22100 4276
rect 21376 4236 22100 4264
rect 21376 4196 21404 4236
rect 22094 4224 22100 4236
rect 22152 4224 22158 4276
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 23301 4267 23359 4273
rect 23301 4264 23313 4267
rect 22244 4236 23313 4264
rect 22244 4224 22250 4236
rect 23301 4233 23313 4236
rect 23347 4233 23359 4267
rect 23301 4227 23359 4233
rect 23937 4267 23995 4273
rect 23937 4233 23949 4267
rect 23983 4264 23995 4267
rect 24394 4264 24400 4276
rect 23983 4236 24400 4264
rect 23983 4233 23995 4236
rect 23937 4227 23995 4233
rect 24394 4224 24400 4236
rect 24452 4224 24458 4276
rect 29178 4264 29184 4276
rect 24504 4236 29184 4264
rect 20496 4168 20541 4196
rect 20732 4168 21404 4196
rect 20496 4156 20502 4168
rect 21726 4156 21732 4208
rect 21784 4196 21790 4208
rect 22462 4196 22468 4208
rect 21784 4168 22468 4196
rect 21784 4156 21790 4168
rect 22462 4156 22468 4168
rect 22520 4156 22526 4208
rect 22925 4199 22983 4205
rect 22925 4196 22937 4199
rect 22572 4168 22937 4196
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15654 4088 15660 4140
rect 15712 4128 15718 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15712 4100 15853 4128
rect 15712 4088 15718 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 18506 4128 18512 4140
rect 18467 4100 18512 4128
rect 15841 4091 15899 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 20622 4128 20628 4140
rect 19668 4100 19713 4128
rect 20535 4100 20628 4128
rect 19668 4088 19674 4100
rect 20622 4088 20628 4100
rect 20680 4128 20686 4140
rect 20806 4128 20812 4140
rect 20680 4100 20812 4128
rect 20680 4088 20686 4100
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 20990 4128 20996 4140
rect 20951 4100 20996 4128
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 13096 4032 14136 4060
rect 14277 4063 14335 4069
rect 12667 4029 12679 4032
rect 12621 4023 12679 4029
rect 14277 4029 14289 4063
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 15197 4063 15255 4069
rect 15197 4029 15209 4063
rect 15243 4060 15255 4063
rect 15378 4060 15384 4072
rect 15243 4032 15384 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3992 8263 3995
rect 9140 3992 9168 4023
rect 8251 3964 9168 3992
rect 10689 3995 10747 4001
rect 8251 3961 8263 3964
rect 8205 3955 8263 3961
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 11054 3992 11060 4004
rect 10735 3964 11060 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3992 12587 3995
rect 12710 3992 12716 4004
rect 12575 3964 12716 3992
rect 12575 3961 12587 3964
rect 12529 3955 12587 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 14292 3992 14320 4023
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 17586 4060 17592 4072
rect 17547 4032 17592 4060
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 18230 4060 18236 4072
rect 17696 4032 18236 4060
rect 17696 3992 17724 4032
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18690 4060 18696 4072
rect 18651 4032 18696 4060
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19484 4032 19529 4060
rect 19484 4020 19490 4032
rect 14292 3964 17724 3992
rect 17865 3995 17923 4001
rect 17865 3961 17877 3995
rect 17911 3961 17923 3995
rect 17865 3955 17923 3961
rect 9398 3924 9404 3936
rect 8128 3896 9404 3924
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 10594 3924 10600 3936
rect 9907 3896 10600 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 10781 3927 10839 3933
rect 10781 3893 10793 3927
rect 10827 3924 10839 3927
rect 12434 3924 12440 3936
rect 10827 3896 12440 3924
rect 10827 3893 10839 3896
rect 10781 3887 10839 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 17880 3924 17908 3955
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 21634 3992 21640 4004
rect 21048 3964 21640 3992
rect 21048 3952 21054 3964
rect 21634 3952 21640 3964
rect 21692 3952 21698 4004
rect 22020 3992 22048 4091
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 22572 4128 22600 4168
rect 22925 4165 22937 4168
rect 22971 4165 22983 4199
rect 24302 4196 24308 4208
rect 24263 4168 24308 4196
rect 22925 4159 22983 4165
rect 24302 4156 24308 4168
rect 24360 4156 24366 4208
rect 22428 4100 22600 4128
rect 22428 4088 22434 4100
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23017 4131 23075 4137
rect 22796 4100 22841 4128
rect 22796 4088 22802 4100
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 23161 4131 23219 4137
rect 23161 4097 23173 4131
rect 23207 4128 23219 4131
rect 23290 4128 23296 4140
rect 23207 4100 23296 4128
rect 23207 4097 23219 4100
rect 23161 4091 23219 4097
rect 23032 4060 23060 4091
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 23382 4088 23388 4140
rect 23440 4128 23446 4140
rect 24504 4128 24532 4236
rect 29178 4224 29184 4236
rect 29236 4224 29242 4276
rect 29362 4224 29368 4276
rect 29420 4264 29426 4276
rect 29549 4267 29607 4273
rect 29549 4264 29561 4267
rect 29420 4236 29561 4264
rect 29420 4224 29426 4236
rect 29549 4233 29561 4236
rect 29595 4264 29607 4267
rect 31757 4267 31815 4273
rect 31757 4264 31769 4267
rect 29595 4236 31769 4264
rect 29595 4233 29607 4236
rect 29549 4227 29607 4233
rect 31757 4233 31769 4236
rect 31803 4233 31815 4267
rect 32306 4264 32312 4276
rect 32267 4236 32312 4264
rect 31757 4227 31815 4233
rect 32306 4224 32312 4236
rect 32364 4224 32370 4276
rect 32582 4224 32588 4276
rect 32640 4264 32646 4276
rect 32677 4267 32735 4273
rect 32677 4264 32689 4267
rect 32640 4236 32689 4264
rect 32640 4224 32646 4236
rect 32677 4233 32689 4236
rect 32723 4233 32735 4267
rect 32677 4227 32735 4233
rect 35621 4267 35679 4273
rect 35621 4233 35633 4267
rect 35667 4264 35679 4267
rect 35894 4264 35900 4276
rect 35667 4236 35900 4264
rect 35667 4233 35679 4236
rect 35621 4227 35679 4233
rect 35894 4224 35900 4236
rect 35952 4264 35958 4276
rect 36722 4264 36728 4276
rect 35952 4236 36728 4264
rect 35952 4224 35958 4236
rect 36722 4224 36728 4236
rect 36780 4264 36786 4276
rect 39390 4264 39396 4276
rect 36780 4236 39396 4264
rect 36780 4224 36786 4236
rect 39390 4224 39396 4236
rect 39448 4224 39454 4276
rect 39485 4267 39543 4273
rect 39485 4233 39497 4267
rect 39531 4233 39543 4267
rect 45922 4264 45928 4276
rect 45883 4236 45928 4264
rect 39485 4227 39543 4233
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 27430 4196 27436 4208
rect 24912 4168 27436 4196
rect 24912 4156 24918 4168
rect 27430 4156 27436 4168
rect 27488 4156 27494 4208
rect 27525 4199 27583 4205
rect 27525 4165 27537 4199
rect 27571 4196 27583 4199
rect 27614 4196 27620 4208
rect 27571 4168 27620 4196
rect 27571 4165 27583 4168
rect 27525 4159 27583 4165
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 28718 4156 28724 4208
rect 28776 4196 28782 4208
rect 28902 4196 28908 4208
rect 28776 4168 28908 4196
rect 28776 4156 28782 4168
rect 28902 4156 28908 4168
rect 28960 4156 28966 4208
rect 28994 4156 29000 4208
rect 29052 4196 29058 4208
rect 35710 4196 35716 4208
rect 29052 4168 35716 4196
rect 29052 4156 29058 4168
rect 35710 4156 35716 4168
rect 35768 4156 35774 4208
rect 37458 4156 37464 4208
rect 37516 4196 37522 4208
rect 37553 4199 37611 4205
rect 37553 4196 37565 4199
rect 37516 4168 37565 4196
rect 37516 4156 37522 4168
rect 37553 4165 37565 4168
rect 37599 4165 37611 4199
rect 38654 4196 38660 4208
rect 38615 4168 38660 4196
rect 37553 4159 37611 4165
rect 38654 4156 38660 4168
rect 38712 4196 38718 4208
rect 39500 4196 39528 4227
rect 45922 4224 45928 4236
rect 45980 4224 45986 4276
rect 53466 4224 53472 4276
rect 53524 4264 53530 4276
rect 54573 4267 54631 4273
rect 54573 4264 54585 4267
rect 53524 4236 54585 4264
rect 53524 4224 53530 4236
rect 54573 4233 54585 4236
rect 54619 4233 54631 4267
rect 54573 4227 54631 4233
rect 40129 4199 40187 4205
rect 40129 4196 40141 4199
rect 38712 4168 40141 4196
rect 38712 4156 38718 4168
rect 40129 4165 40141 4168
rect 40175 4196 40187 4199
rect 41601 4199 41659 4205
rect 41601 4196 41613 4199
rect 40175 4168 41613 4196
rect 40175 4165 40187 4168
rect 40129 4159 40187 4165
rect 41601 4165 41613 4168
rect 41647 4165 41659 4199
rect 41601 4159 41659 4165
rect 42242 4156 42248 4208
rect 42300 4196 42306 4208
rect 42300 4168 44036 4196
rect 42300 4156 42306 4168
rect 25130 4128 25136 4140
rect 23440 4100 24532 4128
rect 25091 4100 25136 4128
rect 23440 4088 23446 4100
rect 25130 4088 25136 4100
rect 25188 4088 25194 4140
rect 25406 4137 25412 4140
rect 25400 4091 25412 4137
rect 25464 4128 25470 4140
rect 25464 4100 25500 4128
rect 25406 4088 25412 4091
rect 25464 4088 25470 4100
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 27246 4128 27252 4140
rect 25832 4100 27252 4128
rect 25832 4088 25838 4100
rect 27246 4088 27252 4100
rect 27304 4088 27310 4140
rect 28537 4131 28595 4137
rect 28537 4128 28549 4131
rect 28460 4100 28549 4128
rect 24210 4060 24216 4072
rect 23032 4032 24216 4060
rect 24210 4020 24216 4032
rect 24268 4020 24274 4072
rect 24397 4063 24455 4069
rect 24397 4029 24409 4063
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4060 24639 4063
rect 24854 4060 24860 4072
rect 24627 4032 24860 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 24412 3992 24440 4023
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 27614 4060 27620 4072
rect 27575 4032 27620 4060
rect 27614 4020 27620 4032
rect 27672 4020 27678 4072
rect 27709 4063 27767 4069
rect 27709 4029 27721 4063
rect 27755 4060 27767 4063
rect 27890 4060 27896 4072
rect 27755 4032 27896 4060
rect 27755 4029 27767 4032
rect 27709 4023 27767 4029
rect 27890 4020 27896 4032
rect 27948 4020 27954 4072
rect 28350 4060 28356 4072
rect 28311 4032 28356 4060
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 25038 3992 25044 4004
rect 22020 3964 24348 3992
rect 24412 3964 25044 3992
rect 13044 3896 17908 3924
rect 18049 3927 18107 3933
rect 13044 3884 13050 3896
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 19978 3924 19984 3936
rect 18095 3896 19984 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 21876 3896 22201 3924
rect 21876 3884 21882 3896
rect 22189 3893 22201 3896
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 23198 3924 23204 3936
rect 22888 3896 23204 3924
rect 22888 3884 22894 3896
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 24320 3924 24348 3964
rect 25038 3952 25044 3964
rect 25096 3952 25102 4004
rect 28460 3992 28488 4100
rect 28537 4097 28549 4100
rect 28583 4097 28595 4131
rect 30633 4131 30691 4137
rect 30633 4128 30645 4131
rect 28537 4091 28595 4097
rect 28966 4100 30645 4128
rect 28626 4020 28632 4072
rect 28684 4060 28690 4072
rect 28966 4060 28994 4100
rect 30633 4097 30645 4100
rect 30679 4097 30691 4131
rect 30633 4091 30691 4097
rect 32769 4131 32827 4137
rect 32769 4097 32781 4131
rect 32815 4128 32827 4131
rect 33226 4128 33232 4140
rect 32815 4100 33232 4128
rect 32815 4097 32827 4100
rect 32769 4091 32827 4097
rect 33226 4088 33232 4100
rect 33284 4088 33290 4140
rect 33502 4088 33508 4140
rect 33560 4128 33566 4140
rect 33597 4131 33655 4137
rect 33597 4128 33609 4131
rect 33560 4100 33609 4128
rect 33560 4088 33566 4100
rect 33597 4097 33609 4100
rect 33643 4097 33655 4131
rect 33597 4091 33655 4097
rect 33686 4088 33692 4140
rect 33744 4128 33750 4140
rect 35342 4128 35348 4140
rect 33744 4100 35348 4128
rect 33744 4088 33750 4100
rect 35342 4088 35348 4100
rect 35400 4088 35406 4140
rect 36262 4128 36268 4140
rect 35728 4100 36268 4128
rect 28684 4032 28994 4060
rect 28684 4020 28690 4032
rect 29454 4020 29460 4072
rect 29512 4060 29518 4072
rect 29641 4063 29699 4069
rect 29641 4060 29653 4063
rect 29512 4032 29653 4060
rect 29512 4020 29518 4032
rect 29641 4029 29653 4032
rect 29687 4029 29699 4063
rect 29641 4023 29699 4029
rect 29730 4020 29736 4072
rect 29788 4060 29794 4072
rect 29788 4032 29833 4060
rect 29788 4020 29794 4032
rect 29914 4020 29920 4072
rect 29972 4060 29978 4072
rect 35728 4069 35756 4100
rect 36262 4088 36268 4100
rect 36320 4088 36326 4140
rect 36446 4128 36452 4140
rect 36407 4100 36452 4128
rect 36446 4088 36452 4100
rect 36504 4088 36510 4140
rect 36998 4088 37004 4140
rect 37056 4128 37062 4140
rect 38930 4128 38936 4140
rect 37056 4100 38936 4128
rect 37056 4088 37062 4100
rect 38930 4088 38936 4100
rect 38988 4088 38994 4140
rect 39298 4128 39304 4140
rect 39259 4100 39304 4128
rect 39298 4088 39304 4100
rect 39356 4088 39362 4140
rect 39942 4088 39948 4140
rect 40000 4128 40006 4140
rect 40865 4131 40923 4137
rect 40865 4128 40877 4131
rect 40000 4100 40877 4128
rect 40000 4088 40006 4100
rect 40865 4097 40877 4100
rect 40911 4097 40923 4131
rect 40865 4091 40923 4097
rect 42518 4088 42524 4140
rect 42576 4128 42582 4140
rect 42613 4131 42671 4137
rect 42613 4128 42625 4131
rect 42576 4100 42625 4128
rect 42576 4088 42582 4100
rect 42613 4097 42625 4100
rect 42659 4097 42671 4131
rect 43254 4128 43260 4140
rect 43215 4100 43260 4128
rect 42613 4091 42671 4097
rect 43254 4088 43260 4100
rect 43312 4088 43318 4140
rect 43625 4131 43683 4137
rect 43625 4097 43637 4131
rect 43671 4128 43683 4131
rect 43714 4128 43720 4140
rect 43671 4100 43720 4128
rect 43671 4097 43683 4100
rect 43625 4091 43683 4097
rect 43714 4088 43720 4100
rect 43772 4088 43778 4140
rect 44008 4128 44036 4168
rect 45094 4156 45100 4208
rect 45152 4196 45158 4208
rect 45152 4168 45197 4196
rect 45152 4156 45158 4168
rect 45738 4156 45744 4208
rect 45796 4196 45802 4208
rect 45833 4199 45891 4205
rect 45833 4196 45845 4199
rect 45796 4168 45845 4196
rect 45796 4156 45802 4168
rect 45833 4165 45845 4168
rect 45879 4165 45891 4199
rect 45833 4159 45891 4165
rect 48866 4156 48872 4208
rect 48924 4196 48930 4208
rect 49145 4199 49203 4205
rect 49145 4196 49157 4199
rect 48924 4168 49157 4196
rect 48924 4156 48930 4168
rect 49145 4165 49157 4168
rect 49191 4165 49203 4199
rect 49145 4159 49203 4165
rect 50614 4156 50620 4208
rect 50672 4196 50678 4208
rect 50709 4199 50767 4205
rect 50709 4196 50721 4199
rect 50672 4168 50721 4196
rect 50672 4156 50678 4168
rect 50709 4165 50721 4168
rect 50755 4165 50767 4199
rect 50709 4159 50767 4165
rect 51350 4156 51356 4208
rect 51408 4196 51414 4208
rect 51537 4199 51595 4205
rect 51537 4196 51549 4199
rect 51408 4168 51549 4196
rect 51408 4156 51414 4168
rect 51537 4165 51549 4168
rect 51583 4165 51595 4199
rect 51537 4159 51595 4165
rect 52454 4156 52460 4208
rect 52512 4196 52518 4208
rect 53009 4199 53067 4205
rect 53009 4196 53021 4199
rect 52512 4168 53021 4196
rect 52512 4156 52518 4168
rect 53009 4165 53021 4168
rect 53055 4165 53067 4199
rect 53009 4159 53067 4165
rect 53098 4156 53104 4208
rect 53156 4196 53162 4208
rect 53745 4199 53803 4205
rect 53745 4196 53757 4199
rect 53156 4168 53757 4196
rect 53156 4156 53162 4168
rect 53745 4165 53757 4168
rect 53791 4165 53803 4199
rect 53745 4159 53803 4165
rect 57882 4156 57888 4208
rect 57940 4196 57946 4208
rect 58161 4199 58219 4205
rect 58161 4196 58173 4199
rect 57940 4168 58173 4196
rect 57940 4156 57946 4168
rect 58161 4165 58173 4168
rect 58207 4165 58219 4199
rect 58161 4159 58219 4165
rect 44361 4131 44419 4137
rect 44008 4126 44312 4128
rect 44361 4126 44373 4131
rect 44008 4100 44373 4126
rect 44284 4098 44373 4100
rect 44361 4097 44373 4098
rect 44407 4097 44419 4131
rect 44361 4091 44419 4097
rect 44542 4088 44548 4140
rect 44600 4128 44606 4140
rect 46569 4131 46627 4137
rect 46569 4128 46581 4131
rect 44600 4126 45048 4128
rect 45204 4126 46581 4128
rect 44600 4100 46581 4126
rect 44600 4088 44606 4100
rect 45020 4098 45232 4100
rect 46569 4097 46581 4100
rect 46615 4097 46627 4131
rect 46750 4128 46756 4140
rect 46711 4100 46756 4128
rect 46569 4091 46627 4097
rect 46750 4088 46756 4100
rect 46808 4088 46814 4140
rect 48222 4128 48228 4140
rect 48183 4100 48228 4128
rect 48222 4088 48228 4100
rect 48280 4088 48286 4140
rect 48406 4128 48412 4140
rect 48367 4100 48412 4128
rect 48406 4088 48412 4100
rect 48464 4088 48470 4140
rect 49234 4088 49240 4140
rect 49292 4128 49298 4140
rect 49329 4131 49387 4137
rect 49329 4128 49341 4131
rect 49292 4100 49341 4128
rect 49292 4088 49298 4100
rect 49329 4097 49341 4100
rect 49375 4097 49387 4131
rect 49329 4091 49387 4097
rect 50798 4088 50804 4140
rect 50856 4128 50862 4140
rect 50893 4131 50951 4137
rect 50893 4128 50905 4131
rect 50856 4100 50905 4128
rect 50856 4088 50862 4100
rect 50893 4097 50905 4100
rect 50939 4097 50951 4131
rect 51718 4128 51724 4140
rect 51679 4100 51724 4128
rect 50893 4091 50951 4097
rect 51718 4088 51724 4100
rect 51776 4088 51782 4140
rect 53190 4128 53196 4140
rect 53151 4100 53196 4128
rect 53190 4088 53196 4100
rect 53248 4088 53254 4140
rect 53282 4088 53288 4140
rect 53340 4128 53346 4140
rect 53929 4131 53987 4137
rect 53929 4128 53941 4131
rect 53340 4100 53941 4128
rect 53340 4088 53346 4100
rect 53929 4097 53941 4100
rect 53975 4097 53987 4131
rect 53929 4091 53987 4097
rect 54110 4088 54116 4140
rect 54168 4128 54174 4140
rect 54389 4131 54447 4137
rect 54389 4128 54401 4131
rect 54168 4100 54401 4128
rect 54168 4088 54174 4100
rect 54389 4097 54401 4100
rect 54435 4097 54447 4131
rect 54389 4091 54447 4097
rect 55125 4131 55183 4137
rect 55125 4097 55137 4131
rect 55171 4097 55183 4131
rect 55125 4091 55183 4097
rect 57241 4131 57299 4137
rect 57241 4097 57253 4131
rect 57287 4128 57299 4131
rect 57974 4128 57980 4140
rect 57287 4100 57980 4128
rect 57287 4097 57299 4100
rect 57241 4091 57299 4097
rect 30377 4063 30435 4069
rect 30377 4060 30389 4063
rect 29972 4032 30389 4060
rect 29972 4020 29978 4032
rect 30377 4029 30389 4032
rect 30423 4029 30435 4063
rect 30377 4023 30435 4029
rect 32861 4063 32919 4069
rect 32861 4029 32873 4063
rect 32907 4060 32919 4063
rect 33873 4063 33931 4069
rect 33873 4060 33885 4063
rect 32907 4032 33885 4060
rect 32907 4029 32919 4032
rect 32861 4023 32919 4029
rect 33873 4029 33885 4032
rect 33919 4029 33931 4063
rect 35713 4063 35771 4069
rect 35713 4060 35725 4063
rect 33873 4023 33931 4029
rect 34624 4032 35725 4060
rect 29748 3992 29776 4020
rect 28460 3964 29776 3992
rect 31754 3952 31760 4004
rect 31812 3992 31818 4004
rect 32876 3992 32904 4023
rect 31812 3964 32904 3992
rect 31812 3952 31818 3964
rect 26513 3927 26571 3933
rect 26513 3924 26525 3927
rect 24320 3896 26525 3924
rect 26513 3893 26525 3896
rect 26559 3893 26571 3927
rect 27154 3924 27160 3936
rect 27115 3896 27160 3924
rect 26513 3887 26571 3893
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 27338 3884 27344 3936
rect 27396 3924 27402 3936
rect 28442 3924 28448 3936
rect 27396 3896 28448 3924
rect 27396 3884 27402 3896
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 28534 3884 28540 3936
rect 28592 3924 28598 3936
rect 28721 3927 28779 3933
rect 28721 3924 28733 3927
rect 28592 3896 28733 3924
rect 28592 3884 28598 3896
rect 28721 3893 28733 3896
rect 28767 3893 28779 3927
rect 29178 3924 29184 3936
rect 29139 3896 29184 3924
rect 28721 3887 28779 3893
rect 29178 3884 29184 3896
rect 29236 3884 29242 3936
rect 29914 3884 29920 3936
rect 29972 3924 29978 3936
rect 34624 3924 34652 4032
rect 35713 4029 35725 4032
rect 35759 4029 35771 4063
rect 35713 4023 35771 4029
rect 35805 4063 35863 4069
rect 35805 4029 35817 4063
rect 35851 4060 35863 4063
rect 35894 4060 35900 4072
rect 35851 4032 35900 4060
rect 35851 4029 35863 4032
rect 35805 4023 35863 4029
rect 35894 4020 35900 4032
rect 35952 4060 35958 4072
rect 36354 4060 36360 4072
rect 35952 4032 36360 4060
rect 35952 4020 35958 4032
rect 36354 4020 36360 4032
rect 36412 4020 36418 4072
rect 36633 4063 36691 4069
rect 36633 4029 36645 4063
rect 36679 4029 36691 4063
rect 36633 4023 36691 4029
rect 34790 3952 34796 4004
rect 34848 3992 34854 4004
rect 36648 3992 36676 4023
rect 38746 4020 38752 4072
rect 38804 4060 38810 4072
rect 40313 4063 40371 4069
rect 40313 4060 40325 4063
rect 38804 4032 40325 4060
rect 38804 4020 38810 4032
rect 40313 4029 40325 4032
rect 40359 4029 40371 4063
rect 40313 4023 40371 4029
rect 40402 4020 40408 4072
rect 40460 4060 40466 4072
rect 41049 4063 41107 4069
rect 41049 4060 41061 4063
rect 40460 4032 41061 4060
rect 40460 4020 40466 4032
rect 41049 4029 41061 4032
rect 41095 4029 41107 4063
rect 41049 4023 41107 4029
rect 41506 4020 41512 4072
rect 41564 4060 41570 4072
rect 42978 4060 42984 4072
rect 41564 4032 42984 4060
rect 41564 4020 41570 4032
rect 42978 4020 42984 4032
rect 43036 4020 43042 4072
rect 43349 4063 43407 4069
rect 43349 4029 43361 4063
rect 43395 4029 43407 4063
rect 43530 4060 43536 4072
rect 43491 4032 43536 4060
rect 43349 4023 43407 4029
rect 37918 3992 37924 4004
rect 34848 3964 36676 3992
rect 36740 3964 37924 3992
rect 34848 3952 34854 3964
rect 29972 3896 34652 3924
rect 35253 3927 35311 3933
rect 29972 3884 29978 3896
rect 35253 3893 35265 3927
rect 35299 3924 35311 3927
rect 35342 3924 35348 3936
rect 35299 3896 35348 3924
rect 35299 3893 35311 3896
rect 35253 3887 35311 3893
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 35618 3884 35624 3936
rect 35676 3924 35682 3936
rect 36740 3924 36768 3964
rect 37918 3952 37924 3964
rect 37976 3952 37982 4004
rect 39114 3992 39120 4004
rect 38028 3964 39120 3992
rect 37642 3924 37648 3936
rect 35676 3896 36768 3924
rect 37603 3896 37648 3924
rect 35676 3884 35682 3896
rect 37642 3884 37648 3896
rect 37700 3884 37706 3936
rect 37734 3884 37740 3936
rect 37792 3924 37798 3936
rect 38028 3924 38056 3964
rect 39114 3952 39120 3964
rect 39172 3992 39178 4004
rect 41138 3992 41144 4004
rect 39172 3964 41144 3992
rect 39172 3952 39178 3964
rect 41138 3952 41144 3964
rect 41196 3992 41202 4004
rect 42794 3992 42800 4004
rect 41196 3964 42800 3992
rect 41196 3952 41202 3964
rect 42794 3952 42800 3964
rect 42852 3952 42858 4004
rect 43364 3992 43392 4023
rect 43530 4020 43536 4032
rect 43588 4060 43594 4072
rect 43806 4060 43812 4072
rect 43588 4032 43812 4060
rect 43588 4020 43594 4032
rect 43806 4020 43812 4032
rect 43864 4020 43870 4072
rect 44450 4020 44456 4072
rect 44508 4060 44514 4072
rect 45281 4063 45339 4069
rect 45281 4060 45293 4063
rect 44508 4032 45293 4060
rect 44508 4020 44514 4032
rect 45281 4029 45293 4032
rect 45327 4029 45339 4063
rect 45281 4023 45339 4029
rect 45370 4020 45376 4072
rect 45428 4060 45434 4072
rect 45428 4032 51074 4060
rect 45428 4020 45434 4032
rect 44542 3992 44548 4004
rect 43364 3964 44548 3992
rect 44542 3952 44548 3964
rect 44600 3952 44606 4004
rect 44726 3952 44732 4004
rect 44784 3992 44790 4004
rect 45646 3992 45652 4004
rect 44784 3964 45652 3992
rect 44784 3952 44790 3964
rect 45646 3952 45652 3964
rect 45704 3952 45710 4004
rect 46566 3952 46572 4004
rect 46624 3992 46630 4004
rect 50890 3992 50896 4004
rect 46624 3964 50896 3992
rect 46624 3952 46630 3964
rect 50890 3952 50896 3964
rect 50948 3952 50954 4004
rect 51046 3992 51074 4032
rect 54294 4020 54300 4072
rect 54352 4060 54358 4072
rect 55140 4060 55168 4091
rect 57974 4088 57980 4100
rect 58032 4088 58038 4140
rect 58342 4128 58348 4140
rect 58303 4100 58348 4128
rect 58342 4088 58348 4100
rect 58400 4088 58406 4140
rect 54352 4032 55168 4060
rect 57057 4063 57115 4069
rect 54352 4020 54358 4032
rect 57057 4029 57069 4063
rect 57103 4060 57115 4063
rect 58250 4060 58256 4072
rect 57103 4032 58256 4060
rect 57103 4029 57115 4032
rect 57057 4023 57115 4029
rect 58250 4020 58256 4032
rect 58308 4020 58314 4072
rect 55306 3992 55312 4004
rect 51046 3964 54708 3992
rect 55267 3964 55312 3992
rect 38746 3924 38752 3936
rect 37792 3896 38056 3924
rect 38707 3896 38752 3924
rect 37792 3884 37798 3896
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 38838 3884 38844 3936
rect 38896 3924 38902 3936
rect 39942 3924 39948 3936
rect 38896 3896 39948 3924
rect 38896 3884 38902 3896
rect 39942 3884 39948 3896
rect 40000 3884 40006 3936
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 41693 3927 41751 3933
rect 41693 3924 41705 3927
rect 41472 3896 41705 3924
rect 41472 3884 41478 3896
rect 41693 3893 41705 3896
rect 41739 3893 41751 3927
rect 42812 3924 42840 3952
rect 43530 3924 43536 3936
rect 42812 3896 43536 3924
rect 41693 3887 41751 3893
rect 43530 3884 43536 3896
rect 43588 3884 43594 3936
rect 43622 3884 43628 3936
rect 43680 3924 43686 3936
rect 44453 3927 44511 3933
rect 44453 3924 44465 3927
rect 43680 3896 44465 3924
rect 43680 3884 43686 3896
rect 44453 3893 44465 3896
rect 44499 3893 44511 3927
rect 44453 3887 44511 3893
rect 48593 3927 48651 3933
rect 48593 3893 48605 3927
rect 48639 3924 48651 3927
rect 51534 3924 51540 3936
rect 48639 3896 51540 3924
rect 48639 3893 48651 3896
rect 48593 3887 48651 3893
rect 51534 3884 51540 3896
rect 51592 3884 51598 3936
rect 54680 3924 54708 3964
rect 55306 3952 55312 3964
rect 55364 3952 55370 4004
rect 57425 3927 57483 3933
rect 57425 3924 57437 3927
rect 54680 3896 57437 3924
rect 57425 3893 57437 3896
rect 57471 3893 57483 3927
rect 57425 3887 57483 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 5718 3720 5724 3732
rect 3252 3692 5724 3720
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 3142 3516 3148 3528
rect 1627 3488 3148 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3252 3525 3280 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 14090 3720 14096 3732
rect 7248 3692 9720 3720
rect 7248 3680 7254 3692
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 5074 3652 5080 3664
rect 4212 3624 5080 3652
rect 4212 3612 4218 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5445 3655 5503 3661
rect 5445 3621 5457 3655
rect 5491 3652 5503 3655
rect 8389 3655 8447 3661
rect 8389 3652 8401 3655
rect 5491 3624 8401 3652
rect 5491 3621 5503 3624
rect 5445 3615 5503 3621
rect 8389 3621 8401 3624
rect 8435 3621 8447 3655
rect 8389 3615 8447 3621
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 9122 3652 9128 3664
rect 8720 3624 9128 3652
rect 8720 3612 8726 3624
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 9692 3661 9720 3692
rect 9876 3692 14096 3720
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3621 9735 3655
rect 9677 3615 9735 3621
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 5994 3584 6000 3596
rect 4755 3556 6000 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7006 3584 7012 3596
rect 6963 3556 7012 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 9876 3584 9904 3692
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 16025 3723 16083 3729
rect 16025 3689 16037 3723
rect 16071 3720 16083 3723
rect 17586 3720 17592 3732
rect 16071 3692 17592 3720
rect 16071 3689 16083 3692
rect 16025 3683 16083 3689
rect 17586 3680 17592 3692
rect 17644 3720 17650 3732
rect 19334 3720 19340 3732
rect 17644 3692 19340 3720
rect 17644 3680 17650 3692
rect 19334 3680 19340 3692
rect 19392 3720 19398 3732
rect 22922 3720 22928 3732
rect 19392 3692 19656 3720
rect 22883 3692 22928 3720
rect 19392 3680 19398 3692
rect 10318 3612 10324 3664
rect 10376 3612 10382 3664
rect 11514 3652 11520 3664
rect 11475 3624 11520 3652
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 11701 3655 11759 3661
rect 11701 3621 11713 3655
rect 11747 3652 11759 3655
rect 11882 3652 11888 3664
rect 11747 3624 11888 3652
rect 11747 3621 11759 3624
rect 11701 3615 11759 3621
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 14918 3652 14924 3664
rect 12406 3624 14924 3652
rect 7340 3556 9904 3584
rect 10336 3584 10364 3612
rect 10597 3587 10655 3593
rect 10336 3556 10548 3584
rect 7340 3544 7346 3556
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 4982 3516 4988 3528
rect 3467 3488 4988 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 7374 3516 7380 3528
rect 5307 3488 7380 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 9950 3516 9956 3528
rect 7515 3488 9956 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10410 3516 10416 3528
rect 10367 3488 10416 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10520 3516 10548 3556
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 12406 3584 12434 3624
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 18138 3652 18144 3664
rect 16816 3624 18144 3652
rect 16816 3612 16822 3624
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 18840 3624 19441 3652
rect 18840 3612 18846 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19429 3615 19487 3621
rect 10643 3556 12434 3584
rect 12621 3587 12679 3593
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 15746 3584 15752 3596
rect 12667 3556 15752 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 17678 3584 17684 3596
rect 17420 3556 17684 3584
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 10520 3488 11253 3516
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 4525 3451 4583 3457
rect 4525 3417 4537 3451
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3448 6055 3451
rect 6043 3420 6684 3448
rect 6043 3417 6055 3420
rect 5997 3411 6055 3417
rect 4540 3380 4568 3411
rect 5902 3380 5908 3392
rect 4540 3352 5908 3380
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6086 3380 6092 3392
rect 6047 3352 6092 3380
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6656 3380 6684 3420
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 6788 3420 6833 3448
rect 7392 3420 8064 3448
rect 6788 3408 6794 3420
rect 7392 3380 7420 3420
rect 7558 3380 7564 3392
rect 6656 3352 7420 3380
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8036 3380 8064 3420
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 8846 3448 8852 3460
rect 8168 3420 8213 3448
rect 8496 3420 8852 3448
rect 8168 3408 8174 3420
rect 8496 3380 8524 3420
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 9401 3451 9459 3457
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10520 3448 10548 3488
rect 11241 3485 11253 3488
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 13170 3516 13176 3528
rect 12391 3488 13176 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13630 3516 13636 3528
rect 13311 3488 13636 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14516 3488 14749 3516
rect 14516 3476 14522 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3516 15071 3519
rect 16577 3519 16635 3525
rect 15059 3488 16528 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 9447 3420 10548 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 12158 3408 12164 3460
rect 12216 3448 12222 3460
rect 13446 3448 13452 3460
rect 12216 3420 13452 3448
rect 12216 3408 12222 3420
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 13541 3451 13599 3457
rect 13541 3417 13553 3451
rect 13587 3448 13599 3451
rect 15749 3451 15807 3457
rect 13587 3420 14780 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 8036 3352 8524 3380
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8662 3380 8668 3392
rect 8619 3352 8668 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 14550 3380 14556 3392
rect 9907 3352 14556 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14752 3380 14780 3420
rect 15749 3417 15761 3451
rect 15795 3448 15807 3451
rect 15838 3448 15844 3460
rect 15795 3420 15844 3448
rect 15795 3417 15807 3420
rect 15749 3411 15807 3417
rect 15838 3408 15844 3420
rect 15896 3448 15902 3460
rect 16206 3448 16212 3460
rect 15896 3420 16212 3448
rect 15896 3408 15902 3420
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 16500 3448 16528 3488
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 17420 3516 17448 3556
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3584 17831 3587
rect 19242 3584 19248 3596
rect 17819 3556 19248 3584
rect 17819 3553 17831 3556
rect 17773 3547 17831 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19628 3584 19656 3692
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 24029 3723 24087 3729
rect 24029 3689 24041 3723
rect 24075 3720 24087 3723
rect 24394 3720 24400 3732
rect 24075 3692 24400 3720
rect 24075 3689 24087 3692
rect 24029 3683 24087 3689
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24578 3720 24584 3732
rect 24539 3692 24584 3720
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 24854 3680 24860 3732
rect 24912 3720 24918 3732
rect 29178 3720 29184 3732
rect 24912 3692 29184 3720
rect 24912 3680 24918 3692
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 31386 3720 31392 3732
rect 29748 3692 31392 3720
rect 19702 3612 19708 3664
rect 19760 3652 19766 3664
rect 23382 3652 23388 3664
rect 19760 3624 20852 3652
rect 19760 3612 19766 3624
rect 19628 3556 19758 3584
rect 16623 3488 17448 3516
rect 17497 3519 17555 3525
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 18046 3516 18052 3528
rect 17543 3488 18052 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18414 3516 18420 3528
rect 18375 3488 18420 3516
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 19334 3516 19340 3528
rect 18739 3488 19340 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 16758 3448 16764 3460
rect 16500 3420 16764 3448
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 16853 3451 16911 3457
rect 16853 3417 16865 3451
rect 16899 3448 16911 3451
rect 18966 3448 18972 3460
rect 16899 3420 18972 3448
rect 16899 3417 16911 3420
rect 16853 3411 16911 3417
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 19730 3448 19758 3556
rect 19978 3544 19984 3596
rect 20036 3544 20042 3596
rect 20824 3584 20852 3624
rect 21836 3624 23388 3652
rect 21836 3584 21864 3624
rect 23382 3612 23388 3624
rect 23440 3612 23446 3664
rect 28350 3612 28356 3664
rect 28408 3652 28414 3664
rect 29748 3652 29776 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 34238 3720 34244 3732
rect 31864 3692 34244 3720
rect 28408 3624 29776 3652
rect 28408 3612 28414 3624
rect 20824 3556 21864 3584
rect 19994 3457 20022 3544
rect 20824 3528 20852 3556
rect 20622 3516 20628 3528
rect 20583 3488 20628 3516
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20806 3516 20812 3528
rect 20719 3488 20812 3516
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20898 3476 20904 3528
rect 20956 3476 20962 3528
rect 21836 3525 21864 3556
rect 22833 3587 22891 3593
rect 22833 3553 22845 3587
rect 22879 3584 22891 3587
rect 23014 3584 23020 3596
rect 22879 3556 23020 3584
rect 22879 3553 22891 3556
rect 22833 3547 22891 3553
rect 23014 3544 23020 3556
rect 23072 3544 23078 3596
rect 23661 3587 23719 3593
rect 23661 3553 23673 3587
rect 23707 3584 23719 3587
rect 24670 3584 24676 3596
rect 23707 3556 24676 3584
rect 23707 3553 23719 3556
rect 23661 3547 23719 3553
rect 24670 3544 24676 3556
rect 24728 3584 24734 3596
rect 25133 3587 25191 3593
rect 25133 3584 25145 3587
rect 24728 3556 25145 3584
rect 24728 3544 24734 3556
rect 25133 3553 25145 3556
rect 25179 3553 25191 3587
rect 25774 3584 25780 3596
rect 25735 3556 25780 3584
rect 25133 3547 25191 3553
rect 21821 3519 21879 3525
rect 21821 3485 21833 3519
rect 21867 3485 21879 3519
rect 21821 3479 21879 3485
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22336 3488 22661 3516
rect 22336 3476 22342 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 22925 3519 22983 3525
rect 22925 3485 22937 3519
rect 22971 3516 22983 3519
rect 23198 3516 23204 3528
rect 22971 3488 23204 3516
rect 22971 3485 22983 3488
rect 22925 3479 22983 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 24854 3516 24860 3528
rect 23891 3488 24860 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 25148 3516 25176 3547
rect 25774 3544 25780 3556
rect 25832 3544 25838 3596
rect 27985 3587 28043 3593
rect 27985 3553 27997 3587
rect 28031 3584 28043 3587
rect 29454 3584 29460 3596
rect 28031 3556 29460 3584
rect 28031 3553 28043 3556
rect 27985 3547 28043 3553
rect 29454 3544 29460 3556
rect 29512 3544 29518 3596
rect 29546 3544 29552 3596
rect 29604 3584 29610 3596
rect 29730 3584 29736 3596
rect 29604 3556 29736 3584
rect 29604 3544 29610 3556
rect 29730 3544 29736 3556
rect 29788 3544 29794 3596
rect 25682 3516 25688 3528
rect 25148 3488 25688 3516
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 26044 3519 26102 3525
rect 26044 3485 26056 3519
rect 26090 3516 26102 3519
rect 27154 3516 27160 3528
rect 26090 3488 27160 3516
rect 26090 3485 26102 3488
rect 26044 3479 26102 3485
rect 27154 3476 27160 3488
rect 27212 3476 27218 3528
rect 27246 3476 27252 3528
rect 27304 3516 27310 3528
rect 27709 3519 27767 3525
rect 27709 3516 27721 3519
rect 27304 3488 27721 3516
rect 27304 3476 27310 3488
rect 27709 3485 27721 3488
rect 27755 3485 27767 3519
rect 29037 3519 29095 3525
rect 29037 3516 29049 3519
rect 27709 3479 27767 3485
rect 28184 3488 29049 3516
rect 19981 3451 20039 3457
rect 19730 3420 19840 3448
rect 19058 3380 19064 3392
rect 14752 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 19702 3380 19708 3392
rect 19663 3352 19708 3380
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 19812 3389 19840 3420
rect 19981 3417 19993 3451
rect 20027 3417 20039 3451
rect 20714 3448 20720 3460
rect 19981 3411 20039 3417
rect 20272 3420 20720 3448
rect 19797 3383 19855 3389
rect 19797 3349 19809 3383
rect 19843 3380 19855 3383
rect 20272 3380 20300 3420
rect 20714 3408 20720 3420
rect 20772 3448 20778 3460
rect 20916 3448 20944 3476
rect 20772 3420 21036 3448
rect 20772 3408 20778 3420
rect 19843 3352 20300 3380
rect 20349 3383 20407 3389
rect 19843 3349 19855 3352
rect 19797 3343 19855 3349
rect 20349 3349 20361 3383
rect 20395 3380 20407 3383
rect 20898 3380 20904 3392
rect 20395 3352 20904 3380
rect 20395 3349 20407 3352
rect 20349 3343 20407 3349
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21008 3389 21036 3420
rect 21082 3408 21088 3460
rect 21140 3448 21146 3460
rect 21177 3451 21235 3457
rect 21177 3448 21189 3451
rect 21140 3420 21189 3448
rect 21140 3408 21146 3420
rect 21177 3417 21189 3420
rect 21223 3417 21235 3451
rect 21634 3448 21640 3460
rect 21595 3420 21640 3448
rect 21177 3411 21235 3417
rect 21634 3408 21640 3420
rect 21692 3408 21698 3460
rect 22023 3451 22081 3457
rect 22023 3448 22035 3451
rect 21836 3420 22035 3448
rect 20993 3383 21051 3389
rect 20993 3349 21005 3383
rect 21039 3380 21051 3383
rect 21836 3380 21864 3420
rect 22023 3417 22035 3420
rect 22069 3417 22081 3451
rect 22023 3411 22081 3417
rect 22186 3408 22192 3460
rect 22244 3448 22250 3460
rect 25041 3451 25099 3457
rect 22244 3420 22289 3448
rect 22244 3408 22250 3420
rect 25041 3417 25053 3451
rect 25087 3448 25099 3451
rect 26970 3448 26976 3460
rect 25087 3420 26976 3448
rect 25087 3417 25099 3420
rect 25041 3411 25099 3417
rect 26970 3408 26976 3420
rect 27028 3408 27034 3460
rect 27522 3408 27528 3460
rect 27580 3448 27586 3460
rect 28184 3448 28212 3488
rect 29037 3485 29049 3488
rect 29083 3516 29095 3519
rect 30926 3516 30932 3528
rect 29083 3488 30932 3516
rect 29083 3485 29095 3488
rect 29037 3479 29095 3485
rect 30926 3476 30932 3488
rect 30984 3516 30990 3528
rect 31864 3516 31892 3692
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 34422 3680 34428 3732
rect 34480 3720 34486 3732
rect 35894 3720 35900 3732
rect 34480 3692 35900 3720
rect 34480 3680 34486 3692
rect 35894 3680 35900 3692
rect 35952 3680 35958 3732
rect 36170 3680 36176 3732
rect 36228 3720 36234 3732
rect 36265 3723 36323 3729
rect 36265 3720 36277 3723
rect 36228 3692 36277 3720
rect 36228 3680 36234 3692
rect 36265 3689 36277 3692
rect 36311 3689 36323 3723
rect 36265 3683 36323 3689
rect 36446 3680 36452 3732
rect 36504 3720 36510 3732
rect 38933 3723 38991 3729
rect 38933 3720 38945 3723
rect 36504 3692 38945 3720
rect 36504 3680 36510 3692
rect 38933 3689 38945 3692
rect 38979 3689 38991 3723
rect 38933 3683 38991 3689
rect 39022 3680 39028 3732
rect 39080 3720 39086 3732
rect 41966 3720 41972 3732
rect 39080 3692 41414 3720
rect 41927 3692 41972 3720
rect 39080 3680 39086 3692
rect 33226 3612 33232 3664
rect 33284 3652 33290 3664
rect 33413 3655 33471 3661
rect 33413 3652 33425 3655
rect 33284 3624 33425 3652
rect 33284 3612 33290 3624
rect 33413 3621 33425 3624
rect 33459 3621 33471 3655
rect 33413 3615 33471 3621
rect 36078 3612 36084 3664
rect 36136 3652 36142 3664
rect 37182 3652 37188 3664
rect 36136 3624 37188 3652
rect 36136 3612 36142 3624
rect 37182 3612 37188 3624
rect 37240 3612 37246 3664
rect 37274 3612 37280 3664
rect 37332 3652 37338 3664
rect 37369 3655 37427 3661
rect 37369 3652 37381 3655
rect 37332 3624 37381 3652
rect 37332 3612 37338 3624
rect 37369 3621 37381 3624
rect 37415 3621 37427 3655
rect 37369 3615 37427 3621
rect 37550 3612 37556 3664
rect 37608 3652 37614 3664
rect 40494 3652 40500 3664
rect 37608 3624 40500 3652
rect 37608 3612 37614 3624
rect 40494 3612 40500 3624
rect 40552 3612 40558 3664
rect 40678 3612 40684 3664
rect 40736 3612 40742 3664
rect 41386 3652 41414 3692
rect 41966 3680 41972 3692
rect 42024 3680 42030 3732
rect 43070 3680 43076 3732
rect 43128 3720 43134 3732
rect 45094 3720 45100 3732
rect 43128 3692 45100 3720
rect 43128 3680 43134 3692
rect 45094 3680 45100 3692
rect 45152 3680 45158 3732
rect 45186 3680 45192 3732
rect 45244 3720 45250 3732
rect 45373 3723 45431 3729
rect 45373 3720 45385 3723
rect 45244 3692 45385 3720
rect 45244 3680 45250 3692
rect 45373 3689 45385 3692
rect 45419 3689 45431 3723
rect 45373 3683 45431 3689
rect 46014 3680 46020 3732
rect 46072 3720 46078 3732
rect 46109 3723 46167 3729
rect 46109 3720 46121 3723
rect 46072 3692 46121 3720
rect 46072 3680 46078 3692
rect 46109 3689 46121 3692
rect 46155 3689 46167 3723
rect 47857 3723 47915 3729
rect 47857 3720 47869 3723
rect 46109 3683 46167 3689
rect 46216 3692 47869 3720
rect 43993 3655 44051 3661
rect 43993 3652 44005 3655
rect 41386 3624 44005 3652
rect 43993 3621 44005 3624
rect 44039 3621 44051 3655
rect 46216 3652 46244 3692
rect 47857 3689 47869 3692
rect 47903 3689 47915 3723
rect 48590 3720 48596 3732
rect 48551 3692 48596 3720
rect 47857 3683 47915 3689
rect 48590 3680 48596 3692
rect 48648 3680 48654 3732
rect 49326 3720 49332 3732
rect 49287 3692 49332 3720
rect 49326 3680 49332 3692
rect 49384 3680 49390 3732
rect 50062 3680 50068 3732
rect 50120 3720 50126 3732
rect 50525 3723 50583 3729
rect 50525 3720 50537 3723
rect 50120 3692 50537 3720
rect 50120 3680 50126 3692
rect 50525 3689 50537 3692
rect 50571 3689 50583 3723
rect 51994 3720 52000 3732
rect 51955 3692 52000 3720
rect 50525 3683 50583 3689
rect 51994 3680 52000 3692
rect 52052 3680 52058 3732
rect 52638 3680 52644 3732
rect 52696 3720 52702 3732
rect 54205 3723 54263 3729
rect 54205 3720 54217 3723
rect 52696 3692 54217 3720
rect 52696 3680 52702 3692
rect 54205 3689 54217 3692
rect 54251 3689 54263 3723
rect 54205 3683 54263 3689
rect 47026 3652 47032 3664
rect 43993 3615 44051 3621
rect 44468 3624 46244 3652
rect 46987 3624 47032 3652
rect 34882 3584 34888 3596
rect 33060 3556 34888 3584
rect 30984 3488 31892 3516
rect 32033 3519 32091 3525
rect 30984 3476 30990 3488
rect 32033 3485 32045 3519
rect 32079 3516 32091 3519
rect 33060 3516 33088 3556
rect 34882 3544 34888 3556
rect 34940 3544 34946 3596
rect 35894 3544 35900 3596
rect 35952 3584 35958 3596
rect 36998 3584 37004 3596
rect 35952 3556 37004 3584
rect 35952 3544 35958 3556
rect 36998 3544 37004 3556
rect 37056 3544 37062 3596
rect 38654 3584 38660 3596
rect 37844 3556 38660 3584
rect 32079 3488 33088 3516
rect 33873 3519 33931 3525
rect 32079 3485 32091 3488
rect 32033 3479 32091 3485
rect 32416 3460 32444 3488
rect 33873 3485 33885 3519
rect 33919 3516 33931 3519
rect 35152 3519 35210 3525
rect 33919 3488 35112 3516
rect 33919 3485 33931 3488
rect 33873 3479 33931 3485
rect 27580 3420 28212 3448
rect 27580 3408 27586 3420
rect 28258 3408 28264 3460
rect 28316 3448 28322 3460
rect 28534 3448 28540 3460
rect 28316 3420 28540 3448
rect 28316 3408 28322 3420
rect 28534 3408 28540 3420
rect 28592 3448 28598 3460
rect 28813 3451 28871 3457
rect 28813 3448 28825 3451
rect 28592 3420 28825 3448
rect 28592 3408 28598 3420
rect 28813 3417 28825 3420
rect 28859 3417 28871 3451
rect 28813 3411 28871 3417
rect 29181 3451 29239 3457
rect 29181 3417 29193 3451
rect 29227 3448 29239 3451
rect 29546 3448 29552 3460
rect 29227 3420 29552 3448
rect 29227 3417 29239 3420
rect 29181 3411 29239 3417
rect 29546 3408 29552 3420
rect 29604 3408 29610 3460
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 32306 3457 32312 3460
rect 30000 3451 30058 3457
rect 30000 3448 30012 3451
rect 29880 3420 30012 3448
rect 29880 3408 29886 3420
rect 30000 3417 30012 3420
rect 30046 3417 30058 3451
rect 32300 3448 32312 3457
rect 32267 3420 32312 3448
rect 30000 3411 30058 3417
rect 32300 3411 32312 3420
rect 32306 3408 32312 3411
rect 32364 3408 32370 3460
rect 32398 3408 32404 3460
rect 32456 3408 32462 3460
rect 32858 3408 32864 3460
rect 32916 3448 32922 3460
rect 34149 3451 34207 3457
rect 34149 3448 34161 3451
rect 32916 3420 34161 3448
rect 32916 3408 32922 3420
rect 34149 3417 34161 3420
rect 34195 3417 34207 3451
rect 35084 3448 35112 3488
rect 35152 3485 35164 3519
rect 35198 3516 35210 3519
rect 36078 3516 36084 3528
rect 35198 3488 36084 3516
rect 35198 3485 35210 3488
rect 35152 3479 35210 3485
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 36722 3516 36728 3528
rect 36683 3488 36728 3516
rect 36722 3476 36728 3488
rect 36780 3476 36786 3528
rect 36906 3525 36912 3528
rect 36873 3519 36912 3525
rect 36873 3485 36885 3519
rect 36873 3479 36912 3485
rect 36906 3476 36912 3479
rect 36964 3476 36970 3528
rect 37231 3519 37289 3525
rect 37231 3485 37243 3519
rect 37277 3516 37289 3519
rect 37734 3516 37740 3528
rect 37277 3488 37740 3516
rect 37277 3485 37289 3488
rect 37231 3479 37289 3485
rect 37734 3476 37740 3488
rect 37792 3476 37798 3528
rect 37844 3525 37872 3556
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 40313 3587 40371 3593
rect 40313 3553 40325 3587
rect 40359 3584 40371 3587
rect 40696 3584 40724 3612
rect 40359 3556 40724 3584
rect 40773 3587 40831 3593
rect 40359 3553 40371 3556
rect 40313 3547 40371 3553
rect 40773 3553 40785 3587
rect 40819 3584 40831 3587
rect 42610 3584 42616 3596
rect 40819 3556 42616 3584
rect 40819 3553 40831 3556
rect 40773 3547 40831 3553
rect 42610 3544 42616 3556
rect 42668 3544 42674 3596
rect 43162 3544 43168 3596
rect 43220 3584 43226 3596
rect 44468 3584 44496 3624
rect 47026 3612 47032 3624
rect 47084 3612 47090 3664
rect 49694 3612 49700 3664
rect 49752 3652 49758 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 49752 3624 52837 3652
rect 49752 3612 49758 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 52825 3615 52883 3621
rect 58253 3655 58311 3661
rect 58253 3621 58265 3655
rect 58299 3621 58311 3655
rect 58253 3615 58311 3621
rect 43220 3556 44496 3584
rect 43220 3544 43226 3556
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 51353 3587 51411 3593
rect 51353 3584 51365 3587
rect 44600 3556 51365 3584
rect 44600 3544 44606 3556
rect 51353 3553 51365 3556
rect 51399 3553 51411 3587
rect 51353 3547 51411 3553
rect 51534 3544 51540 3596
rect 51592 3584 51598 3596
rect 56870 3584 56876 3596
rect 51592 3556 54340 3584
rect 56831 3556 56876 3584
rect 51592 3544 51598 3556
rect 37829 3519 37887 3525
rect 37829 3485 37841 3519
rect 37875 3485 37887 3519
rect 40681 3519 40739 3525
rect 37829 3479 37887 3485
rect 38028 3488 40264 3516
rect 36630 3448 36636 3460
rect 35084 3420 36636 3448
rect 34149 3411 34207 3417
rect 36630 3408 36636 3420
rect 36688 3408 36694 3460
rect 36998 3448 37004 3460
rect 36959 3420 37004 3448
rect 36998 3408 37004 3420
rect 37056 3408 37062 3460
rect 37093 3451 37151 3457
rect 37093 3417 37105 3451
rect 37139 3448 37151 3451
rect 38028 3448 38056 3488
rect 37139 3420 38056 3448
rect 38105 3451 38163 3457
rect 37139 3417 37151 3420
rect 37093 3411 37151 3417
rect 38105 3417 38117 3451
rect 38151 3417 38163 3451
rect 38105 3411 38163 3417
rect 21039 3352 21864 3380
rect 21913 3383 21971 3389
rect 21039 3349 21051 3352
rect 20993 3343 21051 3349
rect 21913 3349 21925 3383
rect 21959 3380 21971 3383
rect 22462 3380 22468 3392
rect 21959 3352 22468 3380
rect 21959 3349 21971 3352
rect 21913 3343 21971 3349
rect 22462 3340 22468 3352
rect 22520 3340 22526 3392
rect 23106 3380 23112 3392
rect 23067 3352 23112 3380
rect 23106 3340 23112 3352
rect 23164 3340 23170 3392
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 23934 3380 23940 3392
rect 23256 3352 23940 3380
rect 23256 3340 23262 3352
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 24949 3383 25007 3389
rect 24949 3349 24961 3383
rect 24995 3380 25007 3383
rect 25222 3380 25228 3392
rect 24995 3352 25228 3380
rect 24995 3349 25007 3352
rect 24949 3343 25007 3349
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 27157 3383 27215 3389
rect 27157 3380 27169 3383
rect 26384 3352 27169 3380
rect 26384 3340 26390 3352
rect 27157 3349 27169 3352
rect 27203 3380 27215 3383
rect 27614 3380 27620 3392
rect 27203 3352 27620 3380
rect 27203 3349 27215 3352
rect 27157 3343 27215 3349
rect 27614 3340 27620 3352
rect 27672 3340 27678 3392
rect 28626 3340 28632 3392
rect 28684 3380 28690 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 28684 3352 28733 3380
rect 28684 3340 28690 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 28905 3383 28963 3389
rect 28905 3349 28917 3383
rect 28951 3380 28963 3383
rect 28994 3380 29000 3392
rect 28951 3352 29000 3380
rect 28951 3349 28963 3352
rect 28905 3343 28963 3349
rect 28994 3340 29000 3352
rect 29052 3340 29058 3392
rect 30190 3340 30196 3392
rect 30248 3380 30254 3392
rect 31113 3383 31171 3389
rect 31113 3380 31125 3383
rect 30248 3352 31125 3380
rect 30248 3340 30254 3352
rect 31113 3349 31125 3352
rect 31159 3349 31171 3383
rect 31113 3343 31171 3349
rect 35250 3340 35256 3392
rect 35308 3380 35314 3392
rect 38120 3380 38148 3411
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 38562 3448 38568 3460
rect 38436 3420 38568 3448
rect 38436 3408 38442 3420
rect 38562 3408 38568 3420
rect 38620 3408 38626 3460
rect 38654 3408 38660 3460
rect 38712 3448 38718 3460
rect 38841 3451 38899 3457
rect 38841 3448 38853 3451
rect 38712 3420 38853 3448
rect 38712 3408 38718 3420
rect 38841 3417 38853 3420
rect 38887 3417 38899 3451
rect 38841 3411 38899 3417
rect 38930 3408 38936 3460
rect 38988 3448 38994 3460
rect 40126 3448 40132 3460
rect 38988 3420 40132 3448
rect 38988 3408 38994 3420
rect 40126 3408 40132 3420
rect 40184 3408 40190 3460
rect 35308 3352 38148 3380
rect 35308 3340 35314 3352
rect 38286 3340 38292 3392
rect 38344 3380 38350 3392
rect 39574 3380 39580 3392
rect 38344 3352 39580 3380
rect 38344 3340 38350 3352
rect 39574 3340 39580 3352
rect 39632 3340 39638 3392
rect 40236 3380 40264 3488
rect 40681 3485 40693 3519
rect 40727 3485 40739 3519
rect 41046 3516 41052 3528
rect 41007 3488 41052 3516
rect 40681 3479 40739 3485
rect 40696 3448 40724 3479
rect 41046 3476 41052 3488
rect 41104 3476 41110 3528
rect 41138 3476 41144 3528
rect 41196 3516 41202 3528
rect 42150 3516 42156 3528
rect 41196 3488 41241 3516
rect 42111 3488 42156 3516
rect 41196 3476 41202 3488
rect 42150 3476 42156 3488
rect 42208 3476 42214 3528
rect 42337 3519 42395 3525
rect 42337 3485 42349 3519
rect 42383 3485 42395 3519
rect 42702 3516 42708 3528
rect 42663 3488 42708 3516
rect 42337 3479 42395 3485
rect 41322 3448 41328 3460
rect 40696 3420 41328 3448
rect 41322 3408 41328 3420
rect 41380 3448 41386 3460
rect 42352 3448 42380 3479
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 42794 3476 42800 3528
rect 42852 3516 42858 3528
rect 42852 3488 42897 3516
rect 42852 3476 42858 3488
rect 43346 3476 43352 3528
rect 43404 3516 43410 3528
rect 43530 3525 43536 3528
rect 43497 3519 43536 3525
rect 43404 3488 43449 3516
rect 43404 3476 43410 3488
rect 43497 3485 43509 3519
rect 43497 3479 43536 3485
rect 43530 3476 43536 3479
rect 43588 3476 43594 3528
rect 43806 3476 43812 3528
rect 43864 3525 43870 3528
rect 43864 3516 43872 3525
rect 45002 3516 45008 3528
rect 43864 3488 43909 3516
rect 44468 3488 45008 3516
rect 43864 3479 43872 3488
rect 43864 3476 43870 3479
rect 43254 3448 43260 3460
rect 41380 3420 43260 3448
rect 41380 3408 41386 3420
rect 43254 3408 43260 3420
rect 43312 3448 43318 3460
rect 43625 3451 43683 3457
rect 43625 3448 43637 3451
rect 43312 3420 43637 3448
rect 43312 3408 43318 3420
rect 43625 3417 43637 3420
rect 43671 3417 43683 3451
rect 43625 3411 43683 3417
rect 43717 3451 43775 3457
rect 43717 3417 43729 3451
rect 43763 3448 43775 3451
rect 44468 3448 44496 3488
rect 45002 3476 45008 3488
rect 45060 3476 45066 3528
rect 46014 3516 46020 3528
rect 45975 3488 46020 3516
rect 46014 3476 46020 3488
rect 46072 3476 46078 3528
rect 48501 3519 48559 3525
rect 48501 3516 48513 3519
rect 46124 3488 48513 3516
rect 43763 3420 44496 3448
rect 43763 3417 43775 3420
rect 43717 3411 43775 3417
rect 44542 3408 44548 3460
rect 44600 3448 44606 3460
rect 45281 3451 45339 3457
rect 45281 3448 45293 3451
rect 44600 3420 45293 3448
rect 44600 3408 44606 3420
rect 45281 3417 45293 3420
rect 45327 3417 45339 3451
rect 45281 3411 45339 3417
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 46124 3448 46152 3488
rect 48501 3485 48513 3488
rect 48547 3485 48559 3519
rect 48501 3479 48559 3485
rect 49142 3476 49148 3528
rect 49200 3516 49206 3528
rect 49200 3488 49464 3516
rect 49200 3476 49206 3488
rect 45520 3420 46152 3448
rect 45520 3408 45526 3420
rect 46658 3408 46664 3460
rect 46716 3448 46722 3460
rect 46845 3451 46903 3457
rect 46845 3448 46857 3451
rect 46716 3420 46857 3448
rect 46716 3408 46722 3420
rect 46845 3417 46857 3420
rect 46891 3417 46903 3451
rect 46845 3411 46903 3417
rect 47118 3408 47124 3460
rect 47176 3448 47182 3460
rect 47765 3451 47823 3457
rect 47765 3448 47777 3451
rect 47176 3420 47777 3448
rect 47176 3408 47182 3420
rect 47765 3417 47777 3420
rect 47811 3417 47823 3451
rect 47765 3411 47823 3417
rect 48130 3408 48136 3460
rect 48188 3448 48194 3460
rect 49237 3451 49295 3457
rect 49237 3448 49249 3451
rect 48188 3420 49249 3448
rect 48188 3408 48194 3420
rect 49237 3417 49249 3420
rect 49283 3417 49295 3451
rect 49237 3411 49295 3417
rect 45186 3380 45192 3392
rect 40236 3352 45192 3380
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 49436 3380 49464 3488
rect 50706 3476 50712 3528
rect 50764 3516 50770 3528
rect 51169 3519 51227 3525
rect 51169 3516 51181 3519
rect 50764 3488 51181 3516
rect 50764 3476 50770 3488
rect 51169 3485 51181 3488
rect 51215 3485 51227 3519
rect 51905 3519 51963 3525
rect 51905 3516 51917 3519
rect 51169 3479 51227 3485
rect 51460 3488 51917 3516
rect 49510 3408 49516 3460
rect 49568 3448 49574 3460
rect 50433 3451 50491 3457
rect 50433 3448 50445 3451
rect 49568 3420 50445 3448
rect 49568 3408 49574 3420
rect 50433 3417 50445 3420
rect 50479 3417 50491 3451
rect 50433 3411 50491 3417
rect 50798 3408 50804 3460
rect 50856 3448 50862 3460
rect 51460 3448 51488 3488
rect 51905 3485 51917 3488
rect 51951 3485 51963 3519
rect 51905 3479 51963 3485
rect 51994 3476 52000 3528
rect 52052 3516 52058 3528
rect 53377 3519 53435 3525
rect 53377 3516 53389 3519
rect 52052 3488 53389 3516
rect 52052 3476 52058 3488
rect 53377 3485 53389 3488
rect 53423 3485 53435 3519
rect 53377 3479 53435 3485
rect 50856 3420 51488 3448
rect 50856 3408 50862 3420
rect 51626 3408 51632 3460
rect 51684 3448 51690 3460
rect 52641 3451 52699 3457
rect 52641 3448 52653 3451
rect 51684 3420 52653 3448
rect 51684 3408 51690 3420
rect 52641 3417 52653 3420
rect 52687 3417 52699 3451
rect 52641 3411 52699 3417
rect 52730 3408 52736 3460
rect 52788 3448 52794 3460
rect 53926 3448 53932 3460
rect 52788 3420 53932 3448
rect 52788 3408 52794 3420
rect 53926 3408 53932 3420
rect 53984 3408 53990 3460
rect 54113 3451 54171 3457
rect 54113 3417 54125 3451
rect 54159 3417 54171 3451
rect 54113 3411 54171 3417
rect 51810 3380 51816 3392
rect 49436 3352 51816 3380
rect 51810 3340 51816 3352
rect 51868 3340 51874 3392
rect 53466 3380 53472 3392
rect 53427 3352 53472 3380
rect 53466 3340 53472 3352
rect 53524 3340 53530 3392
rect 53650 3340 53656 3392
rect 53708 3380 53714 3392
rect 54128 3380 54156 3411
rect 53708 3352 54156 3380
rect 54312 3380 54340 3556
rect 56870 3544 56876 3556
rect 56928 3544 56934 3596
rect 55953 3519 56011 3525
rect 55953 3485 55965 3519
rect 55999 3516 56011 3519
rect 58268 3516 58296 3615
rect 55999 3488 58296 3516
rect 55999 3485 56011 3488
rect 55953 3479 56011 3485
rect 56226 3448 56232 3460
rect 56187 3420 56232 3448
rect 56226 3408 56232 3420
rect 56284 3408 56290 3460
rect 57118 3451 57176 3457
rect 57118 3448 57130 3451
rect 56336 3420 57130 3448
rect 56336 3380 56364 3420
rect 57118 3417 57130 3420
rect 57164 3417 57176 3451
rect 57118 3411 57176 3417
rect 54312 3352 56364 3380
rect 53708 3340 53714 3352
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 4154 3176 4160 3188
rect 3007 3148 4160 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 6546 3176 6552 3188
rect 4479 3148 6552 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9030 3176 9036 3188
rect 8435 3148 9036 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 17678 3176 17684 3188
rect 9140 3148 17684 3176
rect 4798 3108 4804 3120
rect 1596 3080 4804 3108
rect 1596 3049 1624 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 5077 3111 5135 3117
rect 5077 3077 5089 3111
rect 5123 3108 5135 3111
rect 7282 3108 7288 3120
rect 5123 3080 7144 3108
rect 7243 3080 7288 3108
rect 5123 3077 5135 3080
rect 5077 3071 5135 3077
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 1581 3003 1639 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4706 3040 4712 3052
rect 4387 3012 4712 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5815 3043 5873 3049
rect 5815 3009 5827 3043
rect 5861 3040 5873 3043
rect 7116 3040 7144 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 7929 3111 7987 3117
rect 7929 3077 7941 3111
rect 7975 3108 7987 3111
rect 8110 3108 8116 3120
rect 7975 3080 8116 3108
rect 7975 3077 7987 3080
rect 7929 3071 7987 3077
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 9140 3117 9168 3148
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 18782 3176 18788 3188
rect 17828 3148 18788 3176
rect 17828 3136 17834 3148
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 20901 3179 20959 3185
rect 19300 3148 20852 3176
rect 19300 3136 19306 3148
rect 9125 3111 9183 3117
rect 9125 3077 9137 3111
rect 9171 3077 9183 3111
rect 9125 3071 9183 3077
rect 10045 3111 10103 3117
rect 10045 3077 10057 3111
rect 10091 3108 10103 3111
rect 15013 3111 15071 3117
rect 10091 3080 14872 3108
rect 10091 3077 10103 3080
rect 10045 3071 10103 3077
rect 8849 3043 8907 3049
rect 5861 3012 6592 3040
rect 7116 3012 8432 3040
rect 5861 3009 5873 3012
rect 5815 3003 5873 3009
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 6564 2972 6592 3012
rect 8404 2972 8432 3012
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 9214 3040 9220 3052
rect 8895 3012 9220 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10226 3040 10232 3052
rect 9815 3012 10232 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10686 3040 10692 3052
rect 10647 3012 10692 3040
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 12158 3040 12164 3052
rect 12119 3012 12164 3040
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12526 3040 12532 3052
rect 12483 3012 12532 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13722 3040 13728 3052
rect 13127 3012 13728 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13964 3012 14013 3040
rect 13964 3000 13970 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14734 3040 14740 3052
rect 14001 3003 14059 3009
rect 14108 3012 14596 3040
rect 14695 3012 14740 3040
rect 10134 2972 10140 2984
rect 6564 2944 8340 2972
rect 8404 2944 10140 2972
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 8205 2907 8263 2913
rect 8205 2904 8217 2907
rect 6144 2876 8217 2904
rect 6144 2864 6150 2876
rect 8205 2873 8217 2876
rect 8251 2873 8263 2907
rect 8205 2867 8263 2873
rect 3694 2836 3700 2848
rect 3655 2808 3700 2836
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 5166 2836 5172 2848
rect 5127 2808 5172 2836
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5868 2808 5917 2836
rect 5868 2796 5874 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 8312 2836 8340 2944
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 13357 2975 13415 2981
rect 11011 2944 12480 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 12066 2904 12072 2916
rect 9916 2876 12072 2904
rect 9916 2864 9922 2876
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 12452 2904 12480 2944
rect 13357 2941 13369 2975
rect 13403 2972 13415 2975
rect 14108 2972 14136 3012
rect 14274 2972 14280 2984
rect 13403 2944 14136 2972
rect 14235 2944 14280 2972
rect 13403 2941 13415 2944
rect 13357 2935 13415 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14568 2972 14596 3012
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14844 3040 14872 3080
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 16574 3108 16580 3120
rect 15059 3080 16580 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 16758 3068 16764 3120
rect 16816 3108 16822 3120
rect 19061 3111 19119 3117
rect 16816 3080 19012 3108
rect 16816 3068 16822 3080
rect 15194 3040 15200 3052
rect 14844 3012 15200 3040
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 15841 3003 15899 3009
rect 15286 2972 15292 2984
rect 14568 2944 15292 2972
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 15470 2904 15476 2916
rect 12452 2876 15476 2904
rect 15470 2864 15476 2876
rect 15528 2864 15534 2916
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2904 15623 2907
rect 15856 2904 15884 3003
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 18785 3043 18843 3049
rect 17328 3012 18736 3040
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 17328 2972 17356 3012
rect 16163 2944 17356 2972
rect 17405 2975 17463 2981
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 17405 2941 17417 2975
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 16942 2904 16948 2916
rect 15611 2876 16948 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17420 2904 17448 2935
rect 18046 2932 18052 2984
rect 18104 2972 18110 2984
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 18104 2944 18337 2972
rect 18104 2932 18110 2944
rect 18325 2941 18337 2944
rect 18371 2941 18383 2975
rect 18708 2972 18736 3012
rect 18785 3009 18797 3043
rect 18831 3040 18843 3043
rect 18874 3040 18880 3052
rect 18831 3012 18880 3040
rect 18831 3009 18843 3012
rect 18785 3003 18843 3009
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 18984 3040 19012 3080
rect 19061 3077 19073 3111
rect 19107 3108 19119 3111
rect 20438 3108 20444 3120
rect 19107 3080 20444 3108
rect 19107 3077 19119 3080
rect 19061 3071 19119 3077
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 20824 3108 20852 3148
rect 20901 3145 20913 3179
rect 20947 3176 20959 3179
rect 20990 3176 20996 3188
rect 20947 3148 20996 3176
rect 20947 3145 20959 3148
rect 20901 3139 20959 3145
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 23017 3179 23075 3185
rect 21100 3148 22876 3176
rect 21100 3108 21128 3148
rect 20824 3080 21128 3108
rect 21177 3111 21235 3117
rect 21177 3077 21189 3111
rect 21223 3108 21235 3111
rect 21358 3108 21364 3120
rect 21223 3080 21364 3108
rect 21223 3077 21235 3080
rect 21177 3071 21235 3077
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 22097 3111 22155 3117
rect 22097 3108 22109 3111
rect 21508 3080 22109 3108
rect 21508 3068 21514 3080
rect 22097 3077 22109 3080
rect 22143 3108 22155 3111
rect 22554 3108 22560 3120
rect 22143 3080 22560 3108
rect 22143 3077 22155 3080
rect 22097 3071 22155 3077
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 19518 3040 19524 3052
rect 18984 3012 19524 3040
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19702 3040 19708 3052
rect 19663 3012 19708 3040
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 19852 3012 20484 3040
rect 19852 3000 19858 3012
rect 19978 2972 19984 2984
rect 18708 2944 19840 2972
rect 19939 2944 19984 2972
rect 18325 2935 18383 2941
rect 19812 2904 19840 2944
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20346 2904 20352 2916
rect 17420 2876 19748 2904
rect 19812 2876 20352 2904
rect 11054 2836 11060 2848
rect 8312 2808 11060 2836
rect 5905 2799 5963 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 15010 2836 15016 2848
rect 14608 2808 15016 2836
rect 14608 2796 14614 2808
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 19426 2836 19432 2848
rect 15436 2808 19432 2836
rect 15436 2796 15442 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 19720 2836 19748 2876
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 20456 2904 20484 3012
rect 20530 3000 20536 3052
rect 20588 3040 20594 3052
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 20588 3012 20637 3040
rect 20588 3000 20594 3012
rect 20625 3009 20637 3012
rect 20671 3009 20683 3043
rect 20806 3040 20812 3052
rect 20767 3012 20812 3040
rect 20625 3003 20683 3009
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 21033 3043 21091 3049
rect 21033 3009 21045 3043
rect 21079 3009 21091 3043
rect 21033 3003 21091 3009
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21048 2972 21076 3003
rect 21358 2972 21364 2984
rect 20772 2944 21364 2972
rect 20772 2932 20778 2944
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 22848 2972 22876 3148
rect 23017 3145 23029 3179
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 23032 3108 23060 3139
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 23164 3148 23209 3176
rect 23164 3136 23170 3148
rect 23566 3136 23572 3188
rect 23624 3176 23630 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 23624 3148 24409 3176
rect 23624 3136 23630 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 25133 3179 25191 3185
rect 25133 3145 25145 3179
rect 25179 3176 25191 3179
rect 25406 3176 25412 3188
rect 25179 3148 25412 3176
rect 25179 3145 25191 3148
rect 25133 3139 25191 3145
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 25498 3136 25504 3188
rect 25556 3176 25562 3188
rect 25556 3148 25601 3176
rect 25556 3136 25562 3148
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 28721 3179 28779 3185
rect 28721 3176 28733 3179
rect 27488 3148 28733 3176
rect 27488 3136 27494 3148
rect 26326 3108 26332 3120
rect 23032 3080 26332 3108
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 26421 3111 26479 3117
rect 26421 3077 26433 3111
rect 26467 3108 26479 3111
rect 27614 3108 27620 3120
rect 26467 3080 27620 3108
rect 26467 3077 26479 3080
rect 26421 3071 26479 3077
rect 27614 3068 27620 3080
rect 27672 3068 27678 3120
rect 27724 3117 27752 3148
rect 28721 3145 28733 3148
rect 28767 3145 28779 3179
rect 28721 3139 28779 3145
rect 29178 3136 29184 3188
rect 29236 3176 29242 3188
rect 29546 3176 29552 3188
rect 29236 3148 29552 3176
rect 29236 3136 29242 3148
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 29822 3136 29828 3188
rect 29880 3176 29886 3188
rect 29917 3179 29975 3185
rect 29917 3176 29929 3179
rect 29880 3148 29929 3176
rect 29880 3136 29886 3148
rect 29917 3145 29929 3148
rect 29963 3145 29975 3179
rect 29917 3139 29975 3145
rect 30006 3136 30012 3188
rect 30064 3176 30070 3188
rect 30285 3179 30343 3185
rect 30285 3176 30297 3179
rect 30064 3148 30297 3176
rect 30064 3136 30070 3148
rect 30285 3145 30297 3148
rect 30331 3145 30343 3179
rect 32030 3176 32036 3188
rect 30285 3139 30343 3145
rect 30392 3148 32036 3176
rect 27709 3111 27767 3117
rect 27709 3077 27721 3111
rect 27755 3077 27767 3111
rect 27709 3071 27767 3077
rect 28258 3068 28264 3120
rect 28316 3108 28322 3120
rect 28537 3111 28595 3117
rect 28537 3108 28549 3111
rect 28316 3080 28549 3108
rect 28316 3068 28322 3080
rect 28537 3077 28549 3080
rect 28583 3077 28595 3111
rect 28537 3071 28595 3077
rect 28905 3111 28963 3117
rect 28905 3077 28917 3111
rect 28951 3108 28963 3111
rect 30392 3108 30420 3148
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 33226 3136 33232 3188
rect 33284 3176 33290 3188
rect 36078 3176 36084 3188
rect 33284 3148 36084 3176
rect 33284 3136 33290 3148
rect 36078 3136 36084 3148
rect 36136 3136 36142 3188
rect 36262 3176 36268 3188
rect 36223 3148 36268 3176
rect 36262 3136 36268 3148
rect 36320 3136 36326 3188
rect 36446 3136 36452 3188
rect 36504 3176 36510 3188
rect 39482 3176 39488 3188
rect 36504 3148 38792 3176
rect 39443 3148 39488 3176
rect 36504 3136 36510 3148
rect 28951 3080 30420 3108
rect 28951 3077 28963 3080
rect 28905 3071 28963 3077
rect 30466 3068 30472 3120
rect 30524 3068 30530 3120
rect 30742 3068 30748 3120
rect 30800 3108 30806 3120
rect 30800 3080 32444 3108
rect 30800 3068 30806 3080
rect 22922 3000 22928 3052
rect 22980 3040 22986 3052
rect 23290 3040 23296 3052
rect 22980 3012 23025 3040
rect 23251 3012 23296 3040
rect 22980 3000 22986 3012
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 24084 3012 24317 3040
rect 24084 3000 24090 3012
rect 24305 3009 24317 3012
rect 24351 3009 24363 3043
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 24305 3003 24363 3009
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 28350 3040 28356 3052
rect 27540 3012 28356 3040
rect 23750 2972 23756 2984
rect 22848 2944 23756 2972
rect 23750 2932 23756 2944
rect 23808 2932 23814 2984
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2941 24639 2975
rect 25590 2972 25596 2984
rect 25551 2944 25596 2972
rect 24581 2935 24639 2941
rect 20806 2904 20812 2916
rect 20456 2876 20812 2904
rect 20806 2864 20812 2876
rect 20864 2864 20870 2916
rect 22281 2907 22339 2913
rect 22281 2873 22293 2907
rect 22327 2904 22339 2907
rect 22462 2904 22468 2916
rect 22327 2876 22468 2904
rect 22327 2873 22339 2876
rect 22281 2867 22339 2873
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 22738 2904 22744 2916
rect 22699 2876 22744 2904
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 23937 2907 23995 2913
rect 23937 2873 23949 2907
rect 23983 2904 23995 2907
rect 24394 2904 24400 2916
rect 23983 2876 24400 2904
rect 23983 2873 23995 2876
rect 23937 2867 23995 2873
rect 24394 2864 24400 2876
rect 24452 2864 24458 2916
rect 24596 2904 24624 2935
rect 25590 2932 25596 2944
rect 25648 2932 25654 2984
rect 25682 2932 25688 2984
rect 25740 2972 25746 2984
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25740 2944 25789 2972
rect 25740 2932 25746 2944
rect 25777 2941 25789 2944
rect 25823 2972 25835 2975
rect 27540 2972 27568 3012
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 28675 3043 28733 3049
rect 28675 3009 28687 3043
rect 28721 3040 28733 3043
rect 29914 3040 29920 3052
rect 28721 3012 29920 3040
rect 28721 3009 28733 3012
rect 28675 3003 28733 3009
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 30282 3040 30288 3052
rect 30116 3012 30288 3040
rect 30116 2972 30144 3012
rect 30282 3000 30288 3012
rect 30340 3000 30346 3052
rect 25823 2944 27568 2972
rect 28184 2944 30144 2972
rect 25823 2941 25835 2944
rect 25777 2935 25835 2941
rect 25700 2904 25728 2932
rect 28184 2904 28212 2944
rect 30190 2932 30196 2984
rect 30248 2972 30254 2984
rect 30377 2975 30435 2981
rect 30377 2972 30389 2975
rect 30248 2944 30389 2972
rect 30248 2932 30254 2944
rect 30377 2941 30389 2944
rect 30423 2941 30435 2975
rect 30484 2972 30512 3068
rect 31294 3040 31300 3052
rect 31255 3012 31300 3040
rect 31294 3000 31300 3012
rect 31352 3000 31358 3052
rect 32306 3040 32312 3052
rect 32267 3012 32312 3040
rect 32306 3000 32312 3012
rect 32364 3000 32370 3052
rect 32416 3040 32444 3080
rect 32490 3068 32496 3120
rect 32548 3108 32554 3120
rect 33505 3111 33563 3117
rect 33505 3108 33517 3111
rect 32548 3080 33517 3108
rect 32548 3068 32554 3080
rect 33505 3077 33517 3080
rect 33551 3077 33563 3111
rect 33505 3071 33563 3077
rect 33962 3068 33968 3120
rect 34020 3108 34026 3120
rect 35152 3111 35210 3117
rect 34020 3080 35020 3108
rect 34020 3068 34026 3080
rect 33229 3043 33287 3049
rect 33229 3040 33241 3043
rect 32416 3012 33241 3040
rect 33229 3009 33241 3012
rect 33275 3040 33287 3043
rect 34146 3040 34152 3052
rect 33275 3012 34152 3040
rect 33275 3009 33287 3012
rect 33229 3003 33287 3009
rect 34146 3000 34152 3012
rect 34204 3000 34210 3052
rect 34241 3043 34299 3049
rect 34241 3009 34253 3043
rect 34287 3009 34299 3043
rect 34422 3040 34428 3052
rect 34383 3012 34428 3040
rect 34241 3003 34299 3009
rect 30561 2975 30619 2981
rect 30561 2972 30573 2975
rect 30484 2944 30573 2972
rect 30377 2935 30435 2941
rect 30561 2941 30573 2944
rect 30607 2941 30619 2975
rect 30561 2935 30619 2941
rect 31202 2932 31208 2984
rect 31260 2972 31266 2984
rect 31481 2975 31539 2981
rect 31481 2972 31493 2975
rect 31260 2944 31493 2972
rect 31260 2932 31266 2944
rect 31481 2941 31493 2944
rect 31527 2941 31539 2975
rect 31481 2935 31539 2941
rect 31754 2932 31760 2984
rect 31812 2972 31818 2984
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31812 2944 32505 2972
rect 31812 2932 31818 2944
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 32493 2935 32551 2941
rect 28350 2904 28356 2916
rect 24596 2876 25728 2904
rect 26712 2876 28212 2904
rect 28311 2876 28356 2904
rect 22370 2836 22376 2848
rect 19720 2808 22376 2836
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 26712 2836 26740 2876
rect 28350 2864 28356 2876
rect 28408 2864 28414 2916
rect 28626 2864 28632 2916
rect 28684 2904 28690 2916
rect 34256 2904 34284 3003
rect 34422 3000 34428 3012
rect 34480 3000 34486 3052
rect 34882 3040 34888 3052
rect 34843 3012 34888 3040
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 34992 3040 35020 3080
rect 35152 3077 35164 3111
rect 35198 3108 35210 3111
rect 35342 3108 35348 3120
rect 35198 3080 35348 3108
rect 35198 3077 35210 3080
rect 35152 3071 35210 3077
rect 35342 3068 35348 3080
rect 35400 3068 35406 3120
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 38657 3111 38715 3117
rect 38657 3108 38669 3111
rect 35492 3080 38669 3108
rect 35492 3068 35498 3080
rect 38657 3077 38669 3080
rect 38703 3077 38715 3111
rect 38764 3108 38792 3148
rect 39482 3136 39488 3148
rect 39540 3136 39546 3188
rect 40586 3176 40592 3188
rect 40547 3148 40592 3176
rect 40586 3136 40592 3148
rect 40644 3136 40650 3188
rect 41138 3136 41144 3188
rect 41196 3176 41202 3188
rect 44453 3179 44511 3185
rect 41196 3148 44312 3176
rect 41196 3136 41202 3148
rect 41233 3111 41291 3117
rect 41233 3108 41245 3111
rect 38764 3080 41245 3108
rect 38657 3071 38715 3077
rect 41233 3077 41245 3080
rect 41279 3077 41291 3111
rect 41233 3071 41291 3077
rect 41417 3111 41475 3117
rect 41417 3077 41429 3111
rect 41463 3108 41475 3111
rect 41874 3108 41880 3120
rect 41463 3080 41880 3108
rect 41463 3077 41475 3080
rect 41417 3071 41475 3077
rect 41874 3068 41880 3080
rect 41932 3068 41938 3120
rect 42426 3068 42432 3120
rect 42484 3108 42490 3120
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 42484 3080 42625 3108
rect 42484 3068 42490 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 42613 3071 42671 3077
rect 43180 3080 43760 3108
rect 37461 3043 37519 3049
rect 34992 3012 35940 3040
rect 35912 2972 35940 3012
rect 37461 3009 37473 3043
rect 37507 3040 37519 3043
rect 38194 3040 38200 3052
rect 37507 3012 38200 3040
rect 37507 3009 37519 3012
rect 37461 3003 37519 3009
rect 38194 3000 38200 3012
rect 38252 3000 38258 3052
rect 38381 3043 38439 3049
rect 38381 3009 38393 3043
rect 38427 3040 38439 3043
rect 38838 3040 38844 3052
rect 38427 3012 38844 3040
rect 38427 3009 38439 3012
rect 38381 3003 38439 3009
rect 38838 3000 38844 3012
rect 38896 3000 38902 3052
rect 39114 3000 39120 3052
rect 39172 3040 39178 3052
rect 39393 3043 39451 3049
rect 39393 3040 39405 3043
rect 39172 3012 39405 3040
rect 39172 3000 39178 3012
rect 39393 3009 39405 3012
rect 39439 3009 39451 3043
rect 39393 3003 39451 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 40313 3043 40371 3049
rect 40313 3040 40325 3043
rect 39816 3012 40325 3040
rect 39816 3000 39822 3012
rect 40313 3009 40325 3012
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 37645 2975 37703 2981
rect 37645 2972 37657 2975
rect 35912 2944 37657 2972
rect 37645 2941 37657 2944
rect 37691 2941 37703 2975
rect 38286 2972 38292 2984
rect 37645 2935 37703 2941
rect 37752 2944 38292 2972
rect 28684 2876 34284 2904
rect 28684 2864 28690 2876
rect 36538 2864 36544 2916
rect 36596 2904 36602 2916
rect 37752 2904 37780 2944
rect 38286 2932 38292 2944
rect 38344 2932 38350 2984
rect 36596 2876 37780 2904
rect 36596 2864 36602 2876
rect 37826 2864 37832 2916
rect 37884 2904 37890 2916
rect 43180 2904 43208 3080
rect 43254 3000 43260 3052
rect 43312 3040 43318 3052
rect 43622 3040 43628 3052
rect 43312 3012 43357 3040
rect 43583 3012 43628 3040
rect 43312 3000 43318 3012
rect 43622 3000 43628 3012
rect 43680 3000 43686 3052
rect 43349 2975 43407 2981
rect 43349 2941 43361 2975
rect 43395 2941 43407 2975
rect 43732 2972 43760 3080
rect 43806 3000 43812 3052
rect 43864 3040 43870 3052
rect 44284 3049 44312 3148
rect 44453 3145 44465 3179
rect 44499 3176 44511 3179
rect 44634 3176 44640 3188
rect 44499 3148 44640 3176
rect 44499 3145 44511 3148
rect 44453 3139 44511 3145
rect 44634 3136 44640 3148
rect 44692 3136 44698 3188
rect 45186 3176 45192 3188
rect 45147 3148 45192 3176
rect 45186 3136 45192 3148
rect 45244 3136 45250 3188
rect 46382 3176 46388 3188
rect 46343 3148 46388 3176
rect 46382 3136 46388 3148
rect 46440 3136 46446 3188
rect 47394 3136 47400 3188
rect 47452 3176 47458 3188
rect 47949 3179 48007 3185
rect 47949 3176 47961 3179
rect 47452 3148 47961 3176
rect 47452 3136 47458 3148
rect 47949 3145 47961 3148
rect 47995 3145 48007 3179
rect 47949 3139 48007 3145
rect 48038 3136 48044 3188
rect 48096 3176 48102 3188
rect 49789 3179 49847 3185
rect 49789 3176 49801 3179
rect 48096 3148 49801 3176
rect 48096 3136 48102 3148
rect 49789 3145 49801 3148
rect 49835 3145 49847 3179
rect 49789 3139 49847 3145
rect 50246 3136 50252 3188
rect 50304 3176 50310 3188
rect 50706 3176 50712 3188
rect 50304 3148 50712 3176
rect 50304 3136 50310 3148
rect 50706 3136 50712 3148
rect 50764 3136 50770 3188
rect 51258 3176 51264 3188
rect 51219 3148 51264 3176
rect 51258 3136 51264 3148
rect 51316 3136 51322 3188
rect 51810 3136 51816 3188
rect 51868 3176 51874 3188
rect 53834 3176 53840 3188
rect 51868 3148 53052 3176
rect 53795 3148 53840 3176
rect 51868 3136 51874 3148
rect 45462 3108 45468 3120
rect 44468 3080 45468 3108
rect 44468 3052 44496 3080
rect 45462 3068 45468 3080
rect 45520 3068 45526 3120
rect 47486 3068 47492 3120
rect 47544 3108 47550 3120
rect 49697 3111 49755 3117
rect 49697 3108 49709 3111
rect 47544 3080 49709 3108
rect 47544 3068 47550 3080
rect 49697 3077 49709 3080
rect 49743 3077 49755 3111
rect 49697 3071 49755 3077
rect 49878 3068 49884 3120
rect 49936 3108 49942 3120
rect 53024 3117 53052 3148
rect 53834 3136 53840 3148
rect 53892 3136 53898 3188
rect 54754 3176 54760 3188
rect 54715 3148 54760 3176
rect 54754 3136 54760 3148
rect 54812 3136 54818 3188
rect 58250 3176 58256 3188
rect 58211 3148 58256 3176
rect 58250 3136 58256 3148
rect 58308 3136 58314 3188
rect 51905 3111 51963 3117
rect 51905 3108 51917 3111
rect 49936 3080 51917 3108
rect 49936 3068 49942 3080
rect 51905 3077 51917 3080
rect 51951 3077 51963 3111
rect 51905 3071 51963 3077
rect 53009 3111 53067 3117
rect 53009 3077 53021 3111
rect 53055 3077 53067 3111
rect 53650 3108 53656 3120
rect 53009 3071 53067 3077
rect 53116 3080 53656 3108
rect 44269 3043 44327 3049
rect 43864 3012 43909 3040
rect 43864 3000 43870 3012
rect 44269 3009 44281 3043
rect 44315 3009 44327 3043
rect 44269 3003 44327 3009
rect 44450 3000 44456 3052
rect 44508 3000 44514 3052
rect 45097 3043 45155 3049
rect 45097 3009 45109 3043
rect 45143 3009 45155 3043
rect 45097 3003 45155 3009
rect 45112 2972 45140 3003
rect 46106 3000 46112 3052
rect 46164 3040 46170 3052
rect 46293 3043 46351 3049
rect 46293 3040 46305 3043
rect 46164 3012 46305 3040
rect 46164 3000 46170 3012
rect 46293 3009 46305 3012
rect 46339 3009 46351 3043
rect 46293 3003 46351 3009
rect 47026 3000 47032 3052
rect 47084 3040 47090 3052
rect 47857 3043 47915 3049
rect 47857 3040 47869 3043
rect 47084 3012 47869 3040
rect 47084 3000 47090 3012
rect 47857 3009 47869 3012
rect 47903 3009 47915 3043
rect 48130 3040 48136 3052
rect 47857 3003 47915 3009
rect 47964 3012 48136 3040
rect 43732 2944 45140 2972
rect 43349 2935 43407 2941
rect 37884 2876 43208 2904
rect 43364 2904 43392 2935
rect 45278 2932 45284 2984
rect 45336 2972 45342 2984
rect 47964 2972 47992 3012
rect 48130 3000 48136 3012
rect 48188 3000 48194 3052
rect 48590 3000 48596 3052
rect 48648 3040 48654 3052
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 48648 3012 48789 3040
rect 48648 3000 48654 3012
rect 48777 3009 48789 3012
rect 48823 3009 48835 3043
rect 48777 3003 48835 3009
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 50433 3043 50491 3049
rect 50433 3040 50445 3043
rect 49016 3012 50445 3040
rect 49016 3000 49022 3012
rect 50433 3009 50445 3012
rect 50479 3009 50491 3043
rect 51077 3043 51135 3049
rect 51077 3040 51089 3043
rect 50433 3003 50491 3009
rect 50540 3012 51089 3040
rect 45336 2944 47992 2972
rect 45336 2932 45342 2944
rect 48038 2932 48044 2984
rect 48096 2972 48102 2984
rect 50540 2972 50568 3012
rect 51077 3009 51089 3012
rect 51123 3009 51135 3043
rect 51077 3003 51135 3009
rect 51166 3000 51172 3052
rect 51224 3040 51230 3052
rect 53116 3040 53144 3080
rect 53650 3068 53656 3080
rect 53708 3068 53714 3120
rect 55674 3068 55680 3120
rect 55732 3108 55738 3120
rect 55769 3111 55827 3117
rect 55769 3108 55781 3111
rect 55732 3080 55781 3108
rect 55732 3068 55738 3080
rect 55769 3077 55781 3080
rect 55815 3077 55827 3111
rect 58158 3108 58164 3120
rect 58119 3080 58164 3108
rect 55769 3071 55827 3077
rect 58158 3068 58164 3080
rect 58216 3068 58222 3120
rect 51224 3012 53144 3040
rect 51224 3000 51230 3012
rect 53558 3000 53564 3052
rect 53616 3040 53622 3052
rect 53745 3043 53803 3049
rect 53745 3040 53757 3043
rect 53616 3012 53757 3040
rect 53616 3000 53622 3012
rect 53745 3009 53757 3012
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 53834 3000 53840 3052
rect 53892 3040 53898 3052
rect 54665 3043 54723 3049
rect 54665 3040 54677 3043
rect 53892 3012 54677 3040
rect 53892 3000 53898 3012
rect 54665 3009 54677 3012
rect 54711 3009 54723 3043
rect 54665 3003 54723 3009
rect 54938 3000 54944 3052
rect 54996 3040 55002 3052
rect 55493 3043 55551 3049
rect 55493 3040 55505 3043
rect 54996 3012 55505 3040
rect 54996 3000 55002 3012
rect 55493 3009 55505 3012
rect 55539 3009 55551 3043
rect 56413 3043 56471 3049
rect 56413 3040 56425 3043
rect 55493 3003 55551 3009
rect 55600 3012 56425 3040
rect 48096 2944 50568 2972
rect 48096 2932 48102 2944
rect 50890 2932 50896 2984
rect 50948 2972 50954 2984
rect 53193 2975 53251 2981
rect 53193 2972 53205 2975
rect 50948 2944 53205 2972
rect 50948 2932 50954 2944
rect 53193 2941 53205 2944
rect 53239 2941 53251 2975
rect 53193 2935 53251 2941
rect 53374 2932 53380 2984
rect 53432 2972 53438 2984
rect 55600 2972 55628 3012
rect 56413 3009 56425 3012
rect 56459 3009 56471 3043
rect 56413 3003 56471 3009
rect 53432 2944 55628 2972
rect 53432 2932 53438 2944
rect 55766 2932 55772 2984
rect 55824 2972 55830 2984
rect 56597 2975 56655 2981
rect 56597 2972 56609 2975
rect 55824 2944 56609 2972
rect 55824 2932 55830 2944
rect 56597 2941 56609 2944
rect 56643 2941 56655 2975
rect 56597 2935 56655 2941
rect 52089 2907 52147 2913
rect 52089 2904 52101 2907
rect 43364 2876 52101 2904
rect 37884 2864 37890 2876
rect 52089 2873 52101 2876
rect 52135 2873 52147 2907
rect 52089 2867 52147 2873
rect 25188 2808 26740 2836
rect 25188 2796 25194 2808
rect 26786 2796 26792 2848
rect 26844 2836 26850 2848
rect 31662 2836 31668 2848
rect 26844 2808 31668 2836
rect 26844 2796 26850 2808
rect 31662 2796 31668 2808
rect 31720 2796 31726 2848
rect 32030 2796 32036 2848
rect 32088 2836 32094 2848
rect 33410 2836 33416 2848
rect 32088 2808 33416 2836
rect 32088 2796 32094 2808
rect 33410 2796 33416 2808
rect 33468 2796 33474 2848
rect 36998 2796 37004 2848
rect 37056 2836 37062 2848
rect 40126 2836 40132 2848
rect 37056 2808 40132 2836
rect 37056 2796 37062 2808
rect 40126 2796 40132 2808
rect 40184 2796 40190 2848
rect 40862 2796 40868 2848
rect 40920 2836 40926 2848
rect 41598 2836 41604 2848
rect 40920 2808 41604 2836
rect 40920 2796 40926 2808
rect 41598 2796 41604 2808
rect 41656 2796 41662 2848
rect 45278 2796 45284 2848
rect 45336 2836 45342 2848
rect 48958 2836 48964 2848
rect 45336 2808 48964 2836
rect 45336 2796 45342 2808
rect 48958 2796 48964 2808
rect 49016 2796 49022 2848
rect 49050 2796 49056 2848
rect 49108 2836 49114 2848
rect 49108 2808 49153 2836
rect 49108 2796 49114 2808
rect 49694 2796 49700 2848
rect 49752 2836 49758 2848
rect 50525 2839 50583 2845
rect 50525 2836 50537 2839
rect 49752 2808 50537 2836
rect 49752 2796 49758 2808
rect 50525 2805 50537 2808
rect 50571 2805 50583 2839
rect 50525 2799 50583 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9582 2632 9588 2644
rect 8619 2604 9588 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 12710 2632 12716 2644
rect 9692 2604 12716 2632
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 7558 2564 7564 2576
rect 4571 2536 7564 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 7653 2567 7711 2573
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 7834 2564 7840 2576
rect 7699 2536 7840 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8478 2564 8484 2576
rect 8439 2536 8484 2564
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 9692 2496 9720 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 14645 2635 14703 2641
rect 14645 2601 14657 2635
rect 14691 2632 14703 2635
rect 14734 2632 14740 2644
rect 14691 2604 14740 2632
rect 14691 2601 14703 2604
rect 14645 2595 14703 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 18046 2592 18052 2644
rect 18104 2632 18110 2644
rect 18966 2632 18972 2644
rect 18104 2604 18972 2632
rect 18104 2592 18110 2604
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 19702 2592 19708 2644
rect 19760 2632 19766 2644
rect 21450 2632 21456 2644
rect 19760 2604 21456 2632
rect 19760 2592 19766 2604
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 23290 2632 23296 2644
rect 21560 2604 23296 2632
rect 10870 2564 10876 2576
rect 6043 2468 9720 2496
rect 9784 2536 10876 2564
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 9306 2428 9312 2440
rect 3283 2400 9168 2428
rect 9267 2400 9312 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2360 4399 2363
rect 4890 2360 4896 2372
rect 4387 2332 4896 2360
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 5074 2360 5080 2372
rect 5035 2332 5080 2360
rect 5074 2320 5080 2332
rect 5132 2320 5138 2372
rect 5810 2360 5816 2372
rect 5771 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 6730 2360 6736 2372
rect 6691 2332 6736 2360
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 7006 2360 7012 2372
rect 6963 2332 7012 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 7469 2363 7527 2369
rect 7469 2329 7481 2363
rect 7515 2329 7527 2363
rect 8110 2360 8116 2372
rect 8071 2332 8116 2360
rect 7469 2323 7527 2329
rect 3326 2292 3332 2304
rect 3287 2264 3332 2292
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 7484 2292 7512 2323
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 9140 2360 9168 2400
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9784 2437 9812 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 11885 2567 11943 2573
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 14550 2564 14556 2576
rect 11931 2536 14556 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 21560 2564 21588 2604
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 24762 2592 24768 2644
rect 24820 2632 24826 2644
rect 25038 2632 25044 2644
rect 24820 2604 25044 2632
rect 24820 2592 24826 2604
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 25133 2635 25191 2641
rect 25133 2601 25145 2635
rect 25179 2632 25191 2635
rect 25498 2632 25504 2644
rect 25179 2604 25504 2632
rect 25179 2601 25191 2604
rect 25133 2595 25191 2601
rect 25498 2592 25504 2604
rect 25556 2592 25562 2644
rect 29362 2632 29368 2644
rect 26206 2604 29368 2632
rect 22002 2564 22008 2576
rect 15068 2536 21588 2564
rect 21963 2536 22008 2564
rect 15068 2524 15074 2536
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 23014 2564 23020 2576
rect 22975 2536 23020 2564
rect 23014 2524 23020 2536
rect 23072 2524 23078 2576
rect 23106 2524 23112 2576
rect 23164 2564 23170 2576
rect 23164 2536 25513 2564
rect 23164 2524 23170 2536
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 12710 2496 12716 2508
rect 10091 2468 12716 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 18046 2496 18052 2508
rect 14139 2468 18052 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 19208 2468 22416 2496
rect 19208 2456 19214 2468
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2397 9827 2431
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 9769 2391 9827 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 12342 2428 12348 2440
rect 12303 2400 12348 2428
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14792 2400 14933 2428
rect 14792 2388 14798 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 15838 2428 15844 2440
rect 15799 2400 15844 2428
rect 14921 2391 14979 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 16390 2428 16396 2440
rect 16080 2400 16396 2428
rect 16080 2388 16086 2400
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 18506 2428 18512 2440
rect 18463 2400 18512 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 19978 2428 19984 2440
rect 18656 2400 19380 2428
rect 19939 2400 19984 2428
rect 18656 2388 18662 2400
rect 9674 2360 9680 2372
rect 9140 2332 9680 2360
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 10962 2360 10968 2372
rect 10923 2332 10968 2360
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 13354 2360 13360 2372
rect 12667 2332 13360 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 13538 2360 13544 2372
rect 13499 2332 13544 2360
rect 13538 2320 13544 2332
rect 13596 2320 13602 2372
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 15930 2360 15936 2372
rect 15243 2332 15936 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 15930 2320 15936 2332
rect 15988 2320 15994 2372
rect 16114 2360 16120 2372
rect 16075 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 17770 2360 17776 2372
rect 17731 2332 17776 2360
rect 17770 2320 17776 2332
rect 17828 2320 17834 2372
rect 18690 2360 18696 2372
rect 18651 2332 18696 2360
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 14366 2292 14372 2304
rect 7484 2264 14372 2292
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 19242 2292 19248 2304
rect 16899 2264 19248 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19352 2292 19380 2400
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20898 2428 20904 2440
rect 20859 2400 20904 2428
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2428 21143 2431
rect 21131 2400 22232 2428
rect 21131 2397 21143 2400
rect 21085 2391 21143 2397
rect 19518 2320 19524 2372
rect 19576 2360 19582 2372
rect 20070 2360 20076 2372
rect 19576 2332 20076 2360
rect 19576 2320 19582 2332
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 20254 2360 20260 2372
rect 20215 2332 20260 2360
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 22204 2369 22232 2400
rect 22278 2388 22284 2440
rect 22336 2437 22342 2440
rect 22336 2431 22359 2437
rect 22347 2397 22359 2431
rect 22388 2428 22416 2468
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 25485 2496 25513 2536
rect 25590 2524 25596 2576
rect 25648 2564 25654 2576
rect 26206 2564 26234 2604
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 31662 2592 31668 2644
rect 31720 2632 31726 2644
rect 33594 2632 33600 2644
rect 31720 2604 33600 2632
rect 31720 2592 31726 2604
rect 33594 2592 33600 2604
rect 33652 2592 33658 2644
rect 34149 2635 34207 2641
rect 34149 2601 34161 2635
rect 34195 2632 34207 2635
rect 34330 2632 34336 2644
rect 34195 2604 34336 2632
rect 34195 2601 34207 2604
rect 34149 2595 34207 2601
rect 34330 2592 34336 2604
rect 34388 2592 34394 2644
rect 37642 2632 37648 2644
rect 34808 2604 37648 2632
rect 33042 2564 33048 2576
rect 25648 2536 26234 2564
rect 28920 2536 33048 2564
rect 25648 2524 25654 2536
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 22520 2468 24900 2496
rect 25485 2468 25697 2496
rect 22520 2456 22526 2468
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22388 2400 22569 2428
rect 22336 2391 22359 2397
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 23198 2428 23204 2440
rect 23159 2400 23204 2428
rect 22557 2391 22615 2397
rect 22336 2388 22342 2391
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 23339 2431 23397 2437
rect 23339 2397 23351 2431
rect 23385 2428 23397 2431
rect 24872 2428 24900 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 26326 2456 26332 2508
rect 26384 2496 26390 2508
rect 26878 2496 26884 2508
rect 26384 2468 26884 2496
rect 26384 2456 26390 2468
rect 26878 2456 26884 2468
rect 26936 2456 26942 2508
rect 27433 2431 27491 2437
rect 27433 2428 27445 2431
rect 23385 2400 24808 2428
rect 24872 2400 27445 2428
rect 23385 2397 23397 2400
rect 23339 2391 23397 2397
rect 21453 2363 21511 2369
rect 21453 2360 21465 2363
rect 20364 2332 21465 2360
rect 20364 2292 20392 2332
rect 21453 2329 21465 2332
rect 21499 2329 21511 2363
rect 21453 2323 21511 2329
rect 22189 2363 22247 2369
rect 22189 2329 22201 2363
rect 22235 2360 22247 2363
rect 23216 2360 23244 2388
rect 23566 2360 23572 2372
rect 22235 2332 23244 2360
rect 23527 2332 23572 2360
rect 22235 2329 22247 2332
rect 22189 2323 22247 2329
rect 23566 2320 23572 2332
rect 23624 2320 23630 2372
rect 24780 2360 24808 2400
rect 27433 2397 27445 2400
rect 27479 2397 27491 2431
rect 27798 2428 27804 2440
rect 27433 2391 27491 2397
rect 27540 2400 27804 2428
rect 26326 2360 26332 2372
rect 24780 2332 26332 2360
rect 26326 2320 26332 2332
rect 26384 2320 26390 2372
rect 26421 2363 26479 2369
rect 26421 2329 26433 2363
rect 26467 2360 26479 2363
rect 27540 2360 27568 2400
rect 27798 2388 27804 2400
rect 27856 2428 27862 2440
rect 28350 2428 28356 2440
rect 27856 2400 28356 2428
rect 27856 2388 27862 2400
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2428 28779 2431
rect 28920 2428 28948 2536
rect 33042 2524 33048 2536
rect 33100 2524 33106 2576
rect 28997 2499 29055 2505
rect 28997 2465 29009 2499
rect 29043 2496 29055 2499
rect 30374 2496 30380 2508
rect 29043 2468 30380 2496
rect 29043 2465 29055 2468
rect 28997 2459 29055 2465
rect 30374 2456 30380 2468
rect 30432 2456 30438 2508
rect 34808 2496 34836 2604
rect 37642 2592 37648 2604
rect 37700 2592 37706 2644
rect 40218 2632 40224 2644
rect 40179 2604 40224 2632
rect 40218 2592 40224 2604
rect 40276 2592 40282 2644
rect 41322 2632 41328 2644
rect 41283 2604 41328 2632
rect 41322 2592 41328 2604
rect 41380 2592 41386 2644
rect 42794 2632 42800 2644
rect 42755 2604 42800 2632
rect 42794 2592 42800 2604
rect 42852 2592 42858 2644
rect 45830 2632 45836 2644
rect 45791 2604 45836 2632
rect 45830 2592 45836 2604
rect 45888 2592 45894 2644
rect 46934 2632 46940 2644
rect 46895 2604 46940 2632
rect 46934 2592 46940 2604
rect 46992 2592 46998 2644
rect 47946 2632 47952 2644
rect 47907 2604 47952 2632
rect 47946 2592 47952 2604
rect 48004 2592 48010 2644
rect 49053 2635 49111 2641
rect 49053 2601 49065 2635
rect 49099 2632 49111 2635
rect 49418 2632 49424 2644
rect 49099 2604 49424 2632
rect 49099 2601 49111 2604
rect 49053 2595 49111 2601
rect 49418 2592 49424 2604
rect 49476 2592 49482 2644
rect 50154 2592 50160 2644
rect 50212 2632 50218 2644
rect 50525 2635 50583 2641
rect 50525 2632 50537 2635
rect 50212 2604 50537 2632
rect 50212 2592 50218 2604
rect 50525 2601 50537 2604
rect 50571 2601 50583 2635
rect 54018 2632 54024 2644
rect 53979 2604 54024 2632
rect 50525 2595 50583 2601
rect 54018 2592 54024 2604
rect 54076 2592 54082 2644
rect 57974 2592 57980 2644
rect 58032 2632 58038 2644
rect 58253 2635 58311 2641
rect 58253 2632 58265 2635
rect 58032 2604 58265 2632
rect 58032 2592 58038 2604
rect 58253 2601 58265 2604
rect 58299 2601 58311 2635
rect 58253 2595 58311 2601
rect 37274 2564 37280 2576
rect 33428 2468 34836 2496
rect 34900 2536 37280 2564
rect 28767 2400 28948 2428
rect 28767 2397 28779 2400
rect 28721 2391 28779 2397
rect 29270 2388 29276 2440
rect 29328 2428 29334 2440
rect 30101 2431 30159 2437
rect 30101 2428 30113 2431
rect 29328 2400 30113 2428
rect 29328 2388 29334 2400
rect 30101 2397 30113 2400
rect 30147 2397 30159 2431
rect 30101 2391 30159 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2428 31079 2431
rect 31938 2428 31944 2440
rect 31067 2400 31944 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31938 2388 31944 2400
rect 31996 2388 32002 2440
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2428 32367 2431
rect 32766 2428 32772 2440
rect 32355 2400 32772 2428
rect 32355 2397 32367 2400
rect 32309 2391 32367 2397
rect 32766 2388 32772 2400
rect 32824 2388 32830 2440
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2428 33287 2431
rect 33428 2428 33456 2468
rect 33275 2400 33456 2428
rect 33275 2397 33287 2400
rect 33229 2391 33287 2397
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 34149 2431 34207 2437
rect 34149 2428 34161 2431
rect 34112 2400 34161 2428
rect 34112 2388 34118 2400
rect 34149 2397 34161 2400
rect 34195 2397 34207 2431
rect 34149 2391 34207 2397
rect 34238 2388 34244 2440
rect 34296 2428 34302 2440
rect 34900 2437 34928 2536
rect 37274 2524 37280 2536
rect 37332 2524 37338 2576
rect 38470 2564 38476 2576
rect 37384 2536 38476 2564
rect 36078 2496 36084 2508
rect 36039 2468 36084 2496
rect 36078 2456 36084 2468
rect 36136 2456 36142 2508
rect 34333 2431 34391 2437
rect 34333 2428 34345 2431
rect 34296 2400 34345 2428
rect 34296 2388 34302 2400
rect 34333 2397 34345 2400
rect 34379 2397 34391 2431
rect 34333 2391 34391 2397
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2428 35863 2431
rect 37384 2428 37412 2536
rect 38470 2524 38476 2536
rect 38528 2524 38534 2576
rect 38562 2524 38568 2576
rect 38620 2564 38626 2576
rect 38620 2536 44220 2564
rect 38620 2524 38626 2536
rect 38746 2496 38752 2508
rect 37476 2468 38752 2496
rect 37476 2437 37504 2468
rect 38746 2456 38752 2468
rect 38804 2456 38810 2508
rect 40126 2456 40132 2508
rect 40184 2496 40190 2508
rect 40184 2468 42656 2496
rect 40184 2456 40190 2468
rect 35851 2400 37412 2428
rect 37461 2431 37519 2437
rect 35851 2397 35863 2400
rect 35805 2391 35863 2397
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 41414 2428 41420 2440
rect 38427 2400 41420 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 41414 2388 41420 2400
rect 41472 2388 41478 2440
rect 42628 2437 42656 2468
rect 44192 2437 44220 2536
rect 44358 2456 44364 2508
rect 44416 2496 44422 2508
rect 52089 2499 52147 2505
rect 52089 2496 52101 2499
rect 44416 2468 52101 2496
rect 44416 2456 44422 2468
rect 52089 2465 52101 2468
rect 52135 2465 52147 2499
rect 52089 2459 52147 2465
rect 55398 2456 55404 2508
rect 55456 2496 55462 2508
rect 55677 2499 55735 2505
rect 55677 2496 55689 2499
rect 55456 2468 55689 2496
rect 55456 2456 55462 2468
rect 55677 2465 55689 2468
rect 55723 2465 55735 2499
rect 55677 2459 55735 2465
rect 42613 2431 42671 2437
rect 42613 2397 42625 2431
rect 42659 2397 42671 2431
rect 44177 2431 44235 2437
rect 42613 2391 42671 2397
rect 42720 2400 43576 2428
rect 26467 2332 27568 2360
rect 27709 2363 27767 2369
rect 26467 2329 26479 2332
rect 26421 2323 26479 2329
rect 27709 2329 27721 2363
rect 27755 2360 27767 2363
rect 29822 2360 29828 2372
rect 27755 2332 29828 2360
rect 27755 2329 27767 2332
rect 27709 2323 27767 2329
rect 29822 2320 29828 2332
rect 29880 2320 29886 2372
rect 30377 2363 30435 2369
rect 30377 2329 30389 2363
rect 30423 2360 30435 2363
rect 30650 2360 30656 2372
rect 30423 2332 30656 2360
rect 30423 2329 30435 2332
rect 30377 2323 30435 2329
rect 30650 2320 30656 2332
rect 30708 2320 30714 2372
rect 30926 2320 30932 2372
rect 30984 2360 30990 2372
rect 31297 2363 31355 2369
rect 31297 2360 31309 2363
rect 30984 2332 31309 2360
rect 30984 2320 30990 2332
rect 31297 2329 31309 2332
rect 31343 2329 31355 2363
rect 31297 2323 31355 2329
rect 31478 2320 31484 2372
rect 31536 2360 31542 2372
rect 32585 2363 32643 2369
rect 32585 2360 32597 2363
rect 31536 2332 32597 2360
rect 31536 2320 31542 2332
rect 32585 2329 32597 2332
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 33505 2363 33563 2369
rect 33505 2329 33517 2363
rect 33551 2329 33563 2363
rect 33505 2323 33563 2329
rect 21174 2292 21180 2304
rect 19352 2264 20392 2292
rect 21135 2264 21180 2292
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 21269 2295 21327 2301
rect 21269 2261 21281 2295
rect 21315 2292 21327 2295
rect 21358 2292 21364 2304
rect 21315 2264 21364 2292
rect 21315 2261 21327 2264
rect 21269 2255 21327 2261
rect 21358 2252 21364 2264
rect 21416 2292 21422 2304
rect 22373 2295 22431 2301
rect 22373 2292 22385 2295
rect 21416 2264 22385 2292
rect 21416 2252 21422 2264
rect 22373 2261 22385 2264
rect 22419 2292 22431 2295
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 22419 2264 23397 2292
rect 22419 2261 22431 2264
rect 22373 2255 22431 2261
rect 23385 2261 23397 2264
rect 23431 2261 23443 2295
rect 23385 2255 23443 2261
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 25501 2295 25559 2301
rect 25501 2292 25513 2295
rect 23532 2264 25513 2292
rect 23532 2252 23538 2264
rect 25501 2261 25513 2264
rect 25547 2261 25559 2295
rect 25501 2255 25559 2261
rect 25590 2252 25596 2304
rect 25648 2292 25654 2304
rect 26510 2292 26516 2304
rect 25648 2264 25693 2292
rect 26471 2264 26516 2292
rect 25648 2252 25654 2264
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 32030 2252 32036 2304
rect 32088 2292 32094 2304
rect 33520 2292 33548 2323
rect 33778 2320 33784 2372
rect 33836 2360 33842 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 33836 2332 35173 2360
rect 33836 2320 33842 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 35250 2320 35256 2372
rect 35308 2360 35314 2372
rect 37737 2363 37795 2369
rect 37737 2360 37749 2363
rect 35308 2332 37749 2360
rect 35308 2320 35314 2332
rect 37737 2329 37749 2332
rect 37783 2329 37795 2363
rect 38654 2360 38660 2372
rect 38615 2332 38660 2360
rect 37737 2323 37795 2329
rect 38654 2320 38660 2332
rect 38712 2320 38718 2372
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 40129 2363 40187 2369
rect 40129 2360 40141 2363
rect 39264 2332 40141 2360
rect 39264 2320 39270 2332
rect 40129 2329 40141 2332
rect 40175 2329 40187 2363
rect 40129 2323 40187 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 41230 2320 41236 2372
rect 41288 2360 41294 2372
rect 42720 2360 42748 2400
rect 43438 2360 43444 2372
rect 41288 2332 42748 2360
rect 43399 2332 43444 2360
rect 41288 2320 41294 2332
rect 43438 2320 43444 2332
rect 43496 2320 43502 2372
rect 43548 2360 43576 2400
rect 44177 2397 44189 2431
rect 44223 2397 44235 2431
rect 44177 2391 44235 2397
rect 46382 2388 46388 2440
rect 46440 2428 46446 2440
rect 47857 2431 47915 2437
rect 47857 2428 47869 2431
rect 46440 2400 47869 2428
rect 46440 2388 46446 2400
rect 47857 2397 47869 2400
rect 47903 2397 47915 2431
rect 50341 2431 50399 2437
rect 50341 2428 50353 2431
rect 47857 2391 47915 2397
rect 47964 2400 50353 2428
rect 44361 2363 44419 2369
rect 44361 2360 44373 2363
rect 43548 2332 44373 2360
rect 44361 2329 44373 2332
rect 44407 2329 44419 2363
rect 44361 2323 44419 2329
rect 45554 2320 45560 2372
rect 45612 2360 45618 2372
rect 45741 2363 45799 2369
rect 45741 2360 45753 2363
rect 45612 2332 45753 2360
rect 45612 2320 45618 2332
rect 45741 2329 45753 2332
rect 45787 2329 45799 2363
rect 45741 2323 45799 2329
rect 45830 2320 45836 2372
rect 45888 2360 45894 2372
rect 46661 2363 46719 2369
rect 46661 2360 46673 2363
rect 45888 2332 46673 2360
rect 45888 2320 45894 2332
rect 46661 2329 46673 2332
rect 46707 2329 46719 2363
rect 46661 2323 46719 2329
rect 47210 2320 47216 2372
rect 47268 2360 47274 2372
rect 47964 2360 47992 2400
rect 50341 2397 50353 2400
rect 50387 2397 50399 2431
rect 51905 2431 51963 2437
rect 51905 2428 51917 2431
rect 50341 2391 50399 2397
rect 50632 2400 51917 2428
rect 47268 2332 47992 2360
rect 47268 2320 47274 2332
rect 48038 2320 48044 2372
rect 48096 2360 48102 2372
rect 48777 2363 48835 2369
rect 48777 2360 48789 2363
rect 48096 2332 48789 2360
rect 48096 2320 48102 2332
rect 48777 2329 48789 2332
rect 48823 2329 48835 2363
rect 48777 2323 48835 2329
rect 49970 2320 49976 2372
rect 50028 2360 50034 2372
rect 50632 2360 50660 2400
rect 51905 2397 51917 2400
rect 51951 2397 51963 2431
rect 51905 2391 51963 2397
rect 54662 2388 54668 2440
rect 54720 2428 54726 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 54720 2400 55505 2428
rect 54720 2388 54726 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 56410 2428 56416 2440
rect 56371 2400 56416 2428
rect 55493 2391 55551 2397
rect 56410 2388 56416 2400
rect 56468 2388 56474 2440
rect 57882 2388 57888 2440
rect 57940 2428 57946 2440
rect 58161 2431 58219 2437
rect 58161 2428 58173 2431
rect 57940 2400 58173 2428
rect 57940 2388 57946 2400
rect 58161 2397 58173 2400
rect 58207 2397 58219 2431
rect 58161 2391 58219 2397
rect 51169 2363 51227 2369
rect 51169 2360 51181 2363
rect 50028 2332 50660 2360
rect 51092 2332 51181 2360
rect 50028 2320 50034 2332
rect 32088 2264 33548 2292
rect 32088 2252 32094 2264
rect 33594 2252 33600 2304
rect 33652 2292 33658 2304
rect 36725 2295 36783 2301
rect 36725 2292 36737 2295
rect 33652 2264 36737 2292
rect 33652 2252 33658 2264
rect 36725 2261 36737 2264
rect 36771 2261 36783 2295
rect 43530 2292 43536 2304
rect 43491 2264 43536 2292
rect 36725 2255 36783 2261
rect 43530 2252 43536 2264
rect 43588 2252 43594 2304
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 51092 2292 51120 2332
rect 51169 2329 51181 2332
rect 51215 2329 51227 2363
rect 51169 2323 51227 2329
rect 52178 2320 52184 2372
rect 52236 2360 52242 2372
rect 53009 2363 53067 2369
rect 53009 2360 53021 2363
rect 52236 2332 53021 2360
rect 52236 2320 52242 2332
rect 53009 2329 53021 2332
rect 53055 2329 53067 2363
rect 53009 2323 53067 2329
rect 53282 2320 53288 2372
rect 53340 2360 53346 2372
rect 53929 2363 53987 2369
rect 53929 2360 53941 2363
rect 53340 2332 53941 2360
rect 53340 2320 53346 2332
rect 53929 2329 53941 2332
rect 53975 2329 53987 2363
rect 53929 2323 53987 2329
rect 56689 2363 56747 2369
rect 56689 2329 56701 2363
rect 56735 2329 56747 2363
rect 56689 2323 56747 2329
rect 51258 2292 51264 2304
rect 48372 2264 51120 2292
rect 51219 2264 51264 2292
rect 48372 2252 48378 2264
rect 51258 2252 51264 2264
rect 51316 2252 51322 2304
rect 53098 2292 53104 2304
rect 53059 2264 53104 2292
rect 53098 2252 53104 2264
rect 53156 2252 53162 2304
rect 55490 2252 55496 2304
rect 55548 2292 55554 2304
rect 56704 2292 56732 2323
rect 55548 2264 56732 2292
rect 55548 2252 55554 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 9306 2048 9312 2100
rect 9364 2088 9370 2100
rect 17218 2088 17224 2100
rect 9364 2060 17224 2088
rect 9364 2048 9370 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 18690 2048 18696 2100
rect 18748 2088 18754 2100
rect 28994 2088 29000 2100
rect 18748 2060 29000 2088
rect 18748 2048 18754 2060
rect 28994 2048 29000 2060
rect 29052 2048 29058 2100
rect 29362 2048 29368 2100
rect 29420 2088 29426 2100
rect 29420 2060 31754 2088
rect 29420 2048 29426 2060
rect 5810 1980 5816 2032
rect 5868 2020 5874 2032
rect 13262 2020 13268 2032
rect 5868 1992 13268 2020
rect 5868 1980 5874 1992
rect 13262 1980 13268 1992
rect 13320 1980 13326 2032
rect 15562 2020 15568 2032
rect 13464 1992 15568 2020
rect 5074 1912 5080 1964
rect 5132 1952 5138 1964
rect 11882 1952 11888 1964
rect 5132 1924 11888 1952
rect 5132 1912 5138 1924
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 13464 1952 13492 1992
rect 15562 1980 15568 1992
rect 15620 1980 15626 2032
rect 17770 1980 17776 2032
rect 17828 2020 17834 2032
rect 28442 2020 28448 2032
rect 17828 1992 28448 2020
rect 17828 1980 17834 1992
rect 28442 1980 28448 1992
rect 28500 1980 28506 2032
rect 31726 2020 31754 2060
rect 33410 2048 33416 2100
rect 33468 2088 33474 2100
rect 35250 2088 35256 2100
rect 33468 2060 35256 2088
rect 33468 2048 33474 2060
rect 35250 2048 35256 2060
rect 35308 2048 35314 2100
rect 36722 2048 36728 2100
rect 36780 2088 36786 2100
rect 43438 2088 43444 2100
rect 36780 2060 43444 2088
rect 36780 2048 36786 2060
rect 43438 2048 43444 2060
rect 43496 2048 43502 2100
rect 43898 2048 43904 2100
rect 43956 2088 43962 2100
rect 45738 2088 45744 2100
rect 43956 2060 45744 2088
rect 43956 2048 43962 2060
rect 45738 2048 45744 2060
rect 45796 2048 45802 2100
rect 34146 2020 34152 2032
rect 31726 1992 34152 2020
rect 34146 1980 34152 1992
rect 34204 1980 34210 2032
rect 34238 1980 34244 2032
rect 34296 2020 34302 2032
rect 38654 2020 38660 2032
rect 34296 1992 38660 2020
rect 34296 1980 34302 1992
rect 38654 1980 38660 1992
rect 38712 1980 38718 2032
rect 12400 1924 13492 1952
rect 12400 1912 12406 1924
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 22922 1952 22928 1964
rect 13596 1924 22928 1952
rect 13596 1912 13602 1924
rect 22922 1912 22928 1924
rect 22980 1912 22986 1964
rect 31570 1912 31576 1964
rect 31628 1952 31634 1964
rect 51258 1952 51264 1964
rect 31628 1924 51264 1952
rect 31628 1912 31634 1924
rect 51258 1912 51264 1924
rect 51316 1912 51322 1964
rect 7006 1844 7012 1896
rect 7064 1884 7070 1896
rect 12802 1884 12808 1896
rect 7064 1856 12808 1884
rect 7064 1844 7070 1856
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 18414 1844 18420 1896
rect 18472 1884 18478 1896
rect 19886 1884 19892 1896
rect 18472 1856 19892 1884
rect 18472 1844 18478 1856
rect 19886 1844 19892 1856
rect 19944 1844 19950 1896
rect 20254 1844 20260 1896
rect 20312 1884 20318 1896
rect 29270 1884 29276 1896
rect 20312 1856 29276 1884
rect 20312 1844 20318 1856
rect 29270 1844 29276 1856
rect 29328 1844 29334 1896
rect 29638 1844 29644 1896
rect 29696 1884 29702 1896
rect 53098 1884 53104 1896
rect 29696 1856 53104 1884
rect 29696 1844 29702 1856
rect 53098 1844 53104 1856
rect 53156 1844 53162 1896
rect 6730 1776 6736 1828
rect 6788 1816 6794 1828
rect 13538 1816 13544 1828
rect 6788 1788 13544 1816
rect 6788 1776 6794 1788
rect 13538 1776 13544 1788
rect 13596 1776 13602 1828
rect 15930 1776 15936 1828
rect 15988 1816 15994 1828
rect 24578 1816 24584 1828
rect 15988 1788 24584 1816
rect 15988 1776 15994 1788
rect 24578 1776 24584 1788
rect 24636 1776 24642 1828
rect 26510 1776 26516 1828
rect 26568 1816 26574 1828
rect 56410 1816 56416 1828
rect 26568 1788 56416 1816
rect 26568 1776 26574 1788
rect 56410 1776 56416 1788
rect 56468 1776 56474 1828
rect 4890 1708 4896 1760
rect 4948 1748 4954 1760
rect 11330 1748 11336 1760
rect 4948 1720 11336 1748
rect 4948 1708 4954 1720
rect 11330 1708 11336 1720
rect 11388 1708 11394 1760
rect 12710 1708 12716 1760
rect 12768 1748 12774 1760
rect 20438 1748 20444 1760
rect 12768 1720 20444 1748
rect 12768 1708 12774 1720
rect 20438 1708 20444 1720
rect 20496 1708 20502 1760
rect 20622 1708 20628 1760
rect 20680 1748 20686 1760
rect 23474 1748 23480 1760
rect 20680 1720 23480 1748
rect 20680 1708 20686 1720
rect 23474 1708 23480 1720
rect 23532 1708 23538 1760
rect 24210 1708 24216 1760
rect 24268 1748 24274 1760
rect 53466 1748 53472 1760
rect 24268 1720 53472 1748
rect 24268 1708 24274 1720
rect 53466 1708 53472 1720
rect 53524 1708 53530 1760
rect 11422 1680 11428 1692
rect 6886 1652 11428 1680
rect 5166 1572 5172 1624
rect 5224 1612 5230 1624
rect 6886 1612 6914 1652
rect 11422 1640 11428 1652
rect 11480 1640 11486 1692
rect 16114 1640 16120 1692
rect 16172 1680 16178 1692
rect 28166 1680 28172 1692
rect 16172 1652 28172 1680
rect 16172 1640 16178 1652
rect 28166 1640 28172 1652
rect 28224 1640 28230 1692
rect 39482 1640 39488 1692
rect 39540 1680 39546 1692
rect 46014 1680 46020 1692
rect 39540 1652 46020 1680
rect 39540 1640 39546 1652
rect 46014 1640 46020 1652
rect 46072 1640 46078 1692
rect 5224 1584 6914 1612
rect 5224 1572 5230 1584
rect 10962 1572 10968 1624
rect 11020 1612 11026 1624
rect 17954 1612 17960 1624
rect 11020 1584 17960 1612
rect 11020 1572 11026 1584
rect 17954 1572 17960 1584
rect 18012 1572 18018 1624
rect 19242 1572 19248 1624
rect 19300 1612 19306 1624
rect 27890 1612 27896 1624
rect 19300 1584 27896 1612
rect 19300 1572 19306 1584
rect 27890 1572 27896 1584
rect 27948 1572 27954 1624
rect 1578 1504 1584 1556
rect 1636 1544 1642 1556
rect 15102 1544 15108 1556
rect 1636 1516 15108 1544
rect 1636 1504 1642 1516
rect 15102 1504 15108 1516
rect 15160 1504 15166 1556
rect 15838 1504 15844 1556
rect 15896 1544 15902 1556
rect 28258 1544 28264 1556
rect 15896 1516 28264 1544
rect 15896 1504 15902 1516
rect 28258 1504 28264 1516
rect 28316 1504 28322 1556
rect 4706 1436 4712 1488
rect 4764 1476 4770 1488
rect 8294 1476 8300 1488
rect 4764 1448 8300 1476
rect 4764 1436 4770 1448
rect 8294 1436 8300 1448
rect 8352 1436 8358 1488
rect 10594 1436 10600 1488
rect 10652 1476 10658 1488
rect 17402 1476 17408 1488
rect 10652 1448 17408 1476
rect 10652 1436 10658 1448
rect 17402 1436 17408 1448
rect 17460 1436 17466 1488
rect 20346 1436 20352 1488
rect 20404 1476 20410 1488
rect 23198 1476 23204 1488
rect 20404 1448 23204 1476
rect 20404 1436 20410 1448
rect 23198 1436 23204 1448
rect 23256 1436 23262 1488
rect 40770 1476 40776 1488
rect 31726 1448 40776 1476
rect 3326 1368 3332 1420
rect 3384 1408 3390 1420
rect 11146 1408 11152 1420
rect 3384 1380 11152 1408
rect 3384 1368 3390 1380
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 13354 1368 13360 1420
rect 13412 1408 13418 1420
rect 19242 1408 19248 1420
rect 13412 1380 19248 1408
rect 13412 1368 13418 1380
rect 19242 1368 19248 1380
rect 19300 1368 19306 1420
rect 20070 1368 20076 1420
rect 20128 1408 20134 1420
rect 20990 1408 20996 1420
rect 20128 1380 20996 1408
rect 20128 1368 20134 1380
rect 20990 1368 20996 1380
rect 21048 1368 21054 1420
rect 22278 1368 22284 1420
rect 22336 1408 22342 1420
rect 31726 1408 31754 1448
rect 40770 1436 40776 1448
rect 40828 1436 40834 1488
rect 43346 1436 43352 1488
rect 43404 1476 43410 1488
rect 47118 1476 47124 1488
rect 43404 1448 47124 1476
rect 43404 1436 43410 1448
rect 47118 1436 47124 1448
rect 47176 1436 47182 1488
rect 22336 1380 31754 1408
rect 22336 1368 22342 1380
rect 32582 1368 32588 1420
rect 32640 1408 32646 1420
rect 33778 1408 33784 1420
rect 32640 1380 33784 1408
rect 32640 1368 32646 1380
rect 33778 1368 33784 1380
rect 33836 1368 33842 1420
rect 37274 1368 37280 1420
rect 37332 1408 37338 1420
rect 38562 1408 38568 1420
rect 37332 1380 38568 1408
rect 37332 1368 37338 1380
rect 38562 1368 38568 1380
rect 38620 1368 38626 1420
rect 16942 1300 16948 1352
rect 17000 1340 17006 1352
rect 40954 1340 40960 1352
rect 17000 1312 40960 1340
rect 17000 1300 17006 1312
rect 40954 1300 40960 1312
rect 41012 1300 41018 1352
rect 13446 1232 13452 1284
rect 13504 1272 13510 1284
rect 23566 1272 23572 1284
rect 13504 1244 23572 1272
rect 13504 1232 13510 1244
rect 23566 1232 23572 1244
rect 23624 1232 23630 1284
rect 10686 1164 10692 1216
rect 10744 1204 10750 1216
rect 33502 1204 33508 1216
rect 10744 1176 33508 1204
rect 10744 1164 10750 1176
rect 33502 1164 33508 1176
rect 33560 1164 33566 1216
rect 42518 1164 42524 1216
rect 42576 1204 42582 1216
rect 44542 1204 44548 1216
rect 42576 1176 44548 1204
rect 42576 1164 42582 1176
rect 44542 1164 44548 1176
rect 44600 1164 44606 1216
rect 3602 1096 3608 1148
rect 3660 1136 3666 1148
rect 7190 1136 7196 1148
rect 3660 1108 7196 1136
rect 3660 1096 3666 1108
rect 7190 1096 7196 1108
rect 7248 1096 7254 1148
rect 8662 1096 8668 1148
rect 8720 1136 8726 1148
rect 29178 1136 29184 1148
rect 8720 1108 29184 1136
rect 8720 1096 8726 1108
rect 29178 1096 29184 1108
rect 29236 1096 29242 1148
rect 4982 1028 4988 1080
rect 5040 1068 5046 1080
rect 24762 1068 24768 1080
rect 5040 1040 24768 1068
rect 5040 1028 5046 1040
rect 24762 1028 24768 1040
rect 24820 1028 24826 1080
rect 6454 960 6460 1012
rect 6512 1000 6518 1012
rect 24394 1000 24400 1012
rect 6512 972 24400 1000
rect 6512 960 6518 972
rect 24394 960 24400 972
rect 24452 960 24458 1012
rect 5350 892 5356 944
rect 5408 932 5414 944
rect 23382 932 23388 944
rect 5408 904 23388 932
rect 5408 892 5414 904
rect 23382 892 23388 904
rect 23440 892 23446 944
rect 3142 824 3148 876
rect 3200 864 3206 876
rect 22738 864 22744 876
rect 3200 836 22744 864
rect 3200 824 3206 836
rect 22738 824 22744 836
rect 22796 824 22802 876
rect 6178 756 6184 808
rect 6236 796 6242 808
rect 24486 796 24492 808
rect 6236 768 24492 796
rect 6236 756 6242 768
rect 24486 756 24492 768
rect 24544 756 24550 808
rect 4798 688 4804 740
rect 4856 728 4862 740
rect 28626 728 28632 740
rect 4856 700 28632 728
rect 4856 688 4862 700
rect 28626 688 28632 700
rect 28684 688 28690 740
rect 2314 620 2320 672
rect 2372 660 2378 672
rect 21634 660 21640 672
rect 2372 632 21640 660
rect 2372 620 2378 632
rect 21634 620 21640 632
rect 21692 620 21698 672
rect 18966 552 18972 604
rect 19024 592 19030 604
rect 25774 592 25780 604
rect 19024 564 25780 592
rect 19024 552 19030 564
rect 25774 552 25780 564
rect 25832 552 25838 604
rect 18874 484 18880 536
rect 18932 524 18938 536
rect 24210 524 24216 536
rect 18932 496 24216 524
rect 18932 484 18938 496
rect 24210 484 24216 496
rect 24268 484 24274 536
<< via1 >>
rect 41236 61684 41288 61736
rect 51448 61684 51500 61736
rect 24952 61616 25004 61668
rect 40316 61616 40368 61668
rect 40408 61616 40460 61668
rect 42708 61616 42760 61668
rect 28356 61548 28408 61600
rect 40684 61548 40736 61600
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 7656 61344 7708 61396
rect 15292 61344 15344 61396
rect 22836 61344 22888 61396
rect 40408 61344 40460 61396
rect 40684 61344 40736 61396
rect 51448 61387 51500 61396
rect 51448 61353 51457 61387
rect 51457 61353 51491 61387
rect 51491 61353 51500 61387
rect 51448 61344 51500 61353
rect 6276 61276 6328 61328
rect 40316 61276 40368 61328
rect 46756 61276 46808 61328
rect 48964 61276 49016 61328
rect 17408 61208 17460 61260
rect 20628 61208 20680 61260
rect 28264 61208 28316 61260
rect 39580 61208 39632 61260
rect 41144 61208 41196 61260
rect 1676 61183 1728 61192
rect 1676 61149 1685 61183
rect 1685 61149 1719 61183
rect 1719 61149 1728 61183
rect 1676 61140 1728 61149
rect 2780 61183 2832 61192
rect 2780 61149 2789 61183
rect 2789 61149 2823 61183
rect 2823 61149 2832 61183
rect 4712 61183 4764 61192
rect 2780 61140 2832 61149
rect 4712 61149 4721 61183
rect 4721 61149 4755 61183
rect 4755 61149 4764 61183
rect 4712 61140 4764 61149
rect 6000 61140 6052 61192
rect 6644 61183 6696 61192
rect 6644 61149 6653 61183
rect 6653 61149 6687 61183
rect 6687 61149 6696 61183
rect 6644 61140 6696 61149
rect 7564 61183 7616 61192
rect 7564 61149 7573 61183
rect 7573 61149 7607 61183
rect 7607 61149 7616 61183
rect 7564 61140 7616 61149
rect 9220 61183 9272 61192
rect 9220 61149 9229 61183
rect 9229 61149 9263 61183
rect 9263 61149 9272 61183
rect 9220 61140 9272 61149
rect 10232 61183 10284 61192
rect 10232 61149 10241 61183
rect 10241 61149 10275 61183
rect 10275 61149 10284 61183
rect 10232 61140 10284 61149
rect 11152 61140 11204 61192
rect 12072 61183 12124 61192
rect 12072 61149 12081 61183
rect 12081 61149 12115 61183
rect 12115 61149 12124 61183
rect 12072 61140 12124 61149
rect 12808 61183 12860 61192
rect 12808 61149 12817 61183
rect 12817 61149 12851 61183
rect 12851 61149 12860 61183
rect 12808 61140 12860 61149
rect 14924 61183 14976 61192
rect 14924 61149 14933 61183
rect 14933 61149 14967 61183
rect 14967 61149 14976 61183
rect 14924 61140 14976 61149
rect 16120 61183 16172 61192
rect 16120 61149 16129 61183
rect 16129 61149 16163 61183
rect 16163 61149 16172 61183
rect 16120 61140 16172 61149
rect 17132 61183 17184 61192
rect 17132 61149 17141 61183
rect 17141 61149 17175 61183
rect 17175 61149 17184 61183
rect 17132 61140 17184 61149
rect 17960 61183 18012 61192
rect 17960 61149 17969 61183
rect 17969 61149 18003 61183
rect 18003 61149 18012 61183
rect 17960 61140 18012 61149
rect 18696 61183 18748 61192
rect 18696 61149 18705 61183
rect 18705 61149 18739 61183
rect 18739 61149 18748 61183
rect 18696 61140 18748 61149
rect 19800 61183 19852 61192
rect 19800 61149 19809 61183
rect 19809 61149 19843 61183
rect 19843 61149 19852 61183
rect 19800 61140 19852 61149
rect 20720 61140 20772 61192
rect 21272 61183 21324 61192
rect 21272 61149 21281 61183
rect 21281 61149 21315 61183
rect 21315 61149 21324 61183
rect 21272 61140 21324 61149
rect 22376 61183 22428 61192
rect 22376 61149 22385 61183
rect 22385 61149 22419 61183
rect 22419 61149 22428 61183
rect 22376 61140 22428 61149
rect 23664 61140 23716 61192
rect 25136 61140 25188 61192
rect 25872 61140 25924 61192
rect 26608 61140 26660 61192
rect 28080 61140 28132 61192
rect 29828 61183 29880 61192
rect 29828 61149 29837 61183
rect 29837 61149 29871 61183
rect 29871 61149 29880 61183
rect 29828 61140 29880 61149
rect 31208 61183 31260 61192
rect 31208 61149 31217 61183
rect 31217 61149 31251 61183
rect 31251 61149 31260 61183
rect 31208 61140 31260 61149
rect 31760 61140 31812 61192
rect 32496 61140 32548 61192
rect 33508 61140 33560 61192
rect 34244 61140 34296 61192
rect 35072 61140 35124 61192
rect 5540 61072 5592 61124
rect 7840 61115 7892 61124
rect 5724 61047 5776 61056
rect 5724 61013 5733 61047
rect 5733 61013 5767 61047
rect 5767 61013 5776 61047
rect 5724 61004 5776 61013
rect 7840 61081 7849 61115
rect 7849 61081 7883 61115
rect 7883 61081 7892 61115
rect 7840 61072 7892 61081
rect 10508 61072 10560 61124
rect 15200 61115 15252 61124
rect 15200 61081 15209 61115
rect 15209 61081 15243 61115
rect 15243 61081 15252 61115
rect 15200 61072 15252 61081
rect 17500 61072 17552 61124
rect 19984 61115 20036 61124
rect 19984 61081 19993 61115
rect 19993 61081 20027 61115
rect 20027 61081 20036 61115
rect 19984 61072 20036 61081
rect 9312 61047 9364 61056
rect 9312 61013 9321 61047
rect 9321 61013 9355 61047
rect 9355 61013 9364 61047
rect 9312 61004 9364 61013
rect 10324 61047 10376 61056
rect 10324 61013 10333 61047
rect 10333 61013 10367 61047
rect 10367 61013 10376 61047
rect 10324 61004 10376 61013
rect 12164 61047 12216 61056
rect 12164 61013 12173 61047
rect 12173 61013 12207 61047
rect 12207 61013 12216 61047
rect 12164 61004 12216 61013
rect 12900 61047 12952 61056
rect 12900 61013 12909 61047
rect 12909 61013 12943 61047
rect 12943 61013 12952 61047
rect 12900 61004 12952 61013
rect 17316 61047 17368 61056
rect 17316 61013 17325 61047
rect 17325 61013 17359 61047
rect 17359 61013 17368 61047
rect 17316 61004 17368 61013
rect 18604 61004 18656 61056
rect 22284 61072 22336 61124
rect 26884 61072 26936 61124
rect 28448 61115 28500 61124
rect 28448 61081 28457 61115
rect 28457 61081 28491 61115
rect 28491 61081 28500 61115
rect 28448 61072 28500 61081
rect 31576 61115 31628 61124
rect 31576 61081 31585 61115
rect 31585 61081 31619 61115
rect 31619 61081 31628 61115
rect 31576 61072 31628 61081
rect 34704 61072 34756 61124
rect 35900 61140 35952 61192
rect 36912 61140 36964 61192
rect 37648 61140 37700 61192
rect 38660 61140 38712 61192
rect 39488 61140 39540 61192
rect 40132 61140 40184 61192
rect 40960 61140 41012 61192
rect 42064 61140 42116 61192
rect 42800 61140 42852 61192
rect 43628 61140 43680 61192
rect 44548 61140 44600 61192
rect 45560 61140 45612 61192
rect 46112 61140 46164 61192
rect 47216 61140 47268 61192
rect 48320 61140 48372 61192
rect 48688 61140 48740 61192
rect 49700 61140 49752 61192
rect 51080 61140 51132 61192
rect 51632 61140 51684 61192
rect 53196 61183 53248 61192
rect 53196 61149 53205 61183
rect 53205 61149 53239 61183
rect 53239 61149 53248 61183
rect 53196 61140 53248 61149
rect 54116 61183 54168 61192
rect 54116 61149 54125 61183
rect 54125 61149 54159 61183
rect 54159 61149 54168 61183
rect 54116 61140 54168 61149
rect 55496 61183 55548 61192
rect 55496 61149 55505 61183
rect 55505 61149 55539 61183
rect 55539 61149 55548 61183
rect 55496 61140 55548 61149
rect 56048 61140 56100 61192
rect 57520 61140 57572 61192
rect 39764 61072 39816 61124
rect 42892 61115 42944 61124
rect 21456 61004 21508 61056
rect 23756 61004 23808 61056
rect 27344 61047 27396 61056
rect 27344 61013 27353 61047
rect 27353 61013 27387 61047
rect 27387 61013 27396 61047
rect 27344 61004 27396 61013
rect 29920 61047 29972 61056
rect 29920 61013 29929 61047
rect 29929 61013 29963 61047
rect 29963 61013 29972 61047
rect 29920 61004 29972 61013
rect 33508 61004 33560 61056
rect 34244 61004 34296 61056
rect 35348 61004 35400 61056
rect 36084 61004 36136 61056
rect 37280 61004 37332 61056
rect 39120 61047 39172 61056
rect 39120 61013 39129 61047
rect 39129 61013 39163 61047
rect 39163 61013 39172 61047
rect 39120 61004 39172 61013
rect 40316 61004 40368 61056
rect 41696 61047 41748 61056
rect 41696 61013 41705 61047
rect 41705 61013 41739 61047
rect 41739 61013 41748 61047
rect 41696 61004 41748 61013
rect 42892 61081 42901 61115
rect 42901 61081 42935 61115
rect 42935 61081 42944 61115
rect 42892 61072 42944 61081
rect 46940 61072 46992 61124
rect 45376 61047 45428 61056
rect 45376 61013 45385 61047
rect 45385 61013 45419 61047
rect 45419 61013 45428 61047
rect 45376 61004 45428 61013
rect 46112 61047 46164 61056
rect 46112 61013 46121 61047
rect 46121 61013 46155 61047
rect 46155 61013 46164 61047
rect 46112 61004 46164 61013
rect 46848 61047 46900 61056
rect 46848 61013 46857 61047
rect 46857 61013 46891 61047
rect 46891 61013 46900 61047
rect 46848 61004 46900 61013
rect 47584 61004 47636 61056
rect 50068 61004 50120 61056
rect 51816 61004 51868 61056
rect 58348 61115 58400 61124
rect 58348 61081 58357 61115
rect 58357 61081 58391 61115
rect 58391 61081 58400 61115
rect 58348 61072 58400 61081
rect 54300 61047 54352 61056
rect 54300 61013 54309 61047
rect 54309 61013 54343 61047
rect 54343 61013 54352 61047
rect 54300 61004 54352 61013
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 10324 60800 10376 60852
rect 22192 60800 22244 60852
rect 27160 60800 27212 60852
rect 46848 60800 46900 60852
rect 3976 60775 4028 60784
rect 3976 60741 3985 60775
rect 3985 60741 4019 60775
rect 4019 60741 4028 60775
rect 3976 60732 4028 60741
rect 5448 60775 5500 60784
rect 5448 60741 5457 60775
rect 5457 60741 5491 60775
rect 5491 60741 5500 60775
rect 5448 60732 5500 60741
rect 8300 60732 8352 60784
rect 9864 60775 9916 60784
rect 9864 60741 9873 60775
rect 9873 60741 9907 60775
rect 9907 60741 9916 60775
rect 9864 60732 9916 60741
rect 13544 60775 13596 60784
rect 13544 60741 13553 60775
rect 13553 60741 13587 60775
rect 13587 60741 13596 60775
rect 13544 60732 13596 60741
rect 14280 60775 14332 60784
rect 14280 60741 14289 60775
rect 14289 60741 14323 60775
rect 14323 60741 14332 60775
rect 14280 60732 14332 60741
rect 15752 60775 15804 60784
rect 15752 60741 15761 60775
rect 15761 60741 15795 60775
rect 15795 60741 15804 60775
rect 15752 60732 15804 60741
rect 19340 60732 19392 60784
rect 23296 60775 23348 60784
rect 23296 60741 23305 60775
rect 23305 60741 23339 60775
rect 23339 60741 23348 60775
rect 23296 60732 23348 60741
rect 24584 60775 24636 60784
rect 24584 60741 24593 60775
rect 24593 60741 24627 60775
rect 24627 60741 24636 60775
rect 24584 60732 24636 60741
rect 27528 60775 27580 60784
rect 27528 60741 27537 60775
rect 27537 60741 27571 60775
rect 27571 60741 27580 60775
rect 27528 60732 27580 60741
rect 29000 60775 29052 60784
rect 29000 60741 29009 60775
rect 29009 60741 29043 60775
rect 29043 60741 29052 60775
rect 29000 60732 29052 60741
rect 30380 60732 30432 60784
rect 36360 60775 36412 60784
rect 36360 60741 36369 60775
rect 36369 60741 36403 60775
rect 36403 60741 36412 60775
rect 36360 60732 36412 60741
rect 41420 60732 41472 60784
rect 46664 60775 46716 60784
rect 46664 60741 46673 60775
rect 46673 60741 46707 60775
rect 46707 60741 46716 60775
rect 46664 60732 46716 60741
rect 50160 60732 50212 60784
rect 52460 60732 52512 60784
rect 1584 60707 1636 60716
rect 1584 60673 1593 60707
rect 1593 60673 1627 60707
rect 1627 60673 1636 60707
rect 1584 60664 1636 60673
rect 3148 60707 3200 60716
rect 3148 60673 3157 60707
rect 3157 60673 3191 60707
rect 3191 60673 3200 60707
rect 3148 60664 3200 60673
rect 21272 60664 21324 60716
rect 22100 60707 22152 60716
rect 22100 60673 22109 60707
rect 22109 60673 22143 60707
rect 22143 60673 22152 60707
rect 22100 60664 22152 60673
rect 24676 60664 24728 60716
rect 35072 60664 35124 60716
rect 4804 60596 4856 60648
rect 13636 60596 13688 60648
rect 22468 60596 22520 60648
rect 22652 60639 22704 60648
rect 22652 60605 22661 60639
rect 22661 60605 22695 60639
rect 22695 60605 22704 60639
rect 41604 60664 41656 60716
rect 54668 60707 54720 60716
rect 54668 60673 54677 60707
rect 54677 60673 54711 60707
rect 54711 60673 54720 60707
rect 54668 60664 54720 60673
rect 55404 60707 55456 60716
rect 55404 60673 55413 60707
rect 55413 60673 55447 60707
rect 55447 60673 55456 60707
rect 55404 60664 55456 60673
rect 56140 60707 56192 60716
rect 56140 60673 56149 60707
rect 56149 60673 56183 60707
rect 56183 60673 56192 60707
rect 56140 60664 56192 60673
rect 56876 60707 56928 60716
rect 56876 60673 56885 60707
rect 56885 60673 56919 60707
rect 56919 60673 56928 60707
rect 56876 60664 56928 60673
rect 58072 60707 58124 60716
rect 58072 60673 58081 60707
rect 58081 60673 58115 60707
rect 58115 60673 58124 60707
rect 58072 60664 58124 60673
rect 22652 60596 22704 60605
rect 36636 60596 36688 60648
rect 46940 60596 46992 60648
rect 4620 60528 4672 60580
rect 3332 60503 3384 60512
rect 3332 60469 3341 60503
rect 3341 60469 3375 60503
rect 3375 60469 3384 60503
rect 3332 60460 3384 60469
rect 9956 60503 10008 60512
rect 9956 60469 9965 60503
rect 9965 60469 9999 60503
rect 9999 60469 10008 60503
rect 9956 60460 10008 60469
rect 15844 60503 15896 60512
rect 15844 60469 15853 60503
rect 15853 60469 15887 60503
rect 15887 60469 15896 60503
rect 15844 60460 15896 60469
rect 20352 60528 20404 60580
rect 24492 60528 24544 60580
rect 25228 60528 25280 60580
rect 22836 60460 22888 60512
rect 24400 60460 24452 60512
rect 28080 60460 28132 60512
rect 28172 60460 28224 60512
rect 28356 60460 28408 60512
rect 29092 60503 29144 60512
rect 29092 60469 29101 60503
rect 29101 60469 29135 60503
rect 29135 60469 29144 60503
rect 29092 60460 29144 60469
rect 35624 60460 35676 60512
rect 35716 60460 35768 60512
rect 41972 60460 42024 60512
rect 44180 60460 44232 60512
rect 50436 60503 50488 60512
rect 50436 60469 50445 60503
rect 50445 60469 50479 60503
rect 50479 60469 50488 60503
rect 50436 60460 50488 60469
rect 53104 60503 53156 60512
rect 53104 60469 53113 60503
rect 53113 60469 53147 60503
rect 53147 60469 53156 60503
rect 53104 60460 53156 60469
rect 54852 60503 54904 60512
rect 54852 60469 54861 60503
rect 54861 60469 54895 60503
rect 54895 60469 54904 60503
rect 54852 60460 54904 60469
rect 55588 60503 55640 60512
rect 55588 60469 55597 60503
rect 55597 60469 55631 60503
rect 55631 60469 55640 60503
rect 55588 60460 55640 60469
rect 56324 60503 56376 60512
rect 56324 60469 56333 60503
rect 56333 60469 56367 60503
rect 56367 60469 56376 60503
rect 56324 60460 56376 60469
rect 57060 60503 57112 60512
rect 57060 60469 57069 60503
rect 57069 60469 57103 60503
rect 57103 60469 57112 60503
rect 57060 60460 57112 60469
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 9956 60256 10008 60308
rect 19248 60256 19300 60308
rect 6644 60188 6696 60240
rect 13636 60188 13688 60240
rect 15844 60120 15896 60172
rect 2596 60095 2648 60104
rect 2596 60061 2605 60095
rect 2605 60061 2639 60095
rect 2639 60061 2648 60095
rect 2596 60052 2648 60061
rect 6000 60095 6052 60104
rect 6000 60061 6009 60095
rect 6009 60061 6043 60095
rect 6043 60061 6052 60095
rect 6000 60052 6052 60061
rect 6276 60095 6328 60104
rect 6276 60061 6285 60095
rect 6285 60061 6319 60095
rect 6319 60061 6328 60095
rect 6276 60052 6328 60061
rect 7012 60052 7064 60104
rect 1676 60027 1728 60036
rect 1676 59993 1685 60027
rect 1685 59993 1719 60027
rect 1719 59993 1728 60027
rect 1676 59984 1728 59993
rect 2044 60027 2096 60036
rect 2044 59993 2053 60027
rect 2053 59993 2087 60027
rect 2087 59993 2096 60027
rect 2044 59984 2096 59993
rect 3884 59984 3936 60036
rect 6736 59984 6788 60036
rect 19432 60052 19484 60104
rect 19984 60095 20036 60104
rect 19984 60061 19993 60095
rect 19993 60061 20027 60095
rect 20027 60061 20036 60095
rect 19984 60052 20036 60061
rect 20536 60231 20588 60240
rect 20536 60197 20545 60231
rect 20545 60197 20579 60231
rect 20579 60197 20588 60231
rect 20536 60188 20588 60197
rect 22652 60188 22704 60240
rect 22928 60256 22980 60308
rect 25964 60256 26016 60308
rect 26792 60256 26844 60308
rect 29736 60256 29788 60308
rect 30012 60256 30064 60308
rect 58256 60256 58308 60308
rect 25872 60188 25924 60240
rect 26056 60188 26108 60240
rect 21272 60120 21324 60172
rect 26976 60120 27028 60172
rect 21180 60095 21232 60104
rect 21180 60061 21189 60095
rect 21189 60061 21223 60095
rect 21223 60061 21232 60095
rect 22284 60095 22336 60104
rect 21180 60052 21232 60061
rect 22284 60061 22293 60095
rect 22293 60061 22327 60095
rect 22327 60061 22336 60095
rect 22284 60052 22336 60061
rect 22652 60095 22704 60104
rect 22652 60061 22666 60095
rect 22666 60061 22700 60095
rect 22700 60061 22704 60095
rect 22652 60052 22704 60061
rect 23020 60052 23072 60104
rect 23848 60095 23900 60104
rect 23848 60061 23851 60095
rect 23851 60061 23900 60095
rect 23848 60052 23900 60061
rect 23940 60095 23992 60104
rect 23940 60061 23966 60095
rect 23966 60061 23992 60095
rect 23940 60052 23992 60061
rect 24768 60052 24820 60104
rect 25136 60095 25188 60104
rect 25136 60061 25145 60095
rect 25145 60061 25179 60095
rect 25179 60061 25188 60095
rect 25136 60052 25188 60061
rect 25228 60095 25280 60104
rect 25228 60061 25237 60095
rect 25237 60061 25271 60095
rect 25271 60061 25280 60095
rect 25504 60095 25556 60104
rect 25228 60052 25280 60061
rect 25504 60061 25513 60095
rect 25513 60061 25547 60095
rect 25547 60061 25556 60095
rect 25504 60052 25556 60061
rect 2504 59916 2556 59968
rect 17684 59959 17736 59968
rect 17684 59925 17693 59959
rect 17693 59925 17727 59959
rect 17727 59925 17736 59959
rect 17684 59916 17736 59925
rect 22560 60027 22612 60036
rect 22560 59993 22569 60027
rect 22569 59993 22603 60027
rect 22603 59993 22612 60027
rect 22560 59984 22612 59993
rect 22744 59984 22796 60036
rect 23572 60027 23624 60036
rect 23572 59993 23581 60027
rect 23581 59993 23615 60027
rect 23615 59993 23624 60027
rect 23572 59984 23624 59993
rect 24952 59984 25004 60036
rect 25964 60095 26016 60104
rect 25964 60061 25973 60095
rect 25973 60061 26007 60095
rect 26007 60061 26016 60095
rect 25964 60052 26016 60061
rect 26424 60052 26476 60104
rect 26884 60095 26936 60104
rect 26884 60061 26894 60095
rect 26894 60061 26928 60095
rect 26928 60061 26936 60095
rect 27160 60095 27212 60104
rect 26884 60052 26936 60061
rect 27160 60061 27169 60095
rect 27169 60061 27203 60095
rect 27203 60061 27212 60095
rect 27160 60052 27212 60061
rect 27252 60095 27304 60104
rect 27252 60061 27266 60095
rect 27266 60061 27300 60095
rect 27300 60061 27304 60095
rect 28172 60120 28224 60172
rect 27988 60095 28040 60104
rect 27252 60052 27304 60061
rect 27988 60061 27997 60095
rect 27997 60061 28031 60095
rect 28031 60061 28040 60095
rect 27988 60052 28040 60061
rect 28080 60095 28132 60104
rect 28080 60061 28090 60095
rect 28090 60061 28124 60095
rect 28124 60061 28132 60095
rect 28724 60188 28776 60240
rect 28816 60188 28868 60240
rect 28540 60120 28592 60172
rect 29644 60120 29696 60172
rect 30104 60120 30156 60172
rect 28080 60052 28132 60061
rect 28724 60052 28776 60104
rect 29000 60052 29052 60104
rect 29184 60095 29236 60104
rect 29184 60061 29193 60095
rect 29193 60061 29227 60095
rect 29227 60061 29236 60095
rect 29184 60052 29236 60061
rect 28816 59984 28868 60036
rect 29092 59984 29144 60036
rect 30196 60095 30248 60104
rect 30196 60061 30210 60095
rect 30210 60061 30244 60095
rect 30244 60061 30248 60095
rect 33784 60095 33836 60104
rect 30196 60052 30248 60061
rect 33784 60061 33793 60095
rect 33793 60061 33827 60095
rect 33827 60061 33836 60095
rect 33784 60052 33836 60061
rect 34152 60095 34204 60104
rect 34152 60061 34161 60095
rect 34161 60061 34195 60095
rect 34195 60061 34204 60095
rect 34152 60052 34204 60061
rect 37188 60120 37240 60172
rect 56232 60188 56284 60240
rect 41880 60163 41932 60172
rect 41880 60129 41889 60163
rect 41889 60129 41923 60163
rect 41923 60129 41932 60163
rect 41880 60120 41932 60129
rect 53748 60120 53800 60172
rect 30012 60027 30064 60036
rect 30012 59993 30021 60027
rect 30021 59993 30055 60027
rect 30055 59993 30064 60027
rect 30012 59984 30064 59993
rect 36636 60052 36688 60104
rect 41604 60095 41656 60104
rect 41604 60061 41613 60095
rect 41613 60061 41647 60095
rect 41647 60061 41656 60095
rect 41604 60052 41656 60061
rect 41788 60052 41840 60104
rect 41972 60095 42024 60104
rect 41972 60061 41981 60095
rect 41981 60061 42015 60095
rect 42015 60061 42024 60095
rect 41972 60052 42024 60061
rect 35624 59984 35676 60036
rect 43260 60095 43312 60104
rect 43260 60061 43269 60095
rect 43269 60061 43303 60095
rect 43303 60061 43312 60095
rect 43260 60052 43312 60061
rect 56508 60095 56560 60104
rect 42616 60027 42668 60036
rect 42616 59993 42625 60027
rect 42625 59993 42659 60027
rect 42659 59993 42668 60027
rect 42616 59984 42668 59993
rect 56508 60061 56517 60095
rect 56517 60061 56551 60095
rect 56551 60061 56560 60095
rect 56508 60052 56560 60061
rect 57244 60095 57296 60104
rect 57244 60061 57253 60095
rect 57253 60061 57287 60095
rect 57287 60061 57296 60095
rect 57244 60052 57296 60061
rect 57980 60095 58032 60104
rect 57980 60061 57989 60095
rect 57989 60061 58023 60095
rect 58023 60061 58032 60095
rect 57980 60052 58032 60061
rect 50436 59984 50488 60036
rect 58440 59984 58492 60036
rect 25872 59916 25924 59968
rect 26240 59916 26292 59968
rect 26424 59959 26476 59968
rect 26424 59925 26433 59959
rect 26433 59925 26467 59959
rect 26467 59925 26476 59959
rect 26424 59916 26476 59925
rect 27528 59916 27580 59968
rect 29276 59916 29328 59968
rect 30656 59959 30708 59968
rect 30656 59925 30665 59959
rect 30665 59925 30699 59959
rect 30699 59925 30708 59959
rect 30656 59916 30708 59925
rect 33232 59959 33284 59968
rect 33232 59925 33241 59959
rect 33241 59925 33275 59959
rect 33275 59925 33284 59959
rect 33232 59916 33284 59925
rect 41052 59959 41104 59968
rect 41052 59925 41061 59959
rect 41061 59925 41095 59959
rect 41095 59925 41104 59959
rect 41052 59916 41104 59925
rect 56600 59959 56652 59968
rect 56600 59925 56609 59959
rect 56609 59925 56643 59959
rect 56643 59925 56652 59959
rect 56600 59916 56652 59925
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 1768 59644 1820 59696
rect 6736 59687 6788 59696
rect 6736 59653 6745 59687
rect 6745 59653 6779 59687
rect 6779 59653 6788 59687
rect 23572 59712 23624 59764
rect 25504 59712 25556 59764
rect 6736 59644 6788 59653
rect 15292 59644 15344 59696
rect 19248 59644 19300 59696
rect 22652 59644 22704 59696
rect 24584 59687 24636 59696
rect 24584 59653 24593 59687
rect 24593 59653 24627 59687
rect 24627 59653 24636 59687
rect 24584 59644 24636 59653
rect 1584 59619 1636 59628
rect 1584 59585 1593 59619
rect 1593 59585 1627 59619
rect 1627 59585 1636 59619
rect 1584 59576 1636 59585
rect 5540 59576 5592 59628
rect 6828 59619 6880 59628
rect 6828 59585 6837 59619
rect 6837 59585 6871 59619
rect 6871 59585 6880 59619
rect 6828 59576 6880 59585
rect 7012 59576 7064 59628
rect 18788 59619 18840 59628
rect 18788 59585 18797 59619
rect 18797 59585 18831 59619
rect 18831 59585 18840 59619
rect 18788 59576 18840 59585
rect 19156 59619 19208 59628
rect 19156 59585 19170 59619
rect 19170 59585 19204 59619
rect 19204 59585 19208 59619
rect 19156 59576 19208 59585
rect 22192 59576 22244 59628
rect 19432 59508 19484 59560
rect 24768 59576 24820 59628
rect 26792 59712 26844 59764
rect 29184 59712 29236 59764
rect 30656 59712 30708 59764
rect 33784 59712 33836 59764
rect 43260 59712 43312 59764
rect 56232 59712 56284 59764
rect 58256 59755 58308 59764
rect 58256 59721 58265 59755
rect 58265 59721 58299 59755
rect 58299 59721 58308 59755
rect 58256 59712 58308 59721
rect 25872 59687 25924 59696
rect 25872 59653 25881 59687
rect 25881 59653 25915 59687
rect 25915 59653 25924 59687
rect 25872 59644 25924 59653
rect 26976 59644 27028 59696
rect 30104 59644 30156 59696
rect 56416 59644 56468 59696
rect 25780 59619 25832 59628
rect 25780 59585 25789 59619
rect 25789 59585 25823 59619
rect 25823 59585 25832 59619
rect 25780 59576 25832 59585
rect 26240 59576 26292 59628
rect 30012 59576 30064 59628
rect 35532 59576 35584 59628
rect 21088 59440 21140 59492
rect 1768 59415 1820 59424
rect 1768 59381 1777 59415
rect 1777 59381 1811 59415
rect 1811 59381 1820 59415
rect 1768 59372 1820 59381
rect 2320 59372 2372 59424
rect 6828 59372 6880 59424
rect 18512 59415 18564 59424
rect 18512 59381 18521 59415
rect 18521 59381 18555 59415
rect 18555 59381 18564 59415
rect 18512 59372 18564 59381
rect 19156 59372 19208 59424
rect 19248 59372 19300 59424
rect 25136 59440 25188 59492
rect 25596 59440 25648 59492
rect 26148 59508 26200 59560
rect 42708 59551 42760 59560
rect 42708 59517 42717 59551
rect 42717 59517 42751 59551
rect 42751 59517 42760 59551
rect 42708 59508 42760 59517
rect 42800 59508 42852 59560
rect 43260 59619 43312 59628
rect 43260 59585 43269 59619
rect 43269 59585 43303 59619
rect 43303 59585 43312 59619
rect 43260 59576 43312 59585
rect 53104 59576 53156 59628
rect 58164 59619 58216 59628
rect 58164 59585 58173 59619
rect 58173 59585 58207 59619
rect 58207 59585 58216 59619
rect 58164 59576 58216 59585
rect 25780 59440 25832 59492
rect 56324 59440 56376 59492
rect 25964 59372 26016 59424
rect 27988 59372 28040 59424
rect 29828 59372 29880 59424
rect 30012 59372 30064 59424
rect 55588 59372 55640 59424
rect 57152 59372 57204 59424
rect 58992 59372 59044 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 1768 59168 1820 59220
rect 6000 59100 6052 59152
rect 26884 59032 26936 59084
rect 848 58964 900 59016
rect 37188 59007 37240 59016
rect 37188 58973 37197 59007
rect 37197 58973 37231 59007
rect 37231 58973 37240 59007
rect 37188 58964 37240 58973
rect 37280 59007 37332 59016
rect 37280 58973 37289 59007
rect 37289 58973 37323 59007
rect 37323 58973 37332 59007
rect 37556 59007 37608 59016
rect 37280 58964 37332 58973
rect 37556 58973 37565 59007
rect 37565 58973 37599 59007
rect 37599 58973 37608 59007
rect 37556 58964 37608 58973
rect 40776 59007 40828 59016
rect 34520 58896 34572 58948
rect 40776 58973 40785 59007
rect 40785 58973 40819 59007
rect 40819 58973 40828 59007
rect 40776 58964 40828 58973
rect 41236 58964 41288 59016
rect 41420 58964 41472 59016
rect 41880 58964 41932 59016
rect 58348 59100 58400 59152
rect 57152 59007 57204 59016
rect 57152 58973 57161 59007
rect 57161 58973 57195 59007
rect 57195 58973 57204 59007
rect 57152 58964 57204 58973
rect 57888 59007 57940 59016
rect 57888 58973 57897 59007
rect 57897 58973 57931 59007
rect 57931 58973 57940 59007
rect 57888 58964 57940 58973
rect 58532 58896 58584 58948
rect 40868 58828 40920 58880
rect 57336 58871 57388 58880
rect 57336 58837 57345 58871
rect 57345 58837 57379 58871
rect 57379 58837 57388 58871
rect 57336 58828 57388 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 18788 58624 18840 58676
rect 57336 58624 57388 58676
rect 58164 58599 58216 58608
rect 58164 58565 58173 58599
rect 58173 58565 58207 58599
rect 58207 58565 58216 58599
rect 58164 58556 58216 58565
rect 1584 58531 1636 58540
rect 1584 58497 1593 58531
rect 1593 58497 1627 58531
rect 1627 58497 1636 58531
rect 1584 58488 1636 58497
rect 1768 58463 1820 58472
rect 1768 58429 1777 58463
rect 1777 58429 1811 58463
rect 1811 58429 1820 58463
rect 1768 58420 1820 58429
rect 2044 58420 2096 58472
rect 40776 58531 40828 58540
rect 40776 58497 40785 58531
rect 40785 58497 40819 58531
rect 40819 58497 40828 58531
rect 41144 58531 41196 58540
rect 40776 58488 40828 58497
rect 41144 58497 41153 58531
rect 41153 58497 41187 58531
rect 41187 58497 41196 58531
rect 41144 58488 41196 58497
rect 41420 58488 41472 58540
rect 39304 58420 39356 58472
rect 40408 58327 40460 58336
rect 40408 58293 40417 58327
rect 40417 58293 40451 58327
rect 40451 58293 40460 58327
rect 40408 58284 40460 58293
rect 56508 58284 56560 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 52920 57944 52972 57996
rect 1584 57919 1636 57928
rect 1584 57885 1593 57919
rect 1593 57885 1627 57919
rect 1627 57885 1636 57919
rect 1584 57876 1636 57885
rect 17224 57808 17276 57860
rect 57980 57851 58032 57860
rect 57980 57817 57989 57851
rect 57989 57817 58023 57851
rect 58023 57817 58032 57851
rect 57980 57808 58032 57817
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1584 57443 1636 57452
rect 1584 57409 1593 57443
rect 1593 57409 1627 57443
rect 1627 57409 1636 57443
rect 1584 57400 1636 57409
rect 29644 57196 29696 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 26976 56992 27028 57044
rect 34520 56992 34572 57044
rect 28356 56924 28408 56976
rect 1584 56831 1636 56840
rect 1584 56797 1593 56831
rect 1593 56797 1627 56831
rect 1627 56797 1636 56831
rect 1584 56788 1636 56797
rect 22468 56788 22520 56840
rect 33784 56788 33836 56840
rect 25688 56720 25740 56772
rect 27620 56652 27672 56704
rect 33324 56695 33376 56704
rect 33324 56661 33333 56695
rect 33333 56661 33367 56695
rect 33367 56661 33376 56695
rect 33324 56652 33376 56661
rect 35624 56831 35676 56840
rect 35624 56797 35633 56831
rect 35633 56797 35667 56831
rect 35667 56797 35676 56831
rect 35900 56831 35952 56840
rect 35624 56788 35676 56797
rect 35900 56797 35909 56831
rect 35909 56797 35943 56831
rect 35943 56797 35952 56831
rect 35900 56788 35952 56797
rect 35992 56831 36044 56840
rect 35992 56797 36001 56831
rect 36001 56797 36035 56831
rect 36035 56797 36044 56831
rect 35992 56788 36044 56797
rect 52460 56924 52512 56976
rect 56508 56856 56560 56908
rect 57888 56831 57940 56840
rect 57888 56797 57897 56831
rect 57897 56797 57931 56831
rect 57931 56797 57940 56831
rect 57888 56788 57940 56797
rect 58072 56720 58124 56772
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 35624 56448 35676 56500
rect 36452 56448 36504 56500
rect 37188 56448 37240 56500
rect 41420 56448 41472 56500
rect 27620 56380 27672 56432
rect 58164 56423 58216 56432
rect 29276 56355 29328 56364
rect 29276 56321 29285 56355
rect 29285 56321 29319 56355
rect 29319 56321 29328 56355
rect 29276 56312 29328 56321
rect 29644 56355 29696 56364
rect 29644 56321 29653 56355
rect 29653 56321 29687 56355
rect 29687 56321 29696 56355
rect 29644 56312 29696 56321
rect 30012 56312 30064 56364
rect 35532 56312 35584 56364
rect 36452 56355 36504 56364
rect 36452 56321 36461 56355
rect 36461 56321 36495 56355
rect 36495 56321 36504 56355
rect 36452 56312 36504 56321
rect 58164 56389 58173 56423
rect 58173 56389 58207 56423
rect 58207 56389 58216 56423
rect 58164 56380 58216 56389
rect 27344 56244 27396 56296
rect 39948 56244 40000 56296
rect 46756 56312 46808 56364
rect 41420 56287 41472 56296
rect 41420 56253 41429 56287
rect 41429 56253 41463 56287
rect 41463 56253 41472 56287
rect 41420 56244 41472 56253
rect 32404 56108 32456 56160
rect 42248 56108 42300 56160
rect 52460 56108 52512 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 58348 55947 58400 55956
rect 58348 55913 58357 55947
rect 58357 55913 58391 55947
rect 58391 55913 58400 55947
rect 58348 55904 58400 55913
rect 23572 55700 23624 55752
rect 27528 55768 27580 55820
rect 1676 55675 1728 55684
rect 1676 55641 1685 55675
rect 1685 55641 1719 55675
rect 1719 55641 1728 55675
rect 1676 55632 1728 55641
rect 26608 55675 26660 55684
rect 26608 55641 26617 55675
rect 26617 55641 26651 55675
rect 26651 55641 26660 55675
rect 26608 55632 26660 55641
rect 27344 55743 27396 55752
rect 27344 55709 27353 55743
rect 27353 55709 27387 55743
rect 27387 55709 27396 55743
rect 27344 55700 27396 55709
rect 30012 55700 30064 55752
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 1584 55267 1636 55276
rect 1584 55233 1593 55267
rect 1593 55233 1627 55267
rect 1627 55233 1636 55267
rect 1584 55224 1636 55233
rect 39396 55292 39448 55344
rect 39948 55292 40000 55344
rect 40040 55199 40092 55208
rect 40040 55165 40049 55199
rect 40049 55165 40083 55199
rect 40083 55165 40092 55199
rect 40040 55156 40092 55165
rect 41420 55292 41472 55344
rect 44180 55224 44232 55276
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 18052 54680 18104 54732
rect 23572 54723 23624 54732
rect 23572 54689 23581 54723
rect 23581 54689 23615 54723
rect 23615 54689 23624 54723
rect 23572 54680 23624 54689
rect 26056 54680 26108 54732
rect 1676 54587 1728 54596
rect 1676 54553 1685 54587
rect 1685 54553 1719 54587
rect 1719 54553 1728 54587
rect 1676 54544 1728 54553
rect 22836 54587 22888 54596
rect 22836 54553 22845 54587
rect 22845 54553 22879 54587
rect 22879 54553 22888 54587
rect 22836 54544 22888 54553
rect 23940 54612 23992 54664
rect 30012 54612 30064 54664
rect 58348 54655 58400 54664
rect 58348 54621 58357 54655
rect 58357 54621 58391 54655
rect 58391 54621 58400 54655
rect 58348 54612 58400 54621
rect 27528 54476 27580 54528
rect 45376 54476 45428 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1584 54179 1636 54188
rect 1584 54145 1593 54179
rect 1593 54145 1627 54179
rect 1627 54145 1636 54179
rect 1584 54136 1636 54145
rect 10968 53932 11020 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 40868 53660 40920 53712
rect 41880 53660 41932 53712
rect 10968 53592 11020 53644
rect 30012 53524 30064 53576
rect 36452 53524 36504 53576
rect 46112 53592 46164 53644
rect 41420 53524 41472 53576
rect 40408 53388 40460 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 23940 53184 23992 53236
rect 27528 53116 27580 53168
rect 1676 53091 1728 53100
rect 1676 53057 1685 53091
rect 1685 53057 1719 53091
rect 1719 53057 1728 53091
rect 1676 53048 1728 53057
rect 23848 53048 23900 53100
rect 24308 53091 24360 53100
rect 24308 53057 24317 53091
rect 24317 53057 24351 53091
rect 24351 53057 24360 53091
rect 24308 53048 24360 53057
rect 27436 53048 27488 53100
rect 39672 53048 39724 53100
rect 23572 52844 23624 52896
rect 58348 52887 58400 52896
rect 58348 52853 58357 52887
rect 58357 52853 58391 52887
rect 58391 52853 58400 52887
rect 58348 52844 58400 52853
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 1860 52547 1912 52556
rect 1860 52513 1869 52547
rect 1869 52513 1903 52547
rect 1903 52513 1912 52547
rect 1860 52504 1912 52513
rect 34612 52504 34664 52556
rect 35992 52504 36044 52556
rect 1584 52479 1636 52488
rect 1584 52445 1593 52479
rect 1593 52445 1627 52479
rect 1627 52445 1636 52479
rect 1584 52436 1636 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1676 52003 1728 52012
rect 1676 51969 1685 52003
rect 1685 51969 1719 52003
rect 1719 51969 1728 52003
rect 1676 51960 1728 51969
rect 6828 52003 6880 52012
rect 6828 51969 6837 52003
rect 6837 51969 6871 52003
rect 6871 51969 6880 52003
rect 6828 51960 6880 51969
rect 7104 52003 7156 52012
rect 7104 51969 7113 52003
rect 7113 51969 7147 52003
rect 7147 51969 7156 52003
rect 7104 51960 7156 51969
rect 6736 51756 6788 51808
rect 17316 51756 17368 51808
rect 26332 51756 26384 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58348 51391 58400 51400
rect 58348 51357 58357 51391
rect 58357 51357 58391 51391
rect 58391 51357 58400 51391
rect 58348 51348 58400 51357
rect 1676 51323 1728 51332
rect 1676 51289 1685 51323
rect 1685 51289 1719 51323
rect 1719 51289 1728 51323
rect 1676 51280 1728 51289
rect 3976 51280 4028 51332
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4620 51008 4672 51060
rect 3976 50983 4028 50992
rect 3976 50949 3985 50983
rect 3985 50949 4019 50983
rect 4019 50949 4028 50983
rect 3976 50940 4028 50949
rect 3884 50915 3936 50924
rect 3884 50881 3893 50915
rect 3893 50881 3927 50915
rect 3927 50881 3936 50915
rect 3884 50872 3936 50881
rect 7104 50872 7156 50924
rect 7564 50872 7616 50924
rect 2596 50804 2648 50856
rect 5908 50668 5960 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 24216 50328 24268 50380
rect 39304 50328 39356 50380
rect 45008 50260 45060 50312
rect 1676 50235 1728 50244
rect 1676 50201 1685 50235
rect 1685 50201 1719 50235
rect 1719 50201 1728 50235
rect 1676 50192 1728 50201
rect 2044 50192 2096 50244
rect 57888 50124 57940 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 1584 49827 1636 49836
rect 1584 49793 1593 49827
rect 1593 49793 1627 49827
rect 1627 49793 1636 49827
rect 1584 49784 1636 49793
rect 22284 49716 22336 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 1676 49147 1728 49156
rect 1676 49113 1685 49147
rect 1685 49113 1719 49147
rect 1719 49113 1728 49147
rect 1676 49104 1728 49113
rect 7840 49104 7892 49156
rect 34796 49104 34848 49156
rect 41788 49104 41840 49156
rect 54576 49104 54628 49156
rect 57980 49147 58032 49156
rect 57980 49113 57989 49147
rect 57989 49113 58023 49147
rect 58023 49113 58032 49147
rect 57980 49104 58032 49113
rect 15844 49036 15896 49088
rect 51908 49036 51960 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 1676 48739 1728 48748
rect 1676 48705 1685 48739
rect 1685 48705 1719 48739
rect 1719 48705 1728 48739
rect 1676 48696 1728 48705
rect 1952 48560 2004 48612
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 24768 48220 24820 48272
rect 25412 48220 25464 48272
rect 36268 47948 36320 48000
rect 57244 48059 57296 48068
rect 57244 48025 57253 48059
rect 57253 48025 57287 48059
rect 57287 48025 57296 48059
rect 57244 48016 57296 48025
rect 57980 48059 58032 48068
rect 57980 48025 57989 48059
rect 57989 48025 58023 48059
rect 58023 48025 58032 48059
rect 57980 48016 58032 48025
rect 58072 47991 58124 48000
rect 58072 47957 58081 47991
rect 58081 47957 58115 47991
rect 58115 47957 58124 47991
rect 58072 47948 58124 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 46296 47744 46348 47796
rect 58072 47744 58124 47796
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 3332 47540 3384 47592
rect 20260 47540 20312 47592
rect 22192 47540 22244 47592
rect 39396 47540 39448 47592
rect 5448 47472 5500 47524
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 1584 47039 1636 47048
rect 1584 47005 1593 47039
rect 1593 47005 1627 47039
rect 1627 47005 1636 47039
rect 1584 46996 1636 47005
rect 57520 46996 57572 47048
rect 24860 46928 24912 46980
rect 57888 46860 57940 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 1584 46563 1636 46572
rect 1584 46529 1593 46563
rect 1593 46529 1627 46563
rect 1627 46529 1636 46563
rect 1584 46520 1636 46529
rect 19064 46384 19116 46436
rect 39120 46384 39172 46436
rect 20720 46316 20772 46368
rect 34244 46316 34296 46368
rect 54852 46316 54904 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1676 45883 1728 45892
rect 1676 45849 1685 45883
rect 1685 45849 1719 45883
rect 1719 45849 1728 45883
rect 1676 45840 1728 45849
rect 57980 45883 58032 45892
rect 57980 45849 57989 45883
rect 57989 45849 58023 45883
rect 58023 45849 58032 45883
rect 57980 45840 58032 45849
rect 17684 45772 17736 45824
rect 44916 45772 44968 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 17868 45568 17920 45620
rect 7564 45432 7616 45484
rect 17776 45500 17828 45552
rect 17684 45475 17736 45484
rect 17684 45441 17694 45475
rect 17694 45441 17728 45475
rect 17728 45441 17736 45475
rect 17684 45432 17736 45441
rect 18236 45432 18288 45484
rect 20720 45500 20772 45552
rect 24124 45432 24176 45484
rect 39856 45500 39908 45552
rect 36452 45475 36504 45484
rect 36452 45441 36461 45475
rect 36461 45441 36495 45475
rect 36495 45441 36504 45475
rect 36452 45432 36504 45441
rect 37096 45432 37148 45484
rect 19800 45296 19852 45348
rect 30564 45296 30616 45348
rect 37556 45296 37608 45348
rect 18236 45271 18288 45280
rect 18236 45237 18245 45271
rect 18245 45237 18279 45271
rect 18279 45237 18288 45271
rect 18236 45228 18288 45237
rect 18328 45228 18380 45280
rect 20812 45228 20864 45280
rect 21180 45228 21232 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 17776 45024 17828 45076
rect 19800 45024 19852 45076
rect 30564 45024 30616 45076
rect 1584 44863 1636 44872
rect 1584 44829 1593 44863
rect 1593 44829 1627 44863
rect 1627 44829 1636 44863
rect 1584 44820 1636 44829
rect 22836 44820 22888 44872
rect 30748 44820 30800 44872
rect 37648 44863 37700 44872
rect 37648 44829 37657 44863
rect 37657 44829 37691 44863
rect 37691 44829 37700 44863
rect 37648 44820 37700 44829
rect 57060 44888 57112 44940
rect 31024 44752 31076 44804
rect 37096 44752 37148 44804
rect 37372 44684 37424 44736
rect 50896 44820 50948 44872
rect 57244 44795 57296 44804
rect 57244 44761 57253 44795
rect 57253 44761 57287 44795
rect 57287 44761 57296 44795
rect 57244 44752 57296 44761
rect 57888 44752 57940 44804
rect 58256 44727 58308 44736
rect 58256 44693 58265 44727
rect 58265 44693 58299 44727
rect 58299 44693 58308 44727
rect 58256 44684 58308 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 1676 44387 1728 44396
rect 1676 44353 1685 44387
rect 1685 44353 1719 44387
rect 1719 44353 1728 44387
rect 1676 44344 1728 44353
rect 17132 44140 17184 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 35440 43911 35492 43920
rect 35440 43877 35449 43911
rect 35449 43877 35483 43911
rect 35483 43877 35492 43911
rect 35440 43868 35492 43877
rect 17132 43800 17184 43852
rect 1676 43707 1728 43716
rect 1676 43673 1685 43707
rect 1685 43673 1719 43707
rect 1719 43673 1728 43707
rect 1676 43664 1728 43673
rect 34060 43664 34112 43716
rect 33968 43596 34020 43648
rect 35164 43707 35216 43716
rect 35164 43673 35173 43707
rect 35173 43673 35207 43707
rect 35207 43673 35216 43707
rect 50804 43732 50856 43784
rect 35164 43664 35216 43673
rect 36176 43664 36228 43716
rect 58164 43707 58216 43716
rect 58164 43673 58173 43707
rect 58173 43673 58207 43707
rect 58207 43673 58216 43707
rect 58164 43664 58216 43673
rect 36452 43596 36504 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 6736 43392 6788 43444
rect 22008 43392 22060 43444
rect 37188 43392 37240 43444
rect 54300 43392 54352 43444
rect 34244 43367 34296 43376
rect 34244 43333 34253 43367
rect 34253 43333 34287 43367
rect 34287 43333 34296 43367
rect 34244 43324 34296 43333
rect 1584 43299 1636 43308
rect 1584 43265 1593 43299
rect 1593 43265 1627 43299
rect 1627 43265 1636 43299
rect 1584 43256 1636 43265
rect 33968 43299 34020 43308
rect 33968 43265 33977 43299
rect 33977 43265 34011 43299
rect 34011 43265 34020 43299
rect 33968 43256 34020 43265
rect 34060 43256 34112 43308
rect 37372 43256 37424 43308
rect 1768 43095 1820 43104
rect 1768 43061 1777 43095
rect 1777 43061 1811 43095
rect 1811 43061 1820 43095
rect 1768 43052 1820 43061
rect 34520 43095 34572 43104
rect 34520 43061 34529 43095
rect 34529 43061 34563 43095
rect 34563 43061 34572 43095
rect 34520 43052 34572 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 24308 42712 24360 42764
rect 36176 42780 36228 42832
rect 1768 42644 1820 42696
rect 33508 42712 33560 42764
rect 32956 42551 33008 42560
rect 32956 42517 32965 42551
rect 32965 42517 32999 42551
rect 32999 42517 33008 42551
rect 32956 42508 33008 42517
rect 33968 42687 34020 42696
rect 33968 42653 33977 42687
rect 33977 42653 34011 42687
rect 34011 42653 34020 42687
rect 33968 42644 34020 42653
rect 36912 42687 36964 42696
rect 36912 42653 36921 42687
rect 36921 42653 36955 42687
rect 36955 42653 36964 42687
rect 36912 42644 36964 42653
rect 37188 42687 37240 42696
rect 37188 42653 37197 42687
rect 37197 42653 37231 42687
rect 37231 42653 37240 42687
rect 37188 42644 37240 42653
rect 37372 42644 37424 42696
rect 37096 42619 37148 42628
rect 37096 42585 37105 42619
rect 37105 42585 37139 42619
rect 37139 42585 37148 42619
rect 37096 42576 37148 42585
rect 57060 42619 57112 42628
rect 57060 42585 57069 42619
rect 57069 42585 57103 42619
rect 57103 42585 57112 42619
rect 57060 42576 57112 42585
rect 57980 42619 58032 42628
rect 57980 42585 57989 42619
rect 57989 42585 58023 42619
rect 58023 42585 58032 42619
rect 57980 42576 58032 42585
rect 58624 42576 58676 42628
rect 57152 42551 57204 42560
rect 57152 42517 57161 42551
rect 57161 42517 57195 42551
rect 57195 42517 57204 42551
rect 57152 42508 57204 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 23480 42304 23532 42356
rect 37096 42304 37148 42356
rect 1676 42211 1728 42220
rect 1676 42177 1685 42211
rect 1685 42177 1719 42211
rect 1719 42177 1728 42211
rect 1676 42168 1728 42177
rect 5448 42100 5500 42152
rect 20904 42100 20956 42152
rect 5540 42032 5592 42084
rect 5632 41964 5684 42016
rect 42892 42032 42944 42084
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 23756 41692 23808 41744
rect 24124 41624 24176 41676
rect 24032 41556 24084 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 24584 41531 24636 41540
rect 24584 41497 24593 41531
rect 24593 41497 24627 41531
rect 24627 41497 24636 41531
rect 24584 41488 24636 41497
rect 1860 41420 1912 41472
rect 20812 41420 20864 41472
rect 51724 41556 51776 41608
rect 57244 41531 57296 41540
rect 57244 41497 57253 41531
rect 57253 41497 57287 41531
rect 57287 41497 57296 41531
rect 57244 41488 57296 41497
rect 57888 41488 57940 41540
rect 38568 41420 38620 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1676 41123 1728 41132
rect 1676 41089 1685 41123
rect 1685 41089 1719 41123
rect 1719 41089 1728 41123
rect 1676 41080 1728 41089
rect 5540 40944 5592 40996
rect 22376 40944 22428 40996
rect 20536 40876 20588 40928
rect 36820 40876 36872 40928
rect 48964 40876 49016 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 20168 40672 20220 40724
rect 41052 40672 41104 40724
rect 56968 40511 57020 40520
rect 56968 40477 56977 40511
rect 56977 40477 57011 40511
rect 57011 40477 57020 40511
rect 56968 40468 57020 40477
rect 57796 40468 57848 40520
rect 1676 40443 1728 40452
rect 1676 40409 1685 40443
rect 1685 40409 1719 40443
rect 1719 40409 1728 40443
rect 1676 40400 1728 40409
rect 44088 40400 44140 40452
rect 11060 40332 11112 40384
rect 57888 40332 57940 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 15844 40060 15896 40112
rect 19340 40060 19392 40112
rect 26608 40060 26660 40112
rect 30288 40060 30340 40112
rect 33324 40060 33376 40112
rect 38568 40060 38620 40112
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 15844 39516 15896 39568
rect 2320 39423 2372 39432
rect 2320 39389 2329 39423
rect 2329 39389 2363 39423
rect 2363 39389 2372 39423
rect 2320 39380 2372 39389
rect 20628 39423 20680 39432
rect 20628 39389 20637 39423
rect 20637 39389 20671 39423
rect 20671 39389 20680 39423
rect 20628 39380 20680 39389
rect 1676 39355 1728 39364
rect 1676 39321 1685 39355
rect 1685 39321 1719 39355
rect 1719 39321 1728 39355
rect 1676 39312 1728 39321
rect 20536 39312 20588 39364
rect 22100 39380 22152 39432
rect 20812 39355 20864 39364
rect 20812 39321 20821 39355
rect 20821 39321 20855 39355
rect 20855 39321 20864 39355
rect 57060 39355 57112 39364
rect 20812 39312 20864 39321
rect 57060 39321 57069 39355
rect 57069 39321 57103 39355
rect 57103 39321 57112 39355
rect 57060 39312 57112 39321
rect 57980 39355 58032 39364
rect 57980 39321 57989 39355
rect 57989 39321 58023 39355
rect 58023 39321 58032 39355
rect 57980 39312 58032 39321
rect 2596 39244 2648 39296
rect 21364 39244 21416 39296
rect 35532 39244 35584 39296
rect 58072 39287 58124 39296
rect 58072 39253 58081 39287
rect 58081 39253 58115 39287
rect 58115 39253 58124 39287
rect 58072 39244 58124 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 34060 39040 34112 39092
rect 9312 38972 9364 39024
rect 1676 38947 1728 38956
rect 1676 38913 1685 38947
rect 1685 38913 1719 38947
rect 1719 38913 1728 38947
rect 1676 38904 1728 38913
rect 34060 38947 34112 38956
rect 34060 38913 34069 38947
rect 34069 38913 34103 38947
rect 34103 38913 34112 38947
rect 34060 38904 34112 38913
rect 26056 38836 26108 38888
rect 34428 38947 34480 38956
rect 34428 38913 34442 38947
rect 34442 38913 34476 38947
rect 34476 38913 34480 38947
rect 47676 39040 47728 39092
rect 58072 39040 58124 39092
rect 34428 38904 34480 38913
rect 45836 38904 45888 38956
rect 4804 38768 4856 38820
rect 34612 38811 34664 38820
rect 34612 38777 34621 38811
rect 34621 38777 34655 38811
rect 34655 38777 34664 38811
rect 34612 38768 34664 38777
rect 38568 38700 38620 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 22744 38335 22796 38344
rect 22744 38301 22753 38335
rect 22753 38301 22787 38335
rect 22787 38301 22796 38335
rect 22744 38292 22796 38301
rect 22928 38335 22980 38344
rect 22928 38301 22935 38335
rect 22935 38301 22980 38335
rect 22928 38292 22980 38301
rect 23480 38360 23532 38412
rect 23204 38335 23256 38344
rect 23204 38301 23218 38335
rect 23218 38301 23252 38335
rect 23252 38301 23256 38335
rect 23204 38292 23256 38301
rect 49056 38292 49108 38344
rect 1676 38267 1728 38276
rect 1676 38233 1685 38267
rect 1685 38233 1719 38267
rect 1719 38233 1728 38267
rect 1676 38224 1728 38233
rect 11060 38224 11112 38276
rect 23020 38267 23072 38276
rect 19432 38156 19484 38208
rect 23020 38233 23029 38267
rect 23029 38233 23063 38267
rect 23063 38233 23072 38267
rect 23020 38224 23072 38233
rect 58164 38267 58216 38276
rect 58164 38233 58173 38267
rect 58173 38233 58207 38267
rect 58207 38233 58216 38267
rect 58164 38224 58216 38233
rect 23664 38156 23716 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 20904 37995 20956 38004
rect 1676 37859 1728 37868
rect 1676 37825 1685 37859
rect 1685 37825 1719 37859
rect 1719 37825 1728 37859
rect 1676 37816 1728 37825
rect 4804 37859 4856 37868
rect 4804 37825 4813 37859
rect 4813 37825 4847 37859
rect 4847 37825 4856 37859
rect 4804 37816 4856 37825
rect 4988 37859 5040 37868
rect 4988 37825 4997 37859
rect 4997 37825 5031 37859
rect 5031 37825 5040 37859
rect 19248 37859 19300 37868
rect 4988 37816 5040 37825
rect 4068 37680 4120 37732
rect 19248 37825 19257 37859
rect 19257 37825 19291 37859
rect 19291 37825 19300 37859
rect 19248 37816 19300 37825
rect 19432 37884 19484 37936
rect 20904 37961 20913 37995
rect 20913 37961 20947 37995
rect 20947 37961 20956 37995
rect 20904 37952 20956 37961
rect 22928 37952 22980 38004
rect 38016 37952 38068 38004
rect 52000 37952 52052 38004
rect 58256 37952 58308 38004
rect 19524 37859 19576 37868
rect 19524 37825 19533 37859
rect 19533 37825 19567 37859
rect 19567 37825 19576 37859
rect 19524 37816 19576 37825
rect 19708 37859 19760 37868
rect 19708 37825 19741 37859
rect 19741 37825 19760 37859
rect 19708 37816 19760 37825
rect 24308 37816 24360 37868
rect 58072 37859 58124 37868
rect 58072 37825 58081 37859
rect 58081 37825 58115 37859
rect 58115 37825 58124 37859
rect 58072 37816 58124 37825
rect 19708 37680 19760 37732
rect 22560 37680 22612 37732
rect 47952 37748 48004 37800
rect 54024 37680 54076 37732
rect 6736 37612 6788 37664
rect 20076 37612 20128 37664
rect 20536 37655 20588 37664
rect 20536 37621 20545 37655
rect 20545 37621 20579 37655
rect 20579 37621 20588 37655
rect 20536 37612 20588 37621
rect 58256 37655 58308 37664
rect 58256 37621 58265 37655
rect 58265 37621 58299 37655
rect 58299 37621 58308 37655
rect 58256 37612 58308 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 22100 37408 22152 37460
rect 2044 37247 2096 37256
rect 2044 37213 2053 37247
rect 2053 37213 2087 37247
rect 2087 37213 2096 37247
rect 2044 37204 2096 37213
rect 6184 37204 6236 37256
rect 2228 37179 2280 37188
rect 2228 37145 2237 37179
rect 2237 37145 2271 37179
rect 2271 37145 2280 37179
rect 2228 37136 2280 37145
rect 2320 37179 2372 37188
rect 2320 37145 2329 37179
rect 2329 37145 2363 37179
rect 2363 37145 2372 37179
rect 2320 37136 2372 37145
rect 7564 37136 7616 37188
rect 21088 37272 21140 37324
rect 18420 37247 18472 37256
rect 18420 37213 18429 37247
rect 18429 37213 18463 37247
rect 18463 37213 18472 37247
rect 18420 37204 18472 37213
rect 20168 37204 20220 37256
rect 18696 37179 18748 37188
rect 18696 37145 18705 37179
rect 18705 37145 18739 37179
rect 18739 37145 18748 37179
rect 18696 37136 18748 37145
rect 19248 37136 19300 37188
rect 20260 37136 20312 37188
rect 16396 37068 16448 37120
rect 48964 37204 49016 37256
rect 58164 37179 58216 37188
rect 58164 37145 58173 37179
rect 58173 37145 58207 37179
rect 58207 37145 58216 37179
rect 58164 37136 58216 37145
rect 21640 37068 21692 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 2136 36796 2188 36848
rect 2596 36796 2648 36848
rect 6644 36839 6696 36848
rect 1952 36728 2004 36780
rect 2228 36771 2280 36780
rect 2228 36737 2237 36771
rect 2237 36737 2271 36771
rect 2271 36737 2280 36771
rect 2228 36728 2280 36737
rect 2688 36728 2740 36780
rect 3056 36771 3108 36780
rect 3056 36737 3065 36771
rect 3065 36737 3099 36771
rect 3099 36737 3108 36771
rect 3056 36728 3108 36737
rect 6644 36805 6653 36839
rect 6653 36805 6687 36839
rect 6687 36805 6696 36839
rect 6644 36796 6696 36805
rect 7012 36796 7064 36848
rect 18696 36796 18748 36848
rect 19064 36839 19116 36848
rect 19064 36805 19073 36839
rect 19073 36805 19107 36839
rect 19107 36805 19116 36839
rect 19064 36796 19116 36805
rect 6736 36703 6788 36712
rect 6736 36669 6745 36703
rect 6745 36669 6779 36703
rect 6779 36669 6788 36703
rect 6736 36660 6788 36669
rect 17960 36771 18012 36780
rect 17960 36737 17969 36771
rect 17969 36737 18003 36771
rect 18003 36737 18012 36771
rect 17960 36728 18012 36737
rect 7840 36660 7892 36712
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 18144 36660 18196 36712
rect 18880 36728 18932 36780
rect 19248 36728 19300 36780
rect 20076 36728 20128 36780
rect 20444 36703 20496 36712
rect 3240 36567 3292 36576
rect 3240 36533 3249 36567
rect 3249 36533 3283 36567
rect 3283 36533 3292 36567
rect 3240 36524 3292 36533
rect 20444 36669 20453 36703
rect 20453 36669 20487 36703
rect 20487 36669 20496 36703
rect 20444 36660 20496 36669
rect 19156 36592 19208 36644
rect 20536 36592 20588 36644
rect 23756 36728 23808 36780
rect 24308 36728 24360 36780
rect 22836 36660 22888 36712
rect 33968 36796 34020 36848
rect 53656 36728 53708 36780
rect 56600 36728 56652 36780
rect 33140 36660 33192 36712
rect 54576 36703 54628 36712
rect 54576 36669 54585 36703
rect 54585 36669 54619 36703
rect 54619 36669 54628 36703
rect 54576 36660 54628 36669
rect 55128 36592 55180 36644
rect 16672 36524 16724 36576
rect 18880 36524 18932 36576
rect 18972 36524 19024 36576
rect 23848 36524 23900 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 7196 36320 7248 36372
rect 7840 36320 7892 36372
rect 16396 36320 16448 36372
rect 19064 36320 19116 36372
rect 18880 36295 18932 36304
rect 2688 36184 2740 36236
rect 2504 36159 2556 36168
rect 2504 36125 2513 36159
rect 2513 36125 2547 36159
rect 2547 36125 2556 36159
rect 2504 36116 2556 36125
rect 1676 36091 1728 36100
rect 1676 36057 1685 36091
rect 1685 36057 1719 36091
rect 1719 36057 1728 36091
rect 1676 36048 1728 36057
rect 2596 36048 2648 36100
rect 2780 36091 2832 36100
rect 2780 36057 2789 36091
rect 2789 36057 2823 36091
rect 2823 36057 2832 36091
rect 2780 36048 2832 36057
rect 5172 36023 5224 36032
rect 5172 35989 5181 36023
rect 5181 35989 5215 36023
rect 5215 35989 5224 36023
rect 5172 35980 5224 35989
rect 5632 36159 5684 36168
rect 5632 36125 5641 36159
rect 5641 36125 5675 36159
rect 5675 36125 5684 36159
rect 5908 36159 5960 36168
rect 5632 36116 5684 36125
rect 5908 36125 5917 36159
rect 5917 36125 5951 36159
rect 5951 36125 5960 36159
rect 5908 36116 5960 36125
rect 6184 36159 6236 36168
rect 6184 36125 6193 36159
rect 6193 36125 6227 36159
rect 6227 36125 6236 36159
rect 6184 36116 6236 36125
rect 18880 36261 18889 36295
rect 18889 36261 18923 36295
rect 18923 36261 18932 36295
rect 18880 36252 18932 36261
rect 19432 36252 19484 36304
rect 32128 36320 32180 36372
rect 22468 36252 22520 36304
rect 23296 36252 23348 36304
rect 46204 36320 46256 36372
rect 54024 36363 54076 36372
rect 54024 36329 54033 36363
rect 54033 36329 54067 36363
rect 54067 36329 54076 36363
rect 54024 36320 54076 36329
rect 7012 36048 7064 36100
rect 7196 36116 7248 36168
rect 18328 36159 18380 36168
rect 18328 36125 18337 36159
rect 18337 36125 18371 36159
rect 18371 36125 18380 36159
rect 18328 36116 18380 36125
rect 18604 36159 18656 36168
rect 18604 36125 18613 36159
rect 18613 36125 18647 36159
rect 18647 36125 18656 36159
rect 18604 36116 18656 36125
rect 18788 36116 18840 36168
rect 19984 36159 20036 36168
rect 19984 36125 19993 36159
rect 19993 36125 20027 36159
rect 20027 36125 20036 36159
rect 19984 36116 20036 36125
rect 20352 36159 20404 36168
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20352 36116 20404 36125
rect 20536 36116 20588 36168
rect 20720 36116 20772 36168
rect 21088 36159 21140 36168
rect 21088 36125 21097 36159
rect 21097 36125 21131 36159
rect 21131 36125 21140 36159
rect 21088 36116 21140 36125
rect 21364 36159 21416 36168
rect 21364 36125 21373 36159
rect 21373 36125 21407 36159
rect 21407 36125 21416 36159
rect 21364 36116 21416 36125
rect 22468 36159 22520 36168
rect 22468 36125 22477 36159
rect 22477 36125 22511 36159
rect 22511 36125 22520 36159
rect 22468 36116 22520 36125
rect 19892 36048 19944 36100
rect 20812 36048 20864 36100
rect 22284 36048 22336 36100
rect 22836 36159 22888 36168
rect 22836 36125 22845 36159
rect 22845 36125 22879 36159
rect 22879 36125 22888 36159
rect 23664 36159 23716 36168
rect 22836 36116 22888 36125
rect 23664 36125 23673 36159
rect 23673 36125 23707 36159
rect 23707 36125 23716 36159
rect 23664 36116 23716 36125
rect 40776 36184 40828 36236
rect 40684 36159 40736 36168
rect 40684 36125 40693 36159
rect 40693 36125 40727 36159
rect 40727 36125 40736 36159
rect 40684 36116 40736 36125
rect 53472 36159 53524 36168
rect 53472 36125 53481 36159
rect 53481 36125 53515 36159
rect 53515 36125 53524 36159
rect 53472 36116 53524 36125
rect 53748 36159 53800 36168
rect 53748 36125 53757 36159
rect 53757 36125 53791 36159
rect 53791 36125 53800 36159
rect 53748 36116 53800 36125
rect 54576 36116 54628 36168
rect 22652 36091 22704 36100
rect 22652 36057 22661 36091
rect 22661 36057 22695 36091
rect 22695 36057 22704 36091
rect 23480 36091 23532 36100
rect 22652 36048 22704 36057
rect 23480 36057 23489 36091
rect 23489 36057 23523 36091
rect 23523 36057 23532 36091
rect 23480 36048 23532 36057
rect 24032 36091 24084 36100
rect 24032 36057 24041 36091
rect 24041 36057 24075 36091
rect 24075 36057 24084 36091
rect 24032 36048 24084 36057
rect 38568 36048 38620 36100
rect 41696 36048 41748 36100
rect 52828 36048 52880 36100
rect 53656 36091 53708 36100
rect 53656 36057 53665 36091
rect 53665 36057 53699 36091
rect 53699 36057 53708 36091
rect 53656 36048 53708 36057
rect 57980 36091 58032 36100
rect 57980 36057 57989 36091
rect 57989 36057 58023 36091
rect 58023 36057 58032 36091
rect 57980 36048 58032 36057
rect 58348 36091 58400 36100
rect 58348 36057 58357 36091
rect 58357 36057 58391 36091
rect 58391 36057 58400 36091
rect 58348 36048 58400 36057
rect 20168 35980 20220 36032
rect 20720 35980 20772 36032
rect 21548 36023 21600 36032
rect 21548 35989 21557 36023
rect 21557 35989 21591 36023
rect 21591 35989 21600 36023
rect 21548 35980 21600 35989
rect 23664 35980 23716 36032
rect 37280 35980 37332 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 2320 35708 2372 35760
rect 1676 35683 1728 35692
rect 1676 35649 1685 35683
rect 1685 35649 1719 35683
rect 1719 35649 1728 35683
rect 1676 35640 1728 35649
rect 20260 35776 20312 35828
rect 23480 35776 23532 35828
rect 26148 35776 26200 35828
rect 34428 35776 34480 35828
rect 19340 35572 19392 35624
rect 23756 35708 23808 35760
rect 37280 35708 37332 35760
rect 22192 35683 22244 35692
rect 20076 35572 20128 35624
rect 20536 35572 20588 35624
rect 19892 35504 19944 35556
rect 15844 35436 15896 35488
rect 21364 35504 21416 35556
rect 21824 35436 21876 35488
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 24124 35683 24176 35692
rect 24124 35649 24133 35683
rect 24133 35649 24167 35683
rect 24167 35649 24176 35683
rect 24124 35640 24176 35649
rect 33140 35640 33192 35692
rect 23664 35572 23716 35624
rect 36176 35572 36228 35624
rect 40684 35572 40736 35624
rect 35992 35504 36044 35556
rect 22744 35436 22796 35488
rect 23848 35479 23900 35488
rect 23848 35445 23857 35479
rect 23857 35445 23891 35479
rect 23891 35445 23900 35479
rect 23848 35436 23900 35445
rect 23940 35436 23992 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19984 35232 20036 35284
rect 21824 35275 21876 35284
rect 21824 35241 21833 35275
rect 21833 35241 21867 35275
rect 21867 35241 21876 35275
rect 21824 35232 21876 35241
rect 43444 35232 43496 35284
rect 50160 35232 50212 35284
rect 2780 35164 2832 35216
rect 16672 35164 16724 35216
rect 20720 35207 20772 35216
rect 19340 35028 19392 35080
rect 1676 35003 1728 35012
rect 1676 34969 1685 35003
rect 1685 34969 1719 35003
rect 1719 34969 1728 35003
rect 1676 34960 1728 34969
rect 12164 34960 12216 35012
rect 20720 35173 20729 35207
rect 20729 35173 20763 35207
rect 20763 35173 20772 35207
rect 20720 35164 20772 35173
rect 23664 35164 23716 35216
rect 24768 35164 24820 35216
rect 37004 35164 37056 35216
rect 44824 35164 44876 35216
rect 58624 35164 58676 35216
rect 19708 35003 19760 35012
rect 19708 34969 19717 35003
rect 19717 34969 19751 35003
rect 19751 34969 19760 35003
rect 21364 35028 21416 35080
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 22652 35028 22704 35080
rect 24768 35028 24820 35080
rect 35992 35071 36044 35080
rect 19708 34960 19760 34969
rect 21088 34935 21140 34944
rect 21088 34901 21097 34935
rect 21097 34901 21131 34935
rect 21131 34901 21140 34935
rect 21088 34892 21140 34901
rect 26148 34960 26200 35012
rect 22468 34892 22520 34944
rect 35992 35037 36001 35071
rect 36001 35037 36035 35071
rect 36035 35037 36044 35071
rect 35992 35028 36044 35037
rect 36084 35071 36136 35080
rect 36084 35037 36093 35071
rect 36093 35037 36127 35071
rect 36127 35037 36136 35071
rect 36084 35028 36136 35037
rect 36820 35071 36872 35080
rect 36820 35037 36829 35071
rect 36829 35037 36863 35071
rect 36863 35037 36872 35071
rect 36820 35028 36872 35037
rect 40316 35071 40368 35080
rect 37372 34960 37424 35012
rect 40316 35037 40325 35071
rect 40325 35037 40359 35071
rect 40359 35037 40368 35071
rect 40316 35028 40368 35037
rect 40684 35028 40736 35080
rect 47768 35028 47820 35080
rect 40224 35003 40276 35012
rect 40224 34969 40233 35003
rect 40233 34969 40267 35003
rect 40267 34969 40276 35003
rect 40224 34960 40276 34969
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 45100 34892 45152 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 22376 34688 22428 34740
rect 23848 34688 23900 34740
rect 22744 34620 22796 34672
rect 22100 34595 22152 34604
rect 22100 34561 22109 34595
rect 22109 34561 22143 34595
rect 22143 34561 22152 34595
rect 22100 34552 22152 34561
rect 22284 34595 22336 34604
rect 22284 34561 22291 34595
rect 22291 34561 22336 34595
rect 22284 34552 22336 34561
rect 20812 34416 20864 34468
rect 22560 34552 22612 34604
rect 22836 34552 22888 34604
rect 22744 34484 22796 34536
rect 23480 34552 23532 34604
rect 26332 34663 26384 34672
rect 26332 34629 26341 34663
rect 26341 34629 26375 34663
rect 26375 34629 26384 34663
rect 26332 34620 26384 34629
rect 25964 34595 26016 34604
rect 25964 34561 25973 34595
rect 25973 34561 26007 34595
rect 26007 34561 26016 34595
rect 25964 34552 26016 34561
rect 26148 34595 26200 34604
rect 26148 34561 26155 34595
rect 26155 34561 26200 34595
rect 26148 34552 26200 34561
rect 24492 34484 24544 34536
rect 24676 34484 24728 34536
rect 37372 34688 37424 34740
rect 50712 34688 50764 34740
rect 57796 34688 57848 34740
rect 57980 34688 58032 34740
rect 26884 34620 26936 34672
rect 40224 34620 40276 34672
rect 57888 34552 57940 34604
rect 23204 34416 23256 34468
rect 26056 34416 26108 34468
rect 33600 34484 33652 34536
rect 34428 34484 34480 34536
rect 19432 34348 19484 34400
rect 20352 34348 20404 34400
rect 21272 34348 21324 34400
rect 22100 34348 22152 34400
rect 26608 34391 26660 34400
rect 26608 34357 26617 34391
rect 26617 34357 26651 34391
rect 26651 34357 26660 34391
rect 26608 34348 26660 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 20628 33940 20680 33992
rect 31760 34144 31812 34196
rect 21272 33983 21324 33992
rect 21272 33949 21286 33983
rect 21286 33949 21320 33983
rect 21320 33949 21324 33983
rect 22560 34051 22612 34060
rect 22560 34017 22569 34051
rect 22569 34017 22603 34051
rect 22603 34017 22612 34051
rect 22560 34008 22612 34017
rect 21272 33940 21324 33949
rect 22468 33983 22520 33992
rect 22468 33949 22477 33983
rect 22477 33949 22511 33983
rect 22511 33949 22520 33983
rect 22468 33940 22520 33949
rect 35348 33940 35400 33992
rect 1676 33915 1728 33924
rect 1676 33881 1685 33915
rect 1685 33881 1719 33915
rect 1719 33881 1728 33915
rect 1676 33872 1728 33881
rect 20720 33872 20772 33924
rect 35440 33872 35492 33924
rect 35900 33872 35952 33924
rect 57152 33872 57204 33924
rect 22284 33804 22336 33856
rect 49332 33804 49384 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 2136 33532 2188 33584
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 22008 33507 22060 33516
rect 22008 33473 22017 33507
rect 22017 33473 22051 33507
rect 22051 33473 22060 33507
rect 22008 33464 22060 33473
rect 22100 33507 22152 33516
rect 22100 33473 22109 33507
rect 22109 33473 22143 33507
rect 22143 33473 22152 33507
rect 22100 33464 22152 33473
rect 23664 33464 23716 33516
rect 24768 33464 24820 33516
rect 27436 33396 27488 33448
rect 38844 33260 38896 33312
rect 45008 33260 45060 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19432 33056 19484 33108
rect 28356 33056 28408 33108
rect 26608 32988 26660 33040
rect 16948 32920 17000 32972
rect 21088 32920 21140 32972
rect 21640 32920 21692 32972
rect 58164 32963 58216 32972
rect 58164 32929 58173 32963
rect 58173 32929 58207 32963
rect 58207 32929 58216 32963
rect 58164 32920 58216 32929
rect 23664 32852 23716 32904
rect 26700 32895 26752 32904
rect 26700 32861 26709 32895
rect 26709 32861 26743 32895
rect 26743 32861 26752 32895
rect 26700 32852 26752 32861
rect 26976 32895 27028 32904
rect 26976 32861 26985 32895
rect 26985 32861 27019 32895
rect 27019 32861 27028 32895
rect 26976 32852 27028 32861
rect 57704 32852 57756 32904
rect 1676 32827 1728 32836
rect 1676 32793 1685 32827
rect 1685 32793 1719 32827
rect 1719 32793 1728 32827
rect 1676 32784 1728 32793
rect 57060 32827 57112 32836
rect 57060 32793 57069 32827
rect 57069 32793 57103 32827
rect 57103 32793 57112 32827
rect 57060 32784 57112 32793
rect 18144 32716 18196 32768
rect 27160 32759 27212 32768
rect 27160 32725 27169 32759
rect 27169 32725 27203 32759
rect 27203 32725 27212 32759
rect 27160 32716 27212 32725
rect 57152 32759 57204 32768
rect 57152 32725 57161 32759
rect 57161 32725 57195 32759
rect 57195 32725 57204 32759
rect 57152 32716 57204 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 29920 32512 29972 32564
rect 41604 32512 41656 32564
rect 31760 32444 31812 32496
rect 47400 32444 47452 32496
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 15660 32376 15712 32428
rect 24032 32376 24084 32428
rect 26148 32376 26200 32428
rect 53840 32376 53892 32428
rect 25320 32172 25372 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 21824 31968 21876 32020
rect 23020 31968 23072 32020
rect 26056 31968 26108 32020
rect 25504 31900 25556 31952
rect 25964 31900 26016 31952
rect 58440 31900 58492 31952
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 44364 31832 44416 31884
rect 26056 31764 26108 31816
rect 57796 31832 57848 31884
rect 22928 31696 22980 31748
rect 25780 31696 25832 31748
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 19524 31356 19576 31408
rect 25596 31399 25648 31408
rect 25596 31365 25605 31399
rect 25605 31365 25639 31399
rect 25639 31365 25648 31399
rect 25596 31356 25648 31365
rect 26700 31424 26752 31476
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 19432 31288 19484 31340
rect 18236 31220 18288 31272
rect 22652 31288 22704 31340
rect 25228 31288 25280 31340
rect 20076 31263 20128 31272
rect 20076 31229 20085 31263
rect 20085 31229 20119 31263
rect 20119 31229 20128 31263
rect 20076 31220 20128 31229
rect 25780 31331 25832 31340
rect 25780 31297 25794 31331
rect 25794 31297 25828 31331
rect 25828 31297 25832 31331
rect 25780 31288 25832 31297
rect 46940 31288 46992 31340
rect 58072 31331 58124 31340
rect 58072 31297 58081 31331
rect 58081 31297 58115 31331
rect 58115 31297 58124 31331
rect 58072 31288 58124 31297
rect 19708 31195 19760 31204
rect 19708 31161 19717 31195
rect 19717 31161 19751 31195
rect 19751 31161 19760 31195
rect 19708 31152 19760 31161
rect 27712 31152 27764 31204
rect 57152 31152 57204 31204
rect 1768 31127 1820 31136
rect 1768 31093 1777 31127
rect 1777 31093 1811 31127
rect 1811 31093 1820 31127
rect 1768 31084 1820 31093
rect 19432 31084 19484 31136
rect 22652 31084 22704 31136
rect 28264 31084 28316 31136
rect 40960 31084 41012 31136
rect 46480 31084 46532 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1768 30880 1820 30932
rect 19524 30880 19576 30932
rect 19708 30880 19760 30932
rect 25320 30880 25372 30932
rect 25596 30880 25648 30932
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 19616 30719 19668 30728
rect 19616 30685 19623 30719
rect 19623 30685 19668 30719
rect 19616 30676 19668 30685
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 19984 30812 20036 30864
rect 20168 30812 20220 30864
rect 20352 30676 20404 30728
rect 22928 30676 22980 30728
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 22836 30336 22888 30388
rect 24216 30336 24268 30388
rect 5724 30268 5776 30320
rect 17960 30200 18012 30252
rect 23940 30268 23992 30320
rect 24032 30268 24084 30320
rect 24676 30268 24728 30320
rect 25320 30311 25372 30320
rect 25320 30277 25329 30311
rect 25329 30277 25363 30311
rect 25363 30277 25372 30311
rect 25320 30268 25372 30277
rect 24492 30200 24544 30252
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 1768 30175 1820 30184
rect 1768 30141 1777 30175
rect 1777 30141 1811 30175
rect 1811 30141 1820 30175
rect 1768 30132 1820 30141
rect 4068 30132 4120 30184
rect 23664 30132 23716 30184
rect 25688 30132 25740 30184
rect 46388 30200 46440 30252
rect 26332 30064 26384 30116
rect 44732 30132 44784 30184
rect 24308 29996 24360 30048
rect 24768 29996 24820 30048
rect 25136 29996 25188 30048
rect 25872 29996 25924 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 22652 29792 22704 29844
rect 23480 29792 23532 29844
rect 25872 29835 25924 29844
rect 25872 29801 25881 29835
rect 25881 29801 25915 29835
rect 25915 29801 25924 29835
rect 25872 29792 25924 29801
rect 25964 29835 26016 29844
rect 25964 29801 25973 29835
rect 25973 29801 26007 29835
rect 26007 29801 26016 29835
rect 25964 29792 26016 29801
rect 20168 29724 20220 29776
rect 23940 29724 23992 29776
rect 24032 29767 24084 29776
rect 24032 29733 24041 29767
rect 24041 29733 24075 29767
rect 24075 29733 24084 29767
rect 24032 29724 24084 29733
rect 24492 29724 24544 29776
rect 18696 29656 18748 29708
rect 16396 29588 16448 29640
rect 23480 29631 23532 29640
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 23848 29631 23900 29640
rect 23848 29597 23857 29631
rect 23857 29597 23891 29631
rect 23891 29597 23900 29631
rect 23848 29588 23900 29597
rect 24584 29631 24636 29640
rect 24584 29597 24593 29631
rect 24593 29597 24627 29631
rect 24627 29597 24636 29631
rect 24584 29588 24636 29597
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25136 29656 25188 29708
rect 25964 29588 26016 29640
rect 26148 29631 26200 29640
rect 26148 29597 26157 29631
rect 26157 29597 26191 29631
rect 26191 29597 26200 29631
rect 58164 29699 58216 29708
rect 58164 29665 58173 29699
rect 58173 29665 58207 29699
rect 58207 29665 58216 29699
rect 58164 29656 58216 29665
rect 26148 29588 26200 29597
rect 57796 29588 57848 29640
rect 1860 29563 1912 29572
rect 1860 29529 1869 29563
rect 1869 29529 1903 29563
rect 1903 29529 1912 29563
rect 1860 29520 1912 29529
rect 23204 29520 23256 29572
rect 24400 29520 24452 29572
rect 24676 29520 24728 29572
rect 20076 29452 20128 29504
rect 25320 29520 25372 29572
rect 57060 29563 57112 29572
rect 57060 29529 57069 29563
rect 57069 29529 57103 29563
rect 57103 29529 57112 29563
rect 57060 29520 57112 29529
rect 25136 29495 25188 29504
rect 25136 29461 25145 29495
rect 25145 29461 25179 29495
rect 25179 29461 25188 29495
rect 25136 29452 25188 29461
rect 25596 29495 25648 29504
rect 25596 29461 25605 29495
rect 25605 29461 25639 29495
rect 25639 29461 25648 29495
rect 25596 29452 25648 29461
rect 30932 29452 30984 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 23480 29248 23532 29300
rect 48780 29248 48832 29300
rect 17960 29223 18012 29232
rect 17960 29189 17969 29223
rect 17969 29189 18003 29223
rect 18003 29189 18012 29223
rect 17960 29180 18012 29189
rect 24308 29223 24360 29232
rect 24308 29189 24317 29223
rect 24317 29189 24351 29223
rect 24351 29189 24360 29223
rect 24308 29180 24360 29189
rect 25136 29180 25188 29232
rect 17684 29112 17736 29164
rect 18144 29112 18196 29164
rect 20168 29112 20220 29164
rect 23572 29112 23624 29164
rect 25596 29155 25648 29164
rect 25596 29121 25605 29155
rect 25605 29121 25639 29155
rect 25639 29121 25648 29155
rect 25596 29112 25648 29121
rect 24032 29044 24084 29096
rect 25320 29044 25372 29096
rect 25412 29044 25464 29096
rect 26976 29044 27028 29096
rect 24492 28908 24544 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 50988 28500 51040 28552
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 18328 28432 18380 28484
rect 39488 28432 39540 28484
rect 58164 28475 58216 28484
rect 58164 28441 58173 28475
rect 58173 28441 58207 28475
rect 58207 28441 58216 28475
rect 58164 28432 58216 28441
rect 7656 28364 7708 28416
rect 20168 28364 20220 28416
rect 24584 28364 24636 28416
rect 54760 28364 54812 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 1584 28160 1636 28212
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 4988 28024 5040 28076
rect 58072 28067 58124 28076
rect 58072 28033 58081 28067
rect 58081 28033 58115 28067
rect 58115 28033 58124 28067
rect 58072 28024 58124 28033
rect 1768 27999 1820 28008
rect 1768 27965 1777 27999
rect 1777 27965 1811 27999
rect 1811 27965 1820 27999
rect 1768 27956 1820 27965
rect 14464 27888 14516 27940
rect 32772 27820 32824 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 1860 27387 1912 27396
rect 1860 27353 1869 27387
rect 1869 27353 1903 27387
rect 1903 27353 1912 27387
rect 1860 27344 1912 27353
rect 3240 27344 3292 27396
rect 9588 27344 9640 27396
rect 24124 27276 24176 27328
rect 25412 27276 25464 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1584 27072 1636 27124
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 2688 26979 2740 26988
rect 2688 26945 2701 26979
rect 2701 26945 2740 26979
rect 2688 26936 2740 26945
rect 18052 26936 18104 26988
rect 29552 26936 29604 26988
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 6184 26868 6236 26920
rect 20996 26868 21048 26920
rect 23296 26868 23348 26920
rect 55680 26868 55732 26920
rect 15200 26800 15252 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 45652 26324 45704 26376
rect 26332 26256 26384 26308
rect 57060 26299 57112 26308
rect 57060 26265 57069 26299
rect 57069 26265 57103 26299
rect 57103 26265 57112 26299
rect 57060 26256 57112 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 17684 25848 17736 25900
rect 20444 25848 20496 25900
rect 32496 25848 32548 25900
rect 1768 25823 1820 25832
rect 1768 25789 1777 25823
rect 1777 25789 1811 25823
rect 1811 25789 1820 25823
rect 1768 25780 1820 25789
rect 21824 25780 21876 25832
rect 29828 25712 29880 25764
rect 42432 25712 42484 25764
rect 5172 25644 5224 25696
rect 18512 25644 18564 25696
rect 26148 25644 26200 25696
rect 43536 25644 43588 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 2688 25279 2740 25288
rect 2688 25245 2701 25279
rect 2701 25245 2740 25279
rect 2688 25236 2740 25245
rect 39948 25236 40000 25288
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 58164 25211 58216 25220
rect 58164 25177 58173 25211
rect 58173 25177 58207 25211
rect 58207 25177 58216 25211
rect 58164 25168 58216 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 46756 24828 46808 24880
rect 49056 24828 49108 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 58072 24803 58124 24812
rect 58072 24769 58081 24803
rect 58081 24769 58115 24803
rect 58115 24769 58124 24803
rect 58072 24760 58124 24769
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 2688 24692 2740 24744
rect 18696 24692 18748 24744
rect 37924 24556 37976 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24352 1636 24404
rect 6920 24284 6972 24336
rect 40776 24284 40828 24336
rect 50160 24284 50212 24336
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 6920 24148 6972 24200
rect 18420 24216 18472 24268
rect 24952 24216 25004 24268
rect 47584 24216 47636 24268
rect 17224 24148 17276 24200
rect 19984 24148 20036 24200
rect 54024 24148 54076 24200
rect 16856 24080 16908 24132
rect 20260 24080 20312 24132
rect 55220 24080 55272 24132
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 17224 23851 17276 23860
rect 17224 23817 17233 23851
rect 17233 23817 17267 23851
rect 17267 23817 17276 23851
rect 17224 23808 17276 23817
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 18972 23672 19024 23724
rect 17684 23604 17736 23656
rect 15200 23536 15252 23588
rect 18328 23536 18380 23588
rect 18420 23468 18472 23520
rect 20536 23468 20588 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 22284 23264 22336 23316
rect 41144 23264 41196 23316
rect 46480 23264 46532 23316
rect 23020 23196 23072 23248
rect 23296 23196 23348 23248
rect 24400 23196 24452 23248
rect 27620 23128 27672 23180
rect 58164 23171 58216 23180
rect 58164 23137 58173 23171
rect 58173 23137 58207 23171
rect 58207 23137 58216 23171
rect 58164 23128 58216 23137
rect 17684 23060 17736 23112
rect 19340 23060 19392 23112
rect 20076 23060 20128 23112
rect 24676 23060 24728 23112
rect 26608 23103 26660 23112
rect 26608 23069 26617 23103
rect 26617 23069 26651 23103
rect 26651 23069 26660 23103
rect 26608 23060 26660 23069
rect 57612 23060 57664 23112
rect 1860 23035 1912 23044
rect 1860 23001 1869 23035
rect 1869 23001 1903 23035
rect 1903 23001 1912 23035
rect 1860 22992 1912 23001
rect 22468 22992 22520 23044
rect 25504 22992 25556 23044
rect 24584 22924 24636 22976
rect 32588 22924 32640 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 30656 22720 30708 22772
rect 42524 22720 42576 22772
rect 27804 22652 27856 22704
rect 22836 22627 22888 22636
rect 22836 22593 22845 22627
rect 22845 22593 22879 22627
rect 22879 22593 22888 22627
rect 22836 22584 22888 22593
rect 25780 22584 25832 22636
rect 58072 22627 58124 22636
rect 58072 22593 58081 22627
rect 58081 22593 58115 22627
rect 58115 22593 58124 22627
rect 58072 22584 58124 22593
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 17684 22516 17736 22568
rect 23296 22516 23348 22568
rect 27620 22516 27672 22568
rect 28448 22516 28500 22568
rect 25872 22491 25924 22500
rect 25872 22457 25881 22491
rect 25881 22457 25915 22491
rect 25915 22457 25924 22491
rect 25872 22448 25924 22457
rect 22100 22380 22152 22432
rect 26056 22423 26108 22432
rect 26056 22389 26065 22423
rect 26065 22389 26099 22423
rect 26099 22389 26108 22423
rect 26056 22380 26108 22389
rect 27528 22423 27580 22432
rect 27528 22389 27537 22423
rect 27537 22389 27571 22423
rect 27571 22389 27580 22423
rect 27528 22380 27580 22389
rect 32956 22380 33008 22432
rect 34428 22380 34480 22432
rect 38476 22380 38528 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 23572 22176 23624 22228
rect 26516 22176 26568 22228
rect 21732 22108 21784 22160
rect 27436 22108 27488 22160
rect 16120 22040 16172 22092
rect 22468 22083 22520 22092
rect 22468 22049 22477 22083
rect 22477 22049 22511 22083
rect 22511 22049 22520 22083
rect 22468 22040 22520 22049
rect 26424 22040 26476 22092
rect 17684 21972 17736 22024
rect 24584 22015 24636 22024
rect 1860 21947 1912 21956
rect 1860 21913 1869 21947
rect 1869 21913 1903 21947
rect 1903 21913 1912 21947
rect 1860 21904 1912 21913
rect 23020 21904 23072 21956
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 23756 21904 23808 21956
rect 23940 21904 23992 21956
rect 27896 21972 27948 22024
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 55864 21972 55916 22024
rect 20352 21836 20404 21888
rect 27712 21836 27764 21888
rect 41328 21904 41380 21956
rect 58164 21947 58216 21956
rect 58164 21913 58173 21947
rect 58173 21913 58207 21947
rect 58207 21913 58216 21947
rect 58164 21904 58216 21913
rect 28724 21879 28776 21888
rect 28724 21845 28733 21879
rect 28733 21845 28767 21879
rect 28767 21845 28776 21879
rect 28724 21836 28776 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 22836 21632 22888 21684
rect 20904 21607 20956 21616
rect 20904 21573 20913 21607
rect 20913 21573 20947 21607
rect 20947 21573 20956 21607
rect 20904 21564 20956 21573
rect 21180 21564 21232 21616
rect 25872 21632 25924 21684
rect 27712 21632 27764 21684
rect 28172 21632 28224 21684
rect 8208 21496 8260 21548
rect 22652 21496 22704 21548
rect 23020 21496 23072 21548
rect 24124 21496 24176 21548
rect 27528 21564 27580 21616
rect 25596 21496 25648 21548
rect 28724 21496 28776 21548
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 58072 21539 58124 21548
rect 58072 21505 58081 21539
rect 58081 21505 58115 21539
rect 58115 21505 58124 21539
rect 58072 21496 58124 21505
rect 20628 21428 20680 21480
rect 22468 21428 22520 21480
rect 23112 21428 23164 21480
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 21088 21335 21140 21344
rect 21088 21301 21097 21335
rect 21097 21301 21131 21335
rect 21131 21301 21140 21335
rect 21088 21292 21140 21301
rect 21272 21335 21324 21344
rect 21272 21301 21281 21335
rect 21281 21301 21315 21335
rect 21315 21301 21324 21335
rect 21272 21292 21324 21301
rect 26240 21428 26292 21480
rect 23756 21292 23808 21344
rect 26700 21292 26752 21344
rect 28448 21428 28500 21480
rect 28816 21428 28868 21480
rect 28540 21360 28592 21412
rect 28448 21292 28500 21344
rect 29000 21292 29052 21344
rect 40040 21360 40092 21412
rect 42064 21360 42116 21412
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 22008 21088 22060 21140
rect 27344 21088 27396 21140
rect 19248 21020 19300 21072
rect 27160 21020 27212 21072
rect 23388 20952 23440 21004
rect 24676 20952 24728 21004
rect 28908 20952 28960 21004
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 16672 20816 16724 20868
rect 21272 20884 21324 20936
rect 22100 20884 22152 20936
rect 26056 20884 26108 20936
rect 45100 20884 45152 20936
rect 46020 20884 46072 20936
rect 20720 20816 20772 20868
rect 32404 20816 32456 20868
rect 33784 20816 33836 20868
rect 44272 20816 44324 20868
rect 47768 20816 47820 20868
rect 20536 20748 20588 20800
rect 20812 20748 20864 20800
rect 21272 20748 21324 20800
rect 22928 20791 22980 20800
rect 22928 20757 22937 20791
rect 22937 20757 22971 20791
rect 22971 20757 22980 20791
rect 22928 20748 22980 20757
rect 27252 20748 27304 20800
rect 27896 20748 27948 20800
rect 28264 20748 28316 20800
rect 30104 20791 30156 20800
rect 30104 20757 30113 20791
rect 30113 20757 30147 20791
rect 30147 20757 30156 20791
rect 30104 20748 30156 20757
rect 31392 20748 31444 20800
rect 58348 20748 58400 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 20628 20544 20680 20596
rect 20720 20544 20772 20596
rect 14280 20408 14332 20460
rect 18788 20408 18840 20460
rect 19984 20476 20036 20528
rect 19524 20451 19576 20460
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 19524 20417 19533 20451
rect 19533 20417 19567 20451
rect 19567 20417 19576 20451
rect 19524 20408 19576 20417
rect 20260 20451 20312 20460
rect 20260 20417 20294 20451
rect 20294 20417 20312 20451
rect 20260 20408 20312 20417
rect 19432 20340 19484 20392
rect 21272 20544 21324 20596
rect 26424 20587 26476 20596
rect 26424 20553 26433 20587
rect 26433 20553 26467 20587
rect 26467 20553 26476 20587
rect 26424 20544 26476 20553
rect 22100 20476 22152 20528
rect 24124 20476 24176 20528
rect 33508 20544 33560 20596
rect 21916 20408 21968 20460
rect 23572 20451 23624 20460
rect 23572 20417 23581 20451
rect 23581 20417 23615 20451
rect 23615 20417 23624 20451
rect 23572 20408 23624 20417
rect 24584 20408 24636 20460
rect 29736 20476 29788 20528
rect 23480 20340 23532 20392
rect 25136 20340 25188 20392
rect 26700 20408 26752 20460
rect 27436 20408 27488 20460
rect 28448 20451 28500 20460
rect 28448 20417 28457 20451
rect 28457 20417 28491 20451
rect 28491 20417 28500 20451
rect 28448 20408 28500 20417
rect 29000 20408 29052 20460
rect 30656 20451 30708 20460
rect 30656 20417 30679 20451
rect 30679 20417 30708 20451
rect 30656 20408 30708 20417
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 38752 20451 38804 20460
rect 38752 20417 38761 20451
rect 38761 20417 38795 20451
rect 38795 20417 38804 20451
rect 38752 20408 38804 20417
rect 18972 20272 19024 20324
rect 19892 20272 19944 20324
rect 22376 20272 22428 20324
rect 16580 20204 16632 20256
rect 19708 20204 19760 20256
rect 20720 20204 20772 20256
rect 23112 20204 23164 20256
rect 24584 20204 24636 20256
rect 24768 20247 24820 20256
rect 24768 20213 24777 20247
rect 24777 20213 24811 20247
rect 24811 20213 24820 20247
rect 24768 20204 24820 20213
rect 26240 20272 26292 20324
rect 27896 20272 27948 20324
rect 26884 20204 26936 20256
rect 27804 20204 27856 20256
rect 28724 20204 28776 20256
rect 38384 20340 38436 20392
rect 39212 20340 39264 20392
rect 57980 20340 58032 20392
rect 36268 20272 36320 20324
rect 39120 20272 39172 20324
rect 39764 20272 39816 20324
rect 29828 20247 29880 20256
rect 29828 20213 29837 20247
rect 29837 20213 29871 20247
rect 29871 20213 29880 20247
rect 29828 20204 29880 20213
rect 30104 20204 30156 20256
rect 31852 20204 31904 20256
rect 39028 20204 39080 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4068 19796 4120 19848
rect 15016 19796 15068 19848
rect 18052 19796 18104 19848
rect 19708 20000 19760 20052
rect 18604 19975 18656 19984
rect 18604 19941 18613 19975
rect 18613 19941 18647 19975
rect 18647 19941 18656 19975
rect 18604 19932 18656 19941
rect 20904 20000 20956 20052
rect 24124 20000 24176 20052
rect 24584 20000 24636 20052
rect 25228 20000 25280 20052
rect 30380 20000 30432 20052
rect 24860 19864 24912 19916
rect 18972 19796 19024 19848
rect 19432 19796 19484 19848
rect 19892 19796 19944 19848
rect 21180 19796 21232 19848
rect 24676 19796 24728 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 25136 19864 25188 19916
rect 25688 19864 25740 19916
rect 38752 20000 38804 20052
rect 40224 20000 40276 20052
rect 41144 20000 41196 20052
rect 48136 20000 48188 20052
rect 48964 20000 49016 20052
rect 47860 19932 47912 19984
rect 24768 19796 24820 19805
rect 26056 19796 26108 19848
rect 30104 19839 30156 19848
rect 30104 19805 30113 19839
rect 30113 19805 30147 19839
rect 30147 19805 30156 19839
rect 30104 19796 30156 19805
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 17316 19728 17368 19780
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 18512 19728 18564 19780
rect 22468 19728 22520 19780
rect 24584 19771 24636 19780
rect 24584 19737 24593 19771
rect 24593 19737 24627 19771
rect 24627 19737 24636 19771
rect 24584 19728 24636 19737
rect 30564 19864 30616 19916
rect 33048 19796 33100 19848
rect 36268 19796 36320 19848
rect 37464 19796 37516 19848
rect 39212 19796 39264 19848
rect 39764 19864 39816 19916
rect 40316 19796 40368 19848
rect 41420 19864 41472 19916
rect 48872 19864 48924 19916
rect 58164 19907 58216 19916
rect 58164 19873 58173 19907
rect 58173 19873 58207 19907
rect 58207 19873 58216 19907
rect 58164 19864 58216 19873
rect 40868 19796 40920 19848
rect 48596 19796 48648 19848
rect 19064 19660 19116 19712
rect 19524 19660 19576 19712
rect 26792 19660 26844 19712
rect 27620 19660 27672 19712
rect 28816 19660 28868 19712
rect 30288 19703 30340 19712
rect 30288 19669 30297 19703
rect 30297 19669 30331 19703
rect 30331 19669 30340 19703
rect 30288 19660 30340 19669
rect 37372 19728 37424 19780
rect 37740 19728 37792 19780
rect 30840 19660 30892 19712
rect 35532 19660 35584 19712
rect 36452 19660 36504 19712
rect 36820 19703 36872 19712
rect 36820 19669 36829 19703
rect 36829 19669 36863 19703
rect 36863 19669 36872 19703
rect 36820 19660 36872 19669
rect 38844 19660 38896 19712
rect 40776 19660 40828 19712
rect 48504 19703 48556 19712
rect 48504 19669 48513 19703
rect 48513 19669 48547 19703
rect 48547 19669 48556 19703
rect 48504 19660 48556 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 19248 19456 19300 19508
rect 20260 19456 20312 19508
rect 23756 19499 23808 19508
rect 18512 19320 18564 19372
rect 19064 19252 19116 19304
rect 21088 19320 21140 19372
rect 21456 19320 21508 19372
rect 21640 19320 21692 19372
rect 19432 19252 19484 19304
rect 23756 19465 23765 19499
rect 23765 19465 23799 19499
rect 23799 19465 23808 19499
rect 23756 19456 23808 19465
rect 25504 19499 25556 19508
rect 25504 19465 25513 19499
rect 25513 19465 25547 19499
rect 25547 19465 25556 19499
rect 25504 19456 25556 19465
rect 27712 19456 27764 19508
rect 22744 19388 22796 19440
rect 23388 19388 23440 19440
rect 27620 19431 27672 19440
rect 27620 19397 27629 19431
rect 27629 19397 27663 19431
rect 27663 19397 27672 19431
rect 27620 19388 27672 19397
rect 22928 19320 22980 19372
rect 26148 19320 26200 19372
rect 27436 19320 27488 19372
rect 33508 19499 33560 19508
rect 33508 19465 33517 19499
rect 33517 19465 33551 19499
rect 33551 19465 33560 19499
rect 33508 19456 33560 19465
rect 35072 19499 35124 19508
rect 35072 19465 35081 19499
rect 35081 19465 35115 19499
rect 35115 19465 35124 19499
rect 35072 19456 35124 19465
rect 34796 19388 34848 19440
rect 30196 19320 30248 19372
rect 40868 19456 40920 19508
rect 35808 19388 35860 19440
rect 41236 19456 41288 19508
rect 41696 19456 41748 19508
rect 48228 19456 48280 19508
rect 48964 19456 49016 19508
rect 18512 19184 18564 19236
rect 19984 19184 20036 19236
rect 20076 19184 20128 19236
rect 7564 19116 7616 19168
rect 20628 19116 20680 19168
rect 22376 19184 22428 19236
rect 24308 19184 24360 19236
rect 27620 19184 27672 19236
rect 31576 19252 31628 19304
rect 35532 19295 35584 19304
rect 35532 19261 35541 19295
rect 35541 19261 35575 19295
rect 35575 19261 35584 19295
rect 35716 19295 35768 19304
rect 35532 19252 35584 19261
rect 35716 19261 35725 19295
rect 35725 19261 35759 19295
rect 35759 19261 35768 19295
rect 35716 19252 35768 19261
rect 27988 19184 28040 19236
rect 28356 19184 28408 19236
rect 36268 19295 36320 19304
rect 36268 19261 36277 19295
rect 36277 19261 36311 19295
rect 36311 19261 36320 19295
rect 36268 19252 36320 19261
rect 47768 19388 47820 19440
rect 48136 19431 48188 19440
rect 48136 19397 48145 19431
rect 48145 19397 48179 19431
rect 48179 19397 48188 19431
rect 48136 19388 48188 19397
rect 48688 19388 48740 19440
rect 58164 19388 58216 19440
rect 37372 19320 37424 19372
rect 37096 19252 37148 19304
rect 40684 19252 40736 19304
rect 28080 19116 28132 19168
rect 33140 19116 33192 19168
rect 40592 19184 40644 19236
rect 41052 19252 41104 19304
rect 41420 19320 41472 19372
rect 43904 19320 43956 19372
rect 47860 19363 47912 19372
rect 47860 19329 47869 19363
rect 47869 19329 47903 19363
rect 47903 19329 47912 19363
rect 47860 19320 47912 19329
rect 48044 19363 48096 19372
rect 48044 19329 48053 19363
rect 48053 19329 48087 19363
rect 48087 19329 48096 19363
rect 48044 19320 48096 19329
rect 48872 19363 48924 19372
rect 41236 19252 41288 19304
rect 46112 19252 46164 19304
rect 48872 19329 48881 19363
rect 48881 19329 48915 19363
rect 48915 19329 48924 19363
rect 48872 19320 48924 19329
rect 49056 19363 49108 19372
rect 49056 19329 49065 19363
rect 49065 19329 49099 19363
rect 49099 19329 49108 19363
rect 49056 19320 49108 19329
rect 58072 19363 58124 19372
rect 58072 19329 58081 19363
rect 58081 19329 58115 19363
rect 58115 19329 58124 19363
rect 58072 19320 58124 19329
rect 49148 19252 49200 19304
rect 41880 19184 41932 19236
rect 48136 19184 48188 19236
rect 58256 19184 58308 19236
rect 36636 19159 36688 19168
rect 36636 19125 36645 19159
rect 36645 19125 36679 19159
rect 36679 19125 36688 19159
rect 36636 19116 36688 19125
rect 40132 19116 40184 19168
rect 41052 19116 41104 19168
rect 41236 19116 41288 19168
rect 42984 19159 43036 19168
rect 42984 19125 42993 19159
rect 42993 19125 43027 19159
rect 43027 19125 43036 19159
rect 42984 19116 43036 19125
rect 48596 19116 48648 19168
rect 49240 19159 49292 19168
rect 49240 19125 49249 19159
rect 49249 19125 49283 19159
rect 49283 19125 49292 19159
rect 49240 19116 49292 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 15936 18776 15988 18828
rect 17592 18819 17644 18828
rect 16672 18751 16724 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 16764 18708 16816 18760
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 17868 18819 17920 18828
rect 17868 18785 17877 18819
rect 17877 18785 17911 18819
rect 17911 18785 17920 18819
rect 17868 18776 17920 18785
rect 18512 18819 18564 18828
rect 18512 18785 18521 18819
rect 18521 18785 18555 18819
rect 18555 18785 18564 18819
rect 18512 18776 18564 18785
rect 22008 18912 22060 18964
rect 22468 18912 22520 18964
rect 23112 18912 23164 18964
rect 24308 18912 24360 18964
rect 26056 18912 26108 18964
rect 27620 18912 27672 18964
rect 30012 18912 30064 18964
rect 30196 18912 30248 18964
rect 34428 18912 34480 18964
rect 35808 18912 35860 18964
rect 26424 18844 26476 18896
rect 28356 18844 28408 18896
rect 39396 18844 39448 18896
rect 40132 18887 40184 18896
rect 40132 18853 40141 18887
rect 40141 18853 40175 18887
rect 40175 18853 40184 18887
rect 40132 18844 40184 18853
rect 41880 18887 41932 18896
rect 41880 18853 41889 18887
rect 41889 18853 41923 18887
rect 41923 18853 41932 18887
rect 41880 18844 41932 18853
rect 44088 18844 44140 18896
rect 17316 18708 17368 18760
rect 18420 18708 18472 18760
rect 19432 18708 19484 18760
rect 19984 18640 20036 18692
rect 20352 18640 20404 18692
rect 20536 18708 20588 18760
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 23388 18776 23440 18828
rect 26056 18776 26108 18828
rect 24860 18751 24912 18760
rect 24860 18717 24894 18751
rect 24894 18717 24912 18751
rect 24860 18708 24912 18717
rect 26884 18751 26936 18760
rect 26884 18717 26893 18751
rect 26893 18717 26927 18751
rect 26927 18717 26936 18751
rect 26884 18708 26936 18717
rect 28448 18708 28500 18760
rect 29828 18708 29880 18760
rect 33048 18776 33100 18828
rect 38108 18776 38160 18828
rect 34796 18708 34848 18760
rect 34888 18751 34940 18760
rect 34888 18717 34897 18751
rect 34897 18717 34931 18751
rect 34931 18717 34940 18751
rect 34888 18708 34940 18717
rect 35808 18751 35860 18760
rect 18236 18572 18288 18624
rect 21088 18572 21140 18624
rect 21272 18572 21324 18624
rect 23112 18572 23164 18624
rect 27620 18640 27672 18692
rect 30012 18640 30064 18692
rect 24584 18572 24636 18624
rect 26056 18572 26108 18624
rect 26240 18572 26292 18624
rect 30840 18683 30892 18692
rect 30840 18649 30849 18683
rect 30849 18649 30883 18683
rect 30883 18649 30892 18683
rect 30840 18640 30892 18649
rect 33968 18640 34020 18692
rect 34704 18640 34756 18692
rect 35808 18717 35817 18751
rect 35817 18717 35851 18751
rect 35851 18717 35860 18751
rect 35808 18708 35860 18717
rect 38844 18708 38896 18760
rect 39212 18708 39264 18760
rect 40592 18708 40644 18760
rect 40776 18751 40828 18760
rect 40776 18717 40810 18751
rect 40810 18717 40828 18751
rect 40776 18708 40828 18717
rect 42984 18819 43036 18828
rect 42984 18785 42993 18819
rect 42993 18785 43027 18819
rect 43027 18785 43036 18819
rect 42984 18776 43036 18785
rect 43628 18751 43680 18760
rect 43628 18717 43637 18751
rect 43637 18717 43671 18751
rect 43671 18717 43680 18751
rect 43628 18708 43680 18717
rect 43996 18751 44048 18760
rect 43996 18717 44005 18751
rect 44005 18717 44039 18751
rect 44039 18717 44048 18751
rect 43996 18708 44048 18717
rect 45560 18751 45612 18760
rect 40684 18640 40736 18692
rect 43076 18640 43128 18692
rect 44272 18640 44324 18692
rect 45560 18717 45569 18751
rect 45569 18717 45603 18751
rect 45603 18717 45612 18751
rect 45560 18708 45612 18717
rect 49056 18912 49108 18964
rect 48044 18844 48096 18896
rect 46112 18776 46164 18828
rect 48596 18776 48648 18828
rect 48228 18751 48280 18760
rect 48228 18717 48237 18751
rect 48237 18717 48271 18751
rect 48271 18717 48280 18751
rect 48228 18708 48280 18717
rect 48688 18708 48740 18760
rect 49148 18776 49200 18828
rect 57888 18751 57940 18760
rect 57888 18717 57897 18751
rect 57897 18717 57931 18751
rect 57931 18717 57940 18751
rect 57888 18708 57940 18717
rect 46848 18640 46900 18692
rect 48044 18683 48096 18692
rect 48044 18649 48053 18683
rect 48053 18649 48087 18683
rect 48087 18649 48096 18683
rect 48044 18640 48096 18649
rect 48136 18683 48188 18692
rect 48136 18649 48145 18683
rect 48145 18649 48179 18683
rect 48179 18649 48188 18683
rect 48136 18640 48188 18649
rect 49884 18640 49936 18692
rect 50712 18640 50764 18692
rect 58164 18683 58216 18692
rect 58164 18649 58173 18683
rect 58173 18649 58207 18683
rect 58207 18649 58216 18683
rect 58164 18640 58216 18649
rect 30748 18615 30800 18624
rect 30748 18581 30757 18615
rect 30757 18581 30791 18615
rect 30791 18581 30800 18615
rect 30748 18572 30800 18581
rect 34520 18572 34572 18624
rect 38568 18615 38620 18624
rect 38568 18581 38577 18615
rect 38577 18581 38611 18615
rect 38611 18581 38620 18615
rect 38568 18572 38620 18581
rect 39212 18572 39264 18624
rect 42984 18572 43036 18624
rect 45744 18615 45796 18624
rect 45744 18581 45753 18615
rect 45753 18581 45787 18615
rect 45787 18581 45796 18615
rect 45744 18572 45796 18581
rect 45928 18572 45980 18624
rect 48688 18572 48740 18624
rect 49424 18615 49476 18624
rect 49424 18581 49433 18615
rect 49433 18581 49467 18615
rect 49467 18581 49476 18615
rect 49424 18572 49476 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 7564 18368 7616 18420
rect 17132 18368 17184 18420
rect 17500 18368 17552 18420
rect 18512 18368 18564 18420
rect 24308 18368 24360 18420
rect 24400 18368 24452 18420
rect 27068 18368 27120 18420
rect 27896 18368 27948 18420
rect 31392 18411 31444 18420
rect 31392 18377 31401 18411
rect 31401 18377 31435 18411
rect 31435 18377 31444 18411
rect 31392 18368 31444 18377
rect 34796 18368 34848 18420
rect 37188 18368 37240 18420
rect 37464 18411 37516 18420
rect 37464 18377 37473 18411
rect 37473 18377 37507 18411
rect 37507 18377 37516 18411
rect 37464 18368 37516 18377
rect 38844 18368 38896 18420
rect 17868 18300 17920 18352
rect 14188 18232 14240 18284
rect 15752 18232 15804 18284
rect 19984 18300 20036 18352
rect 21272 18300 21324 18352
rect 24032 18300 24084 18352
rect 25872 18300 25924 18352
rect 26424 18300 26476 18352
rect 27528 18300 27580 18352
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 21088 18232 21140 18284
rect 13728 18096 13780 18148
rect 10784 18028 10836 18080
rect 18512 18096 18564 18148
rect 20536 18096 20588 18148
rect 26056 18164 26108 18216
rect 27160 18232 27212 18284
rect 27620 18275 27672 18284
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 27896 18232 27948 18284
rect 28264 18275 28316 18284
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 29828 18232 29880 18284
rect 30656 18232 30708 18284
rect 36636 18300 36688 18352
rect 43628 18368 43680 18420
rect 44272 18411 44324 18420
rect 44272 18377 44281 18411
rect 44281 18377 44315 18411
rect 44315 18377 44324 18411
rect 44272 18368 44324 18377
rect 37280 18232 37332 18284
rect 22192 18139 22244 18148
rect 22192 18105 22201 18139
rect 22201 18105 22235 18139
rect 22235 18105 22244 18139
rect 22192 18096 22244 18105
rect 24032 18096 24084 18148
rect 24676 18096 24728 18148
rect 26148 18096 26200 18148
rect 23756 18028 23808 18080
rect 26884 18028 26936 18080
rect 27436 18164 27488 18216
rect 30472 18164 30524 18216
rect 31116 18164 31168 18216
rect 31576 18207 31628 18216
rect 31576 18173 31585 18207
rect 31585 18173 31619 18207
rect 31619 18173 31628 18207
rect 31576 18164 31628 18173
rect 34244 18164 34296 18216
rect 37924 18207 37976 18216
rect 37924 18173 37933 18207
rect 37933 18173 37967 18207
rect 37967 18173 37976 18207
rect 37924 18164 37976 18173
rect 39028 18275 39080 18284
rect 39028 18241 39062 18275
rect 39062 18241 39080 18275
rect 39028 18232 39080 18241
rect 45928 18368 45980 18420
rect 46756 18368 46808 18420
rect 48136 18368 48188 18420
rect 57704 18368 57756 18420
rect 58256 18411 58308 18420
rect 58256 18377 58265 18411
rect 58265 18377 58299 18411
rect 58299 18377 58308 18411
rect 58256 18368 58308 18377
rect 45744 18343 45796 18352
rect 40316 18232 40368 18284
rect 31760 18096 31812 18148
rect 37556 18096 37608 18148
rect 38660 18164 38712 18216
rect 40132 18164 40184 18216
rect 40868 18164 40920 18216
rect 41236 18207 41288 18216
rect 41236 18173 41245 18207
rect 41245 18173 41279 18207
rect 41279 18173 41288 18207
rect 41236 18164 41288 18173
rect 45744 18309 45778 18343
rect 45778 18309 45796 18343
rect 45744 18300 45796 18309
rect 47492 18300 47544 18352
rect 48228 18300 48280 18352
rect 49240 18300 49292 18352
rect 41696 18275 41748 18284
rect 41696 18241 41705 18275
rect 41705 18241 41739 18275
rect 41739 18241 41748 18275
rect 41696 18232 41748 18241
rect 42800 18232 42852 18284
rect 42892 18207 42944 18216
rect 42892 18173 42901 18207
rect 42901 18173 42935 18207
rect 42935 18173 42944 18207
rect 42892 18164 42944 18173
rect 44180 18164 44232 18216
rect 46848 18232 46900 18284
rect 48136 18207 48188 18216
rect 48136 18173 48145 18207
rect 48145 18173 48179 18207
rect 48179 18173 48188 18207
rect 48136 18164 48188 18173
rect 49424 18232 49476 18284
rect 58072 18275 58124 18284
rect 58072 18241 58081 18275
rect 58081 18241 58115 18275
rect 58115 18241 58124 18275
rect 58072 18232 58124 18241
rect 27804 18028 27856 18080
rect 27896 18028 27948 18080
rect 28356 18028 28408 18080
rect 29000 18028 29052 18080
rect 30840 18028 30892 18080
rect 31024 18071 31076 18080
rect 31024 18037 31033 18071
rect 31033 18037 31067 18071
rect 31067 18037 31076 18071
rect 31024 18028 31076 18037
rect 31392 18028 31444 18080
rect 33140 18028 33192 18080
rect 33508 18071 33560 18080
rect 33508 18037 33517 18071
rect 33517 18037 33551 18071
rect 33551 18037 33560 18071
rect 33508 18028 33560 18037
rect 33876 18028 33928 18080
rect 46204 18028 46256 18080
rect 47032 18028 47084 18080
rect 49700 18028 49752 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 11060 17620 11112 17672
rect 14188 17620 14240 17672
rect 16672 17824 16724 17876
rect 20076 17824 20128 17876
rect 26792 17867 26844 17876
rect 16028 17799 16080 17808
rect 16028 17765 16037 17799
rect 16037 17765 16071 17799
rect 16071 17765 16080 17799
rect 16028 17756 16080 17765
rect 15200 17663 15252 17672
rect 1860 17595 1912 17604
rect 1860 17561 1869 17595
rect 1869 17561 1903 17595
rect 1903 17561 1912 17595
rect 1860 17552 1912 17561
rect 11612 17484 11664 17536
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 17224 17620 17276 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 20720 17620 20772 17672
rect 14832 17552 14884 17604
rect 20904 17756 20956 17808
rect 24400 17756 24452 17808
rect 24584 17799 24636 17808
rect 24584 17765 24593 17799
rect 24593 17765 24627 17799
rect 24627 17765 24636 17799
rect 24584 17756 24636 17765
rect 21456 17688 21508 17740
rect 24492 17688 24544 17740
rect 26792 17833 26801 17867
rect 26801 17833 26835 17867
rect 26835 17833 26844 17867
rect 26792 17824 26844 17833
rect 26884 17824 26936 17876
rect 27896 17824 27948 17876
rect 29184 17824 29236 17876
rect 32496 17824 32548 17876
rect 41144 17824 41196 17876
rect 42800 17824 42852 17876
rect 27896 17688 27948 17740
rect 24584 17620 24636 17672
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 24860 17663 24912 17672
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 24032 17595 24084 17604
rect 15752 17484 15804 17536
rect 16580 17484 16632 17536
rect 16764 17484 16816 17536
rect 23756 17484 23808 17536
rect 24032 17561 24041 17595
rect 24041 17561 24075 17595
rect 24075 17561 24084 17595
rect 24032 17552 24084 17561
rect 26240 17620 26292 17672
rect 26424 17620 26476 17672
rect 41052 17756 41104 17808
rect 44364 17824 44416 17876
rect 45560 17824 45612 17876
rect 51724 17867 51776 17876
rect 28448 17620 28500 17672
rect 28908 17620 28960 17672
rect 31760 17731 31812 17740
rect 31760 17697 31769 17731
rect 31769 17697 31803 17731
rect 31803 17697 31812 17731
rect 31760 17688 31812 17697
rect 30288 17663 30340 17672
rect 30288 17629 30297 17663
rect 30297 17629 30331 17663
rect 30331 17629 30340 17663
rect 30288 17620 30340 17629
rect 31300 17620 31352 17672
rect 33324 17620 33376 17672
rect 29000 17552 29052 17604
rect 34888 17663 34940 17672
rect 34888 17629 34897 17663
rect 34897 17629 34931 17663
rect 34931 17629 34940 17663
rect 34888 17620 34940 17629
rect 35992 17620 36044 17672
rect 37464 17620 37516 17672
rect 38660 17620 38712 17672
rect 40592 17620 40644 17672
rect 42892 17663 42944 17672
rect 26884 17484 26936 17536
rect 27620 17484 27672 17536
rect 28172 17484 28224 17536
rect 28816 17484 28868 17536
rect 29368 17484 29420 17536
rect 33416 17527 33468 17536
rect 33416 17493 33425 17527
rect 33425 17493 33459 17527
rect 33459 17493 33468 17527
rect 33416 17484 33468 17493
rect 33692 17484 33744 17536
rect 34428 17552 34480 17604
rect 36820 17552 36872 17604
rect 37372 17552 37424 17604
rect 38568 17552 38620 17604
rect 41788 17552 41840 17604
rect 42616 17552 42668 17604
rect 42892 17629 42901 17663
rect 42901 17629 42935 17663
rect 42935 17629 42944 17663
rect 42892 17620 42944 17629
rect 44088 17620 44140 17672
rect 42984 17552 43036 17604
rect 43168 17595 43220 17604
rect 43168 17561 43202 17595
rect 43202 17561 43220 17595
rect 43168 17552 43220 17561
rect 44456 17552 44508 17604
rect 45560 17663 45612 17672
rect 45560 17629 45569 17663
rect 45569 17629 45603 17663
rect 45603 17629 45612 17663
rect 45560 17620 45612 17629
rect 46756 17552 46808 17604
rect 51724 17833 51733 17867
rect 51733 17833 51767 17867
rect 51767 17833 51776 17867
rect 51724 17824 51776 17833
rect 48136 17731 48188 17740
rect 48136 17697 48145 17731
rect 48145 17697 48179 17731
rect 48179 17697 48188 17731
rect 48136 17688 48188 17697
rect 47492 17663 47544 17672
rect 47492 17629 47501 17663
rect 47501 17629 47535 17663
rect 47535 17629 47544 17663
rect 47492 17620 47544 17629
rect 48044 17552 48096 17604
rect 48504 17552 48556 17604
rect 48596 17552 48648 17604
rect 37280 17527 37332 17536
rect 37280 17493 37289 17527
rect 37289 17493 37323 17527
rect 37323 17493 37332 17527
rect 37280 17484 37332 17493
rect 37648 17484 37700 17536
rect 39028 17484 39080 17536
rect 39212 17527 39264 17536
rect 39212 17493 39221 17527
rect 39221 17493 39255 17527
rect 39255 17493 39264 17527
rect 39212 17484 39264 17493
rect 40592 17484 40644 17536
rect 41696 17484 41748 17536
rect 46296 17484 46348 17536
rect 49240 17484 49292 17536
rect 49976 17552 50028 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 15200 17280 15252 17332
rect 21180 17280 21232 17332
rect 24124 17323 24176 17332
rect 24124 17289 24133 17323
rect 24133 17289 24167 17323
rect 24167 17289 24176 17323
rect 24124 17280 24176 17289
rect 25780 17280 25832 17332
rect 3700 17212 3752 17264
rect 13728 17212 13780 17264
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 13820 17144 13872 17196
rect 18604 17144 18656 17196
rect 19616 17212 19668 17264
rect 20536 17144 20588 17196
rect 16856 17076 16908 17128
rect 17224 17076 17276 17128
rect 18420 17076 18472 17128
rect 18880 17076 18932 17128
rect 18604 17008 18656 17060
rect 19616 17076 19668 17128
rect 20168 17076 20220 17128
rect 20720 17076 20772 17128
rect 21364 17076 21416 17128
rect 21916 17076 21968 17128
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 24492 17212 24544 17264
rect 25688 17212 25740 17264
rect 22192 17144 22244 17153
rect 27436 17280 27488 17332
rect 29828 17280 29880 17332
rect 30288 17280 30340 17332
rect 34796 17280 34848 17332
rect 26332 17187 26384 17196
rect 26332 17153 26341 17187
rect 26341 17153 26375 17187
rect 26375 17153 26384 17187
rect 26332 17144 26384 17153
rect 27068 17144 27120 17196
rect 27344 17187 27396 17196
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 14924 16940 14976 16992
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 16672 16940 16724 16992
rect 20904 17008 20956 17060
rect 26700 17076 26752 17128
rect 27620 17076 27672 17128
rect 33508 17212 33560 17264
rect 33692 17212 33744 17264
rect 31300 17144 31352 17196
rect 31208 17076 31260 17128
rect 32680 17144 32732 17196
rect 31576 17119 31628 17128
rect 31576 17085 31585 17119
rect 31585 17085 31619 17119
rect 31619 17085 31628 17119
rect 31576 17076 31628 17085
rect 23112 17008 23164 17060
rect 23756 17008 23808 17060
rect 36084 17144 36136 17196
rect 37188 17144 37240 17196
rect 37648 17187 37700 17196
rect 37648 17153 37657 17187
rect 37657 17153 37691 17187
rect 37691 17153 37700 17187
rect 37648 17144 37700 17153
rect 38660 17280 38712 17332
rect 39856 17280 39908 17332
rect 40592 17280 40644 17332
rect 41144 17280 41196 17332
rect 42156 17280 42208 17332
rect 43628 17280 43680 17332
rect 45652 17280 45704 17332
rect 49884 17323 49936 17332
rect 49884 17289 49893 17323
rect 49893 17289 49927 17323
rect 49927 17289 49936 17323
rect 49884 17280 49936 17289
rect 44364 17212 44416 17264
rect 49700 17212 49752 17264
rect 40224 17144 40276 17196
rect 33968 17076 34020 17128
rect 36360 17076 36412 17128
rect 36544 17119 36596 17128
rect 36544 17085 36553 17119
rect 36553 17085 36587 17119
rect 36587 17085 36596 17119
rect 36544 17076 36596 17085
rect 39948 17076 40000 17128
rect 19800 16940 19852 16992
rect 20812 16940 20864 16992
rect 24124 16940 24176 16992
rect 24768 16940 24820 16992
rect 25688 16940 25740 16992
rect 30288 16940 30340 16992
rect 30748 16940 30800 16992
rect 32404 16940 32456 16992
rect 36912 16983 36964 16992
rect 36912 16949 36921 16983
rect 36921 16949 36955 16983
rect 36955 16949 36964 16983
rect 36912 16940 36964 16949
rect 37832 16940 37884 16992
rect 38292 16940 38344 16992
rect 41052 17008 41104 17060
rect 40316 16983 40368 16992
rect 40316 16949 40325 16983
rect 40325 16949 40359 16983
rect 40359 16949 40368 16983
rect 40316 16940 40368 16949
rect 40408 16940 40460 16992
rect 41420 17076 41472 17128
rect 41512 16940 41564 16992
rect 43812 17144 43864 17196
rect 43996 17144 44048 17196
rect 45560 17144 45612 17196
rect 42984 17076 43036 17128
rect 44180 17119 44232 17128
rect 44180 17085 44189 17119
rect 44189 17085 44223 17119
rect 44223 17085 44232 17119
rect 44180 17076 44232 17085
rect 48136 17076 48188 17128
rect 43260 16983 43312 16992
rect 43260 16949 43269 16983
rect 43269 16949 43303 16983
rect 43303 16949 43312 16983
rect 43260 16940 43312 16949
rect 43996 16940 44048 16992
rect 45468 16940 45520 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 30380 16736 30432 16788
rect 30840 16736 30892 16788
rect 36084 16736 36136 16788
rect 16764 16668 16816 16720
rect 14832 16643 14884 16652
rect 14832 16609 14841 16643
rect 14841 16609 14875 16643
rect 14875 16609 14884 16643
rect 14832 16600 14884 16609
rect 16212 16600 16264 16652
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 13176 16532 13228 16584
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 15936 16575 15988 16584
rect 1860 16507 1912 16516
rect 1860 16473 1869 16507
rect 1869 16473 1903 16507
rect 1903 16473 1912 16507
rect 1860 16464 1912 16473
rect 12348 16464 12400 16516
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 19800 16600 19852 16652
rect 18052 16532 18104 16584
rect 18788 16532 18840 16584
rect 19432 16532 19484 16584
rect 20628 16532 20680 16584
rect 18604 16464 18656 16516
rect 23112 16532 23164 16584
rect 23388 16600 23440 16652
rect 11060 16396 11112 16448
rect 18328 16396 18380 16448
rect 22928 16396 22980 16448
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 24032 16532 24084 16584
rect 26056 16668 26108 16720
rect 26700 16668 26752 16720
rect 29368 16668 29420 16720
rect 32680 16668 32732 16720
rect 34980 16668 35032 16720
rect 27620 16600 27672 16652
rect 28724 16600 28776 16652
rect 29736 16643 29788 16652
rect 29736 16609 29745 16643
rect 29745 16609 29779 16643
rect 29779 16609 29788 16643
rect 29736 16600 29788 16609
rect 30748 16600 30800 16652
rect 35716 16600 35768 16652
rect 26884 16575 26936 16584
rect 25044 16464 25096 16516
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 29828 16532 29880 16584
rect 31024 16532 31076 16584
rect 35164 16532 35216 16584
rect 35348 16575 35400 16584
rect 35348 16541 35357 16575
rect 35357 16541 35391 16575
rect 35391 16541 35400 16575
rect 35348 16532 35400 16541
rect 36176 16643 36228 16652
rect 36176 16609 36185 16643
rect 36185 16609 36219 16643
rect 36219 16609 36228 16643
rect 36176 16600 36228 16609
rect 38292 16668 38344 16720
rect 38200 16600 38252 16652
rect 38476 16600 38528 16652
rect 38752 16668 38804 16720
rect 40224 16668 40276 16720
rect 40316 16668 40368 16720
rect 41788 16711 41840 16720
rect 39120 16600 39172 16652
rect 37280 16532 37332 16584
rect 40408 16532 40460 16584
rect 41052 16600 41104 16652
rect 41420 16643 41472 16652
rect 41420 16609 41429 16643
rect 41429 16609 41463 16643
rect 41463 16609 41472 16643
rect 41420 16600 41472 16609
rect 41788 16677 41797 16711
rect 41797 16677 41831 16711
rect 41831 16677 41840 16711
rect 41788 16668 41840 16677
rect 45560 16711 45612 16720
rect 42616 16532 42668 16584
rect 43260 16600 43312 16652
rect 43628 16600 43680 16652
rect 32220 16464 32272 16516
rect 28264 16396 28316 16448
rect 29644 16396 29696 16448
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 33048 16439 33100 16448
rect 33048 16405 33057 16439
rect 33057 16405 33091 16439
rect 33091 16405 33100 16439
rect 33048 16396 33100 16405
rect 34704 16396 34756 16448
rect 34980 16396 35032 16448
rect 35624 16396 35676 16448
rect 39764 16464 39816 16516
rect 40132 16396 40184 16448
rect 41512 16464 41564 16516
rect 40592 16439 40644 16448
rect 40592 16405 40601 16439
rect 40601 16405 40635 16439
rect 40635 16405 40644 16439
rect 40592 16396 40644 16405
rect 41144 16396 41196 16448
rect 41328 16396 41380 16448
rect 43168 16464 43220 16516
rect 44364 16600 44416 16652
rect 45560 16677 45569 16711
rect 45569 16677 45603 16711
rect 45603 16677 45612 16711
rect 45560 16668 45612 16677
rect 46848 16600 46900 16652
rect 44088 16396 44140 16448
rect 48136 16600 48188 16652
rect 48688 16464 48740 16516
rect 58164 16575 58216 16584
rect 58164 16541 58173 16575
rect 58173 16541 58207 16575
rect 58207 16541 58216 16575
rect 58164 16532 58216 16541
rect 57060 16507 57112 16516
rect 46756 16396 46808 16448
rect 57060 16473 57069 16507
rect 57069 16473 57103 16507
rect 57103 16473 57112 16507
rect 57060 16464 57112 16473
rect 49700 16439 49752 16448
rect 49700 16405 49709 16439
rect 49709 16405 49743 16439
rect 49743 16405 49752 16439
rect 49700 16396 49752 16405
rect 50804 16396 50856 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 1584 16192 1636 16244
rect 13176 16192 13228 16244
rect 24492 16192 24544 16244
rect 25044 16235 25096 16244
rect 25044 16201 25053 16235
rect 25053 16201 25087 16235
rect 25087 16201 25096 16235
rect 25044 16192 25096 16201
rect 26884 16192 26936 16244
rect 27988 16192 28040 16244
rect 29276 16192 29328 16244
rect 33048 16192 33100 16244
rect 33692 16235 33744 16244
rect 33692 16201 33701 16235
rect 33701 16201 33735 16235
rect 33735 16201 33744 16235
rect 33692 16192 33744 16201
rect 35624 16235 35676 16244
rect 35624 16201 35633 16235
rect 35633 16201 35667 16235
rect 35667 16201 35676 16235
rect 35624 16192 35676 16201
rect 36176 16192 36228 16244
rect 36452 16235 36504 16244
rect 36452 16201 36461 16235
rect 36461 16201 36495 16235
rect 36495 16201 36504 16235
rect 36452 16192 36504 16201
rect 38108 16192 38160 16244
rect 40040 16192 40092 16244
rect 40316 16192 40368 16244
rect 41052 16192 41104 16244
rect 41696 16235 41748 16244
rect 41696 16201 41705 16235
rect 41705 16201 41739 16235
rect 41739 16201 41748 16235
rect 41696 16192 41748 16201
rect 42984 16192 43036 16244
rect 11152 16124 11204 16176
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 13176 16099 13228 16108
rect 13176 16065 13185 16099
rect 13185 16065 13219 16099
rect 13219 16065 13228 16099
rect 13176 16056 13228 16065
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 15108 16056 15160 16108
rect 17776 16056 17828 16108
rect 18236 16056 18288 16108
rect 22100 16124 22152 16176
rect 22284 16167 22336 16176
rect 22284 16133 22318 16167
rect 22318 16133 22336 16167
rect 22284 16124 22336 16133
rect 22928 16124 22980 16176
rect 27528 16124 27580 16176
rect 27712 16124 27764 16176
rect 29828 16124 29880 16176
rect 32220 16124 32272 16176
rect 4068 15988 4120 16040
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 12164 15920 12216 15972
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13544 15988 13596 16040
rect 16856 15988 16908 16040
rect 21180 15988 21232 16040
rect 27160 16056 27212 16108
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 29644 16056 29696 16108
rect 32312 16099 32364 16108
rect 29828 15988 29880 16040
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32404 16056 32456 16108
rect 34428 16124 34480 16176
rect 34520 16099 34572 16108
rect 34520 16065 34554 16099
rect 34554 16065 34572 16099
rect 34520 16056 34572 16065
rect 35164 16124 35216 16176
rect 40592 16124 40644 16176
rect 41512 16124 41564 16176
rect 44548 16192 44600 16244
rect 48688 16235 48740 16244
rect 37464 16099 37516 16108
rect 13268 15920 13320 15972
rect 14556 15852 14608 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 17868 15852 17920 15904
rect 18236 15852 18288 15904
rect 24216 15920 24268 15972
rect 27620 15920 27672 15972
rect 24032 15852 24084 15904
rect 24492 15852 24544 15904
rect 30104 15852 30156 15904
rect 30656 15895 30708 15904
rect 30656 15861 30665 15895
rect 30665 15861 30699 15895
rect 30699 15861 30708 15895
rect 30656 15852 30708 15861
rect 33692 15988 33744 16040
rect 34244 16031 34296 16040
rect 34244 15997 34253 16031
rect 34253 15997 34287 16031
rect 34287 15997 34296 16031
rect 34244 15988 34296 15997
rect 35624 15988 35676 16040
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 37556 16056 37608 16108
rect 38200 16056 38252 16108
rect 39764 16099 39816 16108
rect 39764 16065 39773 16099
rect 39773 16065 39807 16099
rect 39807 16065 39816 16099
rect 40224 16099 40276 16108
rect 39764 16056 39816 16065
rect 40224 16065 40233 16099
rect 40233 16065 40267 16099
rect 40267 16065 40276 16099
rect 40224 16056 40276 16065
rect 40408 16099 40460 16108
rect 40408 16065 40417 16099
rect 40417 16065 40451 16099
rect 40451 16065 40460 16099
rect 40408 16056 40460 16065
rect 38660 15988 38712 16040
rect 39120 15988 39172 16040
rect 41788 16031 41840 16040
rect 33416 15852 33468 15904
rect 33968 15852 34020 15904
rect 36176 15920 36228 15972
rect 37188 15920 37240 15972
rect 39212 15920 39264 15972
rect 41788 15997 41797 16031
rect 41797 15997 41831 16031
rect 41831 15997 41840 16031
rect 41788 15988 41840 15997
rect 42156 16056 42208 16108
rect 43996 16056 44048 16108
rect 44272 16124 44324 16176
rect 45468 16124 45520 16176
rect 48688 16201 48697 16235
rect 48697 16201 48731 16235
rect 48731 16201 48740 16235
rect 48688 16192 48740 16201
rect 49976 16192 50028 16244
rect 40040 15920 40092 15972
rect 43168 15920 43220 15972
rect 37740 15852 37792 15904
rect 40592 15895 40644 15904
rect 40592 15861 40601 15895
rect 40601 15861 40635 15895
rect 40635 15861 40644 15895
rect 40592 15852 40644 15861
rect 41328 15895 41380 15904
rect 41328 15861 41337 15895
rect 41337 15861 41371 15895
rect 41371 15861 41380 15895
rect 41328 15852 41380 15861
rect 43444 15895 43496 15904
rect 43444 15861 43453 15895
rect 43453 15861 43487 15895
rect 43487 15861 43496 15895
rect 43444 15852 43496 15861
rect 45744 16056 45796 16108
rect 46480 16056 46532 16108
rect 49700 16124 49752 16176
rect 46204 16031 46256 16040
rect 46204 15997 46213 16031
rect 46213 15997 46247 16031
rect 46247 15997 46256 16031
rect 46204 15988 46256 15997
rect 46848 15988 46900 16040
rect 48872 16056 48924 16108
rect 49240 16056 49292 16108
rect 49424 15988 49476 16040
rect 57796 15920 57848 15972
rect 44180 15852 44232 15904
rect 46572 15895 46624 15904
rect 46572 15861 46581 15895
rect 46581 15861 46615 15895
rect 46615 15861 46624 15895
rect 46572 15852 46624 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 17868 15648 17920 15700
rect 17316 15580 17368 15632
rect 18236 15580 18288 15632
rect 20536 15580 20588 15632
rect 23480 15580 23532 15632
rect 24768 15580 24820 15632
rect 25228 15580 25280 15632
rect 26516 15580 26568 15632
rect 27160 15648 27212 15700
rect 41788 15648 41840 15700
rect 42892 15691 42944 15700
rect 42892 15657 42901 15691
rect 42901 15657 42935 15691
rect 42935 15657 42944 15691
rect 42892 15648 42944 15657
rect 45744 15691 45796 15700
rect 45744 15657 45753 15691
rect 45753 15657 45787 15691
rect 45787 15657 45796 15691
rect 45744 15648 45796 15657
rect 48136 15691 48188 15700
rect 48136 15657 48145 15691
rect 48145 15657 48179 15691
rect 48179 15657 48188 15691
rect 48136 15648 48188 15657
rect 2412 15512 2464 15564
rect 16396 15512 16448 15564
rect 17776 15512 17828 15564
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 13912 15444 13964 15496
rect 14556 15444 14608 15496
rect 16580 15487 16632 15496
rect 16304 15376 16356 15428
rect 16580 15453 16589 15487
rect 16589 15453 16623 15487
rect 16623 15453 16632 15487
rect 16580 15444 16632 15453
rect 19432 15444 19484 15496
rect 25136 15512 25188 15564
rect 26056 15512 26108 15564
rect 28080 15555 28132 15564
rect 28080 15521 28089 15555
rect 28089 15521 28123 15555
rect 28123 15521 28132 15555
rect 28080 15512 28132 15521
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 25044 15444 25096 15496
rect 29000 15444 29052 15496
rect 27160 15376 27212 15428
rect 19984 15308 20036 15360
rect 20904 15351 20956 15360
rect 20904 15317 20913 15351
rect 20913 15317 20947 15351
rect 20947 15317 20956 15351
rect 20904 15308 20956 15317
rect 25044 15308 25096 15360
rect 25228 15308 25280 15360
rect 25504 15351 25556 15360
rect 25504 15317 25513 15351
rect 25513 15317 25547 15351
rect 25547 15317 25556 15351
rect 25504 15308 25556 15317
rect 25872 15308 25924 15360
rect 28448 15376 28500 15428
rect 31300 15580 31352 15632
rect 31484 15580 31536 15632
rect 33416 15580 33468 15632
rect 34060 15580 34112 15632
rect 29920 15512 29972 15564
rect 30932 15444 30984 15496
rect 32312 15444 32364 15496
rect 31576 15376 31628 15428
rect 31852 15376 31904 15428
rect 27528 15308 27580 15360
rect 29460 15308 29512 15360
rect 30564 15308 30616 15360
rect 30748 15351 30800 15360
rect 30748 15317 30757 15351
rect 30757 15317 30791 15351
rect 30791 15317 30800 15351
rect 30748 15308 30800 15317
rect 31484 15308 31536 15360
rect 34428 15512 34480 15564
rect 34060 15487 34112 15496
rect 34060 15453 34069 15487
rect 34069 15453 34103 15487
rect 34103 15453 34112 15487
rect 34060 15444 34112 15453
rect 34704 15444 34756 15496
rect 35072 15487 35124 15496
rect 35072 15453 35081 15487
rect 35081 15453 35115 15487
rect 35115 15453 35124 15487
rect 35072 15444 35124 15453
rect 37556 15580 37608 15632
rect 39948 15580 40000 15632
rect 35440 15512 35492 15564
rect 36912 15512 36964 15564
rect 38108 15555 38160 15564
rect 34888 15308 34940 15360
rect 35348 15308 35400 15360
rect 36084 15308 36136 15360
rect 36636 15308 36688 15360
rect 38108 15521 38117 15555
rect 38117 15521 38151 15555
rect 38151 15521 38160 15555
rect 38108 15512 38160 15521
rect 37740 15444 37792 15496
rect 41052 15512 41104 15564
rect 39212 15444 39264 15496
rect 39856 15444 39908 15496
rect 38844 15376 38896 15428
rect 41512 15444 41564 15496
rect 44088 15444 44140 15496
rect 44548 15444 44600 15496
rect 45192 15487 45244 15496
rect 45192 15453 45201 15487
rect 45201 15453 45235 15487
rect 45235 15453 45244 15487
rect 45192 15444 45244 15453
rect 46664 15444 46716 15496
rect 38752 15308 38804 15360
rect 40132 15376 40184 15428
rect 44364 15376 44416 15428
rect 46756 15376 46808 15428
rect 48872 15512 48924 15564
rect 47124 15444 47176 15496
rect 49424 15487 49476 15496
rect 49424 15453 49433 15487
rect 49433 15453 49467 15487
rect 49467 15453 49476 15487
rect 49424 15444 49476 15453
rect 47216 15376 47268 15428
rect 48044 15376 48096 15428
rect 49792 15444 49844 15496
rect 56508 15444 56560 15496
rect 58164 15419 58216 15428
rect 40316 15308 40368 15360
rect 40592 15308 40644 15360
rect 43260 15308 43312 15360
rect 46204 15308 46256 15360
rect 58164 15385 58173 15419
rect 58173 15385 58207 15419
rect 58207 15385 58216 15419
rect 58164 15376 58216 15385
rect 50712 15351 50764 15360
rect 50712 15317 50721 15351
rect 50721 15317 50755 15351
rect 50755 15317 50764 15351
rect 50712 15308 50764 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 11244 14968 11296 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 2412 14943 2464 14952
rect 2412 14909 2421 14943
rect 2421 14909 2455 14943
rect 2455 14909 2464 14943
rect 2412 14900 2464 14909
rect 8208 14900 8260 14952
rect 13912 14968 13964 15020
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 16028 15104 16080 15156
rect 17040 15104 17092 15156
rect 25136 15147 25188 15156
rect 18328 15036 18380 15088
rect 20904 15036 20956 15088
rect 14004 14968 14056 14977
rect 17960 14968 18012 15020
rect 10416 14832 10468 14884
rect 16856 14900 16908 14952
rect 17224 14900 17276 14952
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 15384 14832 15436 14884
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22468 15036 22520 15088
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 28356 15104 28408 15156
rect 30840 15147 30892 15156
rect 30840 15113 30849 15147
rect 30849 15113 30883 15147
rect 30883 15113 30892 15147
rect 30840 15104 30892 15113
rect 30932 15104 30984 15156
rect 36176 15104 36228 15156
rect 36636 15104 36688 15156
rect 38844 15104 38896 15156
rect 39120 15104 39172 15156
rect 41788 15104 41840 15156
rect 44272 15104 44324 15156
rect 44456 15104 44508 15156
rect 29000 15036 29052 15088
rect 31024 15036 31076 15088
rect 32772 15079 32824 15088
rect 32772 15045 32781 15079
rect 32781 15045 32815 15079
rect 32815 15045 32824 15079
rect 33968 15079 34020 15088
rect 32772 15036 32824 15045
rect 33968 15045 34002 15079
rect 34002 15045 34020 15079
rect 33968 15036 34020 15045
rect 34336 15036 34388 15088
rect 22100 14968 22152 14977
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 30656 14968 30708 15020
rect 25596 14900 25648 14952
rect 30564 14900 30616 14952
rect 31116 14900 31168 14952
rect 32036 14968 32088 15020
rect 36084 15036 36136 15088
rect 37464 15036 37516 15088
rect 38016 15036 38068 15088
rect 39396 15036 39448 15088
rect 39580 15036 39632 15088
rect 39856 15036 39908 15088
rect 41328 15036 41380 15088
rect 13452 14764 13504 14816
rect 15568 14764 15620 14816
rect 20904 14764 20956 14816
rect 22284 14764 22336 14816
rect 22836 14764 22888 14816
rect 23388 14764 23440 14816
rect 25504 14832 25556 14884
rect 23572 14764 23624 14816
rect 31208 14832 31260 14884
rect 27344 14764 27396 14816
rect 27804 14764 27856 14816
rect 28080 14764 28132 14816
rect 28908 14764 28960 14816
rect 31484 14832 31536 14884
rect 32956 14900 33008 14952
rect 33692 14943 33744 14952
rect 33692 14909 33701 14943
rect 33701 14909 33735 14943
rect 33735 14909 33744 14943
rect 33692 14900 33744 14909
rect 35532 14900 35584 14952
rect 31576 14764 31628 14816
rect 35624 14832 35676 14884
rect 36176 14900 36228 14952
rect 36820 14968 36872 15020
rect 36452 14900 36504 14952
rect 36636 14900 36688 14952
rect 37188 14900 37240 14952
rect 37648 15011 37700 15020
rect 37648 14977 37657 15011
rect 37657 14977 37691 15011
rect 37691 14977 37700 15011
rect 37648 14968 37700 14977
rect 39120 14968 39172 15020
rect 38108 14900 38160 14952
rect 38752 14832 38804 14884
rect 39304 14943 39356 14952
rect 39304 14909 39313 14943
rect 39313 14909 39347 14943
rect 39347 14909 39356 14943
rect 39304 14900 39356 14909
rect 38844 14807 38896 14816
rect 38844 14773 38853 14807
rect 38853 14773 38887 14807
rect 38887 14773 38896 14807
rect 38844 14764 38896 14773
rect 39212 14764 39264 14816
rect 40316 14764 40368 14816
rect 40592 14764 40644 14816
rect 40776 14764 40828 14816
rect 42340 14968 42392 15020
rect 42616 14900 42668 14952
rect 43444 14968 43496 15020
rect 43628 15011 43680 15020
rect 43628 14977 43637 15011
rect 43637 14977 43671 15011
rect 43671 14977 43680 15011
rect 43628 14968 43680 14977
rect 44088 14968 44140 15020
rect 44180 14968 44232 15020
rect 44732 15011 44784 15020
rect 44732 14977 44766 15011
rect 44766 14977 44784 15011
rect 44732 14968 44784 14977
rect 45468 14968 45520 15020
rect 46664 15036 46716 15088
rect 47492 15036 47544 15088
rect 48228 15036 48280 15088
rect 50712 15036 50764 15088
rect 43720 14832 43772 14884
rect 55864 14968 55916 15020
rect 47124 14764 47176 14816
rect 57612 14900 57664 14952
rect 49792 14875 49844 14884
rect 49792 14841 49801 14875
rect 49801 14841 49835 14875
rect 49835 14841 49844 14875
rect 49792 14832 49844 14841
rect 50988 14832 51040 14884
rect 49700 14764 49752 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 11428 14560 11480 14612
rect 13452 14560 13504 14612
rect 24584 14603 24636 14612
rect 13912 14424 13964 14476
rect 15200 14424 15252 14476
rect 15936 14424 15988 14476
rect 8944 14356 8996 14408
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 11612 14356 11664 14408
rect 13728 14356 13780 14408
rect 16856 14424 16908 14476
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 20904 14492 20956 14544
rect 22100 14492 22152 14544
rect 24308 14492 24360 14544
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 25596 14560 25648 14612
rect 22652 14424 22704 14476
rect 26608 14492 26660 14544
rect 30748 14560 30800 14612
rect 34704 14560 34756 14612
rect 36176 14560 36228 14612
rect 37096 14560 37148 14612
rect 37556 14560 37608 14612
rect 42340 14560 42392 14612
rect 42708 14603 42760 14612
rect 42708 14569 42717 14603
rect 42717 14569 42751 14603
rect 42751 14569 42760 14603
rect 42708 14560 42760 14569
rect 46756 14603 46808 14612
rect 46756 14569 46765 14603
rect 46765 14569 46799 14603
rect 46799 14569 46808 14603
rect 46756 14560 46808 14569
rect 30932 14492 30984 14544
rect 31116 14535 31168 14544
rect 31116 14501 31125 14535
rect 31125 14501 31159 14535
rect 31159 14501 31168 14535
rect 31116 14492 31168 14501
rect 33876 14492 33928 14544
rect 34244 14492 34296 14544
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 22836 14356 22888 14408
rect 23112 14356 23164 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 28356 14424 28408 14476
rect 28540 14467 28592 14476
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 28540 14424 28592 14433
rect 29368 14424 29420 14476
rect 34336 14424 34388 14476
rect 34704 14424 34756 14476
rect 25504 14356 25556 14408
rect 29828 14356 29880 14408
rect 33876 14356 33928 14408
rect 10968 14220 11020 14272
rect 13084 14220 13136 14272
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 16028 14220 16080 14272
rect 17132 14220 17184 14272
rect 25596 14288 25648 14340
rect 30012 14331 30064 14340
rect 30012 14297 30046 14331
rect 30046 14297 30064 14331
rect 30012 14288 30064 14297
rect 31300 14288 31352 14340
rect 33968 14288 34020 14340
rect 34796 14356 34848 14408
rect 35716 14424 35768 14476
rect 36636 14492 36688 14544
rect 37188 14492 37240 14544
rect 41328 14492 41380 14544
rect 41420 14492 41472 14544
rect 38016 14467 38068 14476
rect 38016 14433 38025 14467
rect 38025 14433 38059 14467
rect 38059 14433 38068 14467
rect 38016 14424 38068 14433
rect 39212 14424 39264 14476
rect 36360 14356 36412 14408
rect 36176 14288 36228 14340
rect 36636 14331 36688 14340
rect 35624 14220 35676 14272
rect 36084 14220 36136 14272
rect 36268 14220 36320 14272
rect 36636 14297 36645 14331
rect 36645 14297 36679 14331
rect 36679 14297 36688 14331
rect 36636 14288 36688 14297
rect 37740 14356 37792 14408
rect 38844 14356 38896 14408
rect 40224 14399 40276 14408
rect 40224 14365 40233 14399
rect 40233 14365 40267 14399
rect 40267 14365 40276 14399
rect 40224 14356 40276 14365
rect 40776 14424 40828 14476
rect 41512 14424 41564 14476
rect 41236 14399 41288 14408
rect 41236 14365 41245 14399
rect 41245 14365 41279 14399
rect 41279 14365 41288 14399
rect 41236 14356 41288 14365
rect 41328 14399 41380 14408
rect 41328 14365 41337 14399
rect 41337 14365 41371 14399
rect 41371 14365 41380 14399
rect 41328 14356 41380 14365
rect 37464 14288 37516 14340
rect 38752 14288 38804 14340
rect 40592 14288 40644 14340
rect 41052 14288 41104 14340
rect 41880 14356 41932 14408
rect 42708 14356 42760 14408
rect 43260 14399 43312 14408
rect 43260 14365 43269 14399
rect 43269 14365 43303 14399
rect 43303 14365 43312 14399
rect 43260 14356 43312 14365
rect 43352 14288 43404 14340
rect 43812 14356 43864 14408
rect 44088 14492 44140 14544
rect 44824 14492 44876 14544
rect 44180 14399 44232 14408
rect 44180 14365 44189 14399
rect 44189 14365 44223 14399
rect 44223 14365 44232 14399
rect 44180 14356 44232 14365
rect 44456 14424 44508 14476
rect 46756 14424 46808 14476
rect 56508 14560 56560 14612
rect 45468 14356 45520 14408
rect 57980 14399 58032 14408
rect 57980 14365 57989 14399
rect 57989 14365 58023 14399
rect 58023 14365 58032 14399
rect 57980 14356 58032 14365
rect 38660 14220 38712 14272
rect 39396 14263 39448 14272
rect 39396 14229 39405 14263
rect 39405 14229 39439 14263
rect 39439 14229 39448 14263
rect 39396 14220 39448 14229
rect 39672 14220 39724 14272
rect 43720 14220 43772 14272
rect 44456 14288 44508 14340
rect 44364 14220 44416 14272
rect 44824 14220 44876 14272
rect 46572 14288 46624 14340
rect 48136 14288 48188 14340
rect 46848 14220 46900 14272
rect 58072 14263 58124 14272
rect 58072 14229 58081 14263
rect 58081 14229 58115 14263
rect 58115 14229 58124 14263
rect 58072 14220 58124 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 11060 14016 11112 14068
rect 12440 14016 12492 14068
rect 10692 13991 10744 14000
rect 10692 13957 10701 13991
rect 10701 13957 10735 13991
rect 10735 13957 10744 13991
rect 10692 13948 10744 13957
rect 12164 13948 12216 14000
rect 12256 13923 12308 13932
rect 12256 13889 12265 13923
rect 12265 13889 12299 13923
rect 12299 13889 12308 13923
rect 12256 13880 12308 13889
rect 15936 14016 15988 14068
rect 17224 14016 17276 14068
rect 17408 14016 17460 14068
rect 13084 13948 13136 14000
rect 13544 13880 13596 13932
rect 15292 13880 15344 13932
rect 16212 13880 16264 13932
rect 16488 13880 16540 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 26792 13948 26844 14000
rect 19248 13880 19300 13932
rect 24308 13923 24360 13932
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 11428 13812 11480 13864
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 12072 13812 12124 13864
rect 12532 13812 12584 13864
rect 12624 13812 12676 13864
rect 14740 13812 14792 13864
rect 22192 13812 22244 13864
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 7840 13744 7892 13796
rect 13728 13744 13780 13796
rect 13912 13744 13964 13796
rect 16028 13744 16080 13796
rect 18052 13744 18104 13796
rect 10048 13676 10100 13728
rect 12900 13676 12952 13728
rect 14464 13676 14516 13728
rect 14648 13676 14700 13728
rect 18236 13676 18288 13728
rect 21824 13744 21876 13796
rect 22376 13744 22428 13796
rect 24308 13889 24317 13923
rect 24317 13889 24351 13923
rect 24351 13889 24360 13923
rect 24308 13880 24360 13889
rect 25228 13880 25280 13932
rect 30012 13948 30064 14000
rect 30196 13991 30248 14000
rect 30196 13957 30230 13991
rect 30230 13957 30248 13991
rect 30196 13948 30248 13957
rect 31024 13948 31076 14000
rect 29828 13880 29880 13932
rect 36268 14016 36320 14068
rect 37096 14016 37148 14068
rect 37372 14016 37424 14068
rect 38660 14016 38712 14068
rect 34336 13948 34388 14000
rect 29276 13812 29328 13864
rect 32956 13880 33008 13932
rect 34888 13880 34940 13932
rect 35247 13923 35299 13932
rect 35247 13889 35279 13923
rect 35279 13889 35299 13923
rect 35247 13880 35299 13889
rect 37280 13880 37332 13932
rect 37556 13923 37608 13932
rect 37556 13889 37565 13923
rect 37565 13889 37599 13923
rect 37599 13889 37608 13923
rect 37556 13880 37608 13889
rect 38016 13880 38068 13932
rect 39672 13948 39724 14000
rect 40408 14016 40460 14068
rect 40776 14016 40828 14068
rect 41880 14059 41932 14068
rect 41236 13948 41288 14000
rect 41052 13880 41104 13932
rect 41604 13991 41656 14000
rect 41604 13957 41613 13991
rect 41613 13957 41647 13991
rect 41647 13957 41656 13991
rect 41604 13948 41656 13957
rect 41880 14025 41889 14059
rect 41889 14025 41923 14059
rect 41923 14025 41932 14059
rect 41880 14016 41932 14025
rect 43628 14016 43680 14068
rect 44732 14059 44784 14068
rect 44732 14025 44741 14059
rect 44741 14025 44775 14059
rect 44775 14025 44784 14059
rect 44732 14016 44784 14025
rect 48136 14059 48188 14068
rect 30932 13812 30984 13864
rect 33876 13812 33928 13864
rect 34796 13812 34848 13864
rect 36084 13812 36136 13864
rect 37464 13812 37516 13864
rect 28172 13744 28224 13796
rect 40408 13812 40460 13864
rect 40776 13812 40828 13864
rect 22652 13676 22704 13728
rect 23112 13676 23164 13728
rect 25228 13676 25280 13728
rect 25504 13719 25556 13728
rect 25504 13685 25513 13719
rect 25513 13685 25547 13719
rect 25547 13685 25556 13719
rect 25504 13676 25556 13685
rect 31116 13676 31168 13728
rect 34244 13676 34296 13728
rect 34336 13676 34388 13728
rect 41052 13744 41104 13796
rect 41328 13744 41380 13796
rect 43720 13948 43772 14000
rect 43352 13923 43404 13932
rect 43352 13889 43361 13923
rect 43361 13889 43395 13923
rect 43395 13889 43404 13923
rect 43352 13880 43404 13889
rect 44088 13880 44140 13932
rect 43812 13812 43864 13864
rect 43996 13812 44048 13864
rect 46848 13991 46900 14000
rect 46848 13957 46857 13991
rect 46857 13957 46891 13991
rect 46891 13957 46900 13991
rect 46848 13948 46900 13957
rect 44824 13880 44876 13932
rect 46664 13923 46716 13932
rect 46664 13889 46673 13923
rect 46673 13889 46707 13923
rect 46707 13889 46716 13923
rect 46664 13880 46716 13889
rect 46756 13880 46808 13932
rect 47492 13880 47544 13932
rect 48136 14025 48145 14059
rect 48145 14025 48179 14059
rect 48179 14025 48188 14059
rect 48136 14016 48188 14025
rect 48228 14016 48280 14068
rect 57244 14016 57296 14068
rect 48872 13880 48924 13932
rect 50804 13812 50856 13864
rect 40408 13676 40460 13728
rect 41512 13676 41564 13728
rect 49240 13676 49292 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 12808 13404 12860 13456
rect 16028 13447 16080 13456
rect 11612 13336 11664 13388
rect 13544 13379 13596 13388
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 13912 13336 13964 13388
rect 14464 13336 14516 13388
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11888 13268 11940 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 12900 13268 12952 13320
rect 14096 13268 14148 13320
rect 14556 13268 14608 13320
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 16212 13472 16264 13524
rect 18972 13404 19024 13456
rect 21916 13472 21968 13524
rect 25504 13472 25556 13524
rect 28172 13472 28224 13524
rect 31944 13472 31996 13524
rect 33232 13472 33284 13524
rect 35440 13472 35492 13524
rect 35808 13472 35860 13524
rect 38384 13472 38436 13524
rect 41052 13472 41104 13524
rect 45192 13472 45244 13524
rect 32312 13404 32364 13456
rect 32864 13404 32916 13456
rect 34336 13404 34388 13456
rect 34796 13404 34848 13456
rect 36268 13404 36320 13456
rect 37096 13404 37148 13456
rect 37740 13404 37792 13456
rect 40316 13404 40368 13456
rect 40408 13404 40460 13456
rect 40684 13404 40736 13456
rect 41420 13404 41472 13456
rect 41512 13404 41564 13456
rect 43444 13404 43496 13456
rect 14924 13336 14976 13388
rect 19432 13379 19484 13388
rect 15016 13268 15068 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 16212 13268 16264 13320
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 11060 13132 11112 13184
rect 12348 13132 12400 13184
rect 12992 13132 13044 13184
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 13912 13132 13964 13184
rect 14096 13132 14148 13184
rect 14832 13132 14884 13184
rect 16028 13200 16080 13252
rect 16856 13268 16908 13320
rect 17500 13268 17552 13320
rect 17960 13268 18012 13320
rect 19432 13345 19441 13379
rect 19441 13345 19475 13379
rect 19475 13345 19484 13379
rect 19432 13336 19484 13345
rect 26056 13336 26108 13388
rect 27988 13336 28040 13388
rect 29920 13336 29972 13388
rect 21640 13268 21692 13320
rect 21916 13268 21968 13320
rect 22468 13268 22520 13320
rect 25136 13268 25188 13320
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 26700 13268 26752 13320
rect 17408 13200 17460 13252
rect 18052 13200 18104 13252
rect 18788 13200 18840 13252
rect 20260 13200 20312 13252
rect 20904 13200 20956 13252
rect 20812 13175 20864 13184
rect 20812 13141 20821 13175
rect 20821 13141 20855 13175
rect 20855 13141 20864 13175
rect 20812 13132 20864 13141
rect 21456 13132 21508 13184
rect 32680 13336 32732 13388
rect 33600 13311 33652 13320
rect 24308 13132 24360 13184
rect 26148 13132 26200 13184
rect 27528 13132 27580 13184
rect 28264 13132 28316 13184
rect 30104 13132 30156 13184
rect 30380 13200 30432 13252
rect 33600 13277 33609 13311
rect 33609 13277 33643 13311
rect 33643 13277 33652 13311
rect 33600 13268 33652 13277
rect 35164 13379 35216 13388
rect 35164 13345 35173 13379
rect 35173 13345 35207 13379
rect 35207 13345 35216 13379
rect 35164 13336 35216 13345
rect 40132 13336 40184 13388
rect 37280 13311 37332 13320
rect 32956 13243 33008 13252
rect 32956 13209 32965 13243
rect 32965 13209 32999 13243
rect 32999 13209 33008 13243
rect 32956 13200 33008 13209
rect 33416 13243 33468 13252
rect 33416 13209 33425 13243
rect 33425 13209 33459 13243
rect 33459 13209 33468 13243
rect 33416 13200 33468 13209
rect 34980 13200 35032 13252
rect 35532 13200 35584 13252
rect 37280 13277 37289 13311
rect 37289 13277 37323 13311
rect 37323 13277 37332 13311
rect 37280 13268 37332 13277
rect 37740 13268 37792 13320
rect 38384 13268 38436 13320
rect 40040 13311 40092 13320
rect 34244 13132 34296 13184
rect 38660 13200 38712 13252
rect 38844 13200 38896 13252
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 43628 13336 43680 13388
rect 57520 13336 57572 13388
rect 58164 13379 58216 13388
rect 58164 13345 58173 13379
rect 58173 13345 58207 13379
rect 58207 13345 58216 13379
rect 58164 13336 58216 13345
rect 39764 13200 39816 13252
rect 40776 13268 40828 13320
rect 41052 13311 41104 13320
rect 41052 13277 41061 13311
rect 41061 13277 41095 13311
rect 41095 13277 41104 13311
rect 41052 13268 41104 13277
rect 41144 13268 41196 13320
rect 41420 13268 41472 13320
rect 41972 13268 42024 13320
rect 35808 13132 35860 13184
rect 39948 13132 40000 13184
rect 41420 13132 41472 13184
rect 42156 13311 42208 13320
rect 42156 13277 42165 13311
rect 42165 13277 42199 13311
rect 42199 13277 42208 13311
rect 42156 13268 42208 13277
rect 51080 13268 51132 13320
rect 57060 13243 57112 13252
rect 57060 13209 57069 13243
rect 57069 13209 57103 13243
rect 57103 13209 57112 13243
rect 57060 13200 57112 13209
rect 48964 13132 49016 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 12624 12928 12676 12980
rect 13176 12928 13228 12980
rect 15660 12928 15712 12980
rect 15752 12928 15804 12980
rect 12716 12860 12768 12912
rect 13544 12860 13596 12912
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 11888 12792 11940 12844
rect 12440 12792 12492 12844
rect 13728 12792 13780 12844
rect 14740 12860 14792 12912
rect 17408 12860 17460 12912
rect 18236 12928 18288 12980
rect 26976 12928 27028 12980
rect 27344 12928 27396 12980
rect 16856 12792 16908 12844
rect 17316 12792 17368 12844
rect 17960 12835 18012 12844
rect 17960 12801 17987 12835
rect 17987 12801 18012 12835
rect 17960 12792 18012 12801
rect 18236 12792 18288 12844
rect 20260 12860 20312 12912
rect 22284 12903 22336 12912
rect 22284 12869 22318 12903
rect 22318 12869 22336 12903
rect 22284 12860 22336 12869
rect 25044 12860 25096 12912
rect 26056 12860 26108 12912
rect 26516 12860 26568 12912
rect 27620 12928 27672 12980
rect 10692 12767 10744 12776
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 10968 12699 11020 12708
rect 10968 12665 10977 12699
rect 10977 12665 11011 12699
rect 11011 12665 11020 12699
rect 10968 12656 11020 12665
rect 12348 12699 12400 12708
rect 12348 12665 12357 12699
rect 12357 12665 12391 12699
rect 12391 12665 12400 12699
rect 12348 12656 12400 12665
rect 13544 12724 13596 12776
rect 14188 12724 14240 12776
rect 14556 12724 14608 12776
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 13728 12656 13780 12708
rect 15844 12656 15896 12708
rect 13820 12588 13872 12640
rect 13912 12588 13964 12640
rect 14740 12588 14792 12640
rect 14832 12588 14884 12640
rect 18604 12724 18656 12776
rect 20260 12724 20312 12776
rect 20352 12724 20404 12776
rect 20812 12724 20864 12776
rect 18052 12588 18104 12640
rect 20720 12656 20772 12708
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 26424 12792 26476 12844
rect 24216 12724 24268 12776
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27804 12860 27856 12912
rect 32496 12903 32548 12912
rect 27344 12792 27396 12801
rect 28172 12835 28224 12844
rect 28172 12801 28181 12835
rect 28181 12801 28215 12835
rect 28215 12801 28224 12835
rect 28172 12792 28224 12801
rect 28264 12792 28316 12844
rect 32496 12869 32505 12903
rect 32505 12869 32539 12903
rect 32539 12869 32548 12903
rect 32496 12860 32548 12869
rect 32588 12903 32640 12912
rect 32588 12869 32597 12903
rect 32597 12869 32631 12903
rect 32631 12869 32640 12903
rect 36452 12903 36504 12912
rect 32588 12860 32640 12869
rect 36452 12869 36461 12903
rect 36461 12869 36495 12903
rect 36495 12869 36504 12903
rect 36452 12860 36504 12869
rect 37096 12860 37148 12912
rect 40960 12903 41012 12912
rect 40960 12869 40969 12903
rect 40969 12869 41003 12903
rect 41003 12869 41012 12903
rect 40960 12860 41012 12869
rect 46664 12928 46716 12980
rect 51908 12860 51960 12912
rect 31392 12767 31444 12776
rect 31392 12733 31401 12767
rect 31401 12733 31435 12767
rect 31435 12733 31444 12767
rect 31392 12724 31444 12733
rect 31484 12767 31536 12776
rect 31484 12733 31493 12767
rect 31493 12733 31527 12767
rect 31527 12733 31536 12767
rect 31484 12724 31536 12733
rect 23480 12656 23532 12708
rect 27344 12656 27396 12708
rect 29736 12656 29788 12708
rect 23388 12631 23440 12640
rect 23388 12597 23397 12631
rect 23397 12597 23431 12631
rect 23431 12597 23440 12631
rect 23388 12588 23440 12597
rect 27574 12588 27626 12640
rect 32956 12792 33008 12844
rect 34796 12792 34848 12844
rect 35808 12792 35860 12844
rect 36084 12835 36136 12844
rect 36084 12801 36093 12835
rect 36093 12801 36127 12835
rect 36127 12801 36136 12835
rect 36084 12792 36136 12801
rect 36544 12792 36596 12844
rect 36820 12792 36872 12844
rect 39672 12835 39724 12844
rect 39672 12801 39681 12835
rect 39681 12801 39715 12835
rect 39715 12801 39724 12835
rect 39672 12792 39724 12801
rect 39948 12792 40000 12844
rect 40684 12835 40736 12844
rect 40684 12801 40693 12835
rect 40693 12801 40727 12835
rect 40727 12801 40736 12835
rect 40684 12792 40736 12801
rect 40776 12792 40828 12844
rect 41328 12792 41380 12844
rect 41880 12835 41932 12844
rect 41880 12801 41889 12835
rect 41889 12801 41923 12835
rect 41923 12801 41932 12835
rect 41880 12792 41932 12801
rect 35164 12724 35216 12776
rect 37372 12724 37424 12776
rect 37740 12767 37792 12776
rect 37740 12733 37749 12767
rect 37749 12733 37783 12767
rect 37783 12733 37792 12767
rect 37740 12724 37792 12733
rect 38936 12767 38988 12776
rect 38936 12733 38945 12767
rect 38945 12733 38979 12767
rect 38979 12733 38988 12767
rect 38936 12724 38988 12733
rect 39764 12724 39816 12776
rect 32864 12699 32916 12708
rect 32864 12665 32873 12699
rect 32873 12665 32907 12699
rect 32907 12665 32916 12699
rect 32864 12656 32916 12665
rect 32680 12588 32732 12640
rect 37280 12656 37332 12708
rect 35440 12631 35492 12640
rect 35440 12597 35449 12631
rect 35449 12597 35483 12631
rect 35483 12597 35492 12631
rect 35440 12588 35492 12597
rect 35808 12588 35860 12640
rect 39120 12656 39172 12708
rect 39580 12656 39632 12708
rect 41420 12724 41472 12776
rect 42064 12724 42116 12776
rect 43076 12767 43128 12776
rect 43076 12733 43085 12767
rect 43085 12733 43119 12767
rect 43119 12733 43128 12767
rect 43076 12724 43128 12733
rect 43168 12767 43220 12776
rect 43168 12733 43177 12767
rect 43177 12733 43211 12767
rect 43211 12733 43220 12767
rect 43168 12724 43220 12733
rect 43352 12724 43404 12776
rect 39948 12631 40000 12640
rect 39948 12597 39957 12631
rect 39957 12597 39991 12631
rect 39991 12597 40000 12631
rect 39948 12588 40000 12597
rect 40500 12588 40552 12640
rect 41512 12656 41564 12708
rect 50068 12656 50120 12708
rect 41788 12588 41840 12640
rect 42892 12588 42944 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10048 12384 10100 12436
rect 12900 12384 12952 12436
rect 14004 12384 14056 12436
rect 14556 12384 14608 12436
rect 17960 12384 18012 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 10692 12316 10744 12368
rect 11980 12316 12032 12368
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 1860 12223 1912 12232
rect 1860 12189 1869 12223
rect 1869 12189 1903 12223
rect 1903 12189 1912 12223
rect 1860 12180 1912 12189
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 13452 12180 13504 12232
rect 12440 12155 12492 12164
rect 12440 12121 12449 12155
rect 12449 12121 12483 12155
rect 12483 12121 12492 12155
rect 12440 12112 12492 12121
rect 12624 12155 12676 12164
rect 12624 12121 12649 12155
rect 12649 12121 12676 12155
rect 12624 12112 12676 12121
rect 12992 12112 13044 12164
rect 14556 12291 14608 12300
rect 14556 12257 14565 12291
rect 14565 12257 14599 12291
rect 14599 12257 14608 12291
rect 14556 12248 14608 12257
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 14832 12291 14884 12300
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 15384 12291 15436 12300
rect 14832 12248 14884 12257
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 15936 12248 15988 12300
rect 16304 12248 16356 12300
rect 17224 12248 17276 12300
rect 21272 12384 21324 12436
rect 24584 12384 24636 12436
rect 20720 12316 20772 12368
rect 32220 12384 32272 12436
rect 33232 12384 33284 12436
rect 34060 12384 34112 12436
rect 36084 12384 36136 12436
rect 36544 12384 36596 12436
rect 39120 12427 39172 12436
rect 28724 12316 28776 12368
rect 23480 12248 23532 12300
rect 29368 12248 29420 12300
rect 31576 12248 31628 12300
rect 31668 12248 31720 12300
rect 33784 12248 33836 12300
rect 34060 12248 34112 12300
rect 15016 12180 15068 12232
rect 15108 12180 15160 12232
rect 16488 12180 16540 12232
rect 16856 12180 16908 12232
rect 19248 12180 19300 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 15200 12112 15252 12164
rect 15476 12112 15528 12164
rect 13820 12044 13872 12096
rect 15844 12044 15896 12096
rect 16120 12044 16172 12096
rect 16304 12112 16356 12164
rect 20260 12112 20312 12164
rect 24584 12223 24636 12232
rect 22008 12112 22060 12164
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 25136 12180 25188 12232
rect 29828 12180 29880 12232
rect 31024 12180 31076 12232
rect 33416 12180 33468 12232
rect 33876 12180 33928 12232
rect 34244 12180 34296 12232
rect 27344 12112 27396 12164
rect 29920 12112 29972 12164
rect 30012 12112 30064 12164
rect 20444 12044 20496 12096
rect 23112 12044 23164 12096
rect 27712 12044 27764 12096
rect 29184 12044 29236 12096
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 31484 12044 31536 12096
rect 31944 12044 31996 12096
rect 32496 12087 32548 12096
rect 32496 12053 32505 12087
rect 32505 12053 32539 12087
rect 32539 12053 32548 12087
rect 32496 12044 32548 12053
rect 32956 12112 33008 12164
rect 35164 12316 35216 12368
rect 35440 12316 35492 12368
rect 35532 12316 35584 12368
rect 36268 12316 36320 12368
rect 37280 12316 37332 12368
rect 37648 12316 37700 12368
rect 34520 12248 34572 12300
rect 35440 12180 35492 12232
rect 35624 12291 35676 12300
rect 35624 12257 35633 12291
rect 35633 12257 35667 12291
rect 35667 12257 35676 12291
rect 35624 12248 35676 12257
rect 36084 12248 36136 12300
rect 35716 12223 35768 12232
rect 35716 12189 35725 12223
rect 35725 12189 35759 12223
rect 35759 12189 35768 12223
rect 35716 12180 35768 12189
rect 35808 12180 35860 12232
rect 38016 12291 38068 12300
rect 38016 12257 38025 12291
rect 38025 12257 38059 12291
rect 38059 12257 38068 12291
rect 38016 12248 38068 12257
rect 39120 12393 39129 12427
rect 39129 12393 39163 12427
rect 39163 12393 39172 12427
rect 39120 12384 39172 12393
rect 41420 12384 41472 12436
rect 43628 12384 43680 12436
rect 36452 12180 36504 12232
rect 37924 12223 37976 12232
rect 37924 12189 37933 12223
rect 37933 12189 37967 12223
rect 37967 12189 37976 12223
rect 37924 12180 37976 12189
rect 38108 12180 38160 12232
rect 38844 12223 38896 12232
rect 38844 12189 38853 12223
rect 38853 12189 38887 12223
rect 38887 12189 38896 12223
rect 38844 12180 38896 12189
rect 39764 12180 39816 12232
rect 34888 12044 34940 12096
rect 35072 12087 35124 12096
rect 35072 12053 35081 12087
rect 35081 12053 35115 12087
rect 35115 12053 35124 12087
rect 35072 12044 35124 12053
rect 35256 12087 35308 12096
rect 35256 12053 35265 12087
rect 35265 12053 35299 12087
rect 35299 12053 35308 12087
rect 35256 12044 35308 12053
rect 41052 12112 41104 12164
rect 39580 12044 39632 12096
rect 40132 12044 40184 12096
rect 40868 12044 40920 12096
rect 42708 12248 42760 12300
rect 41788 12223 41840 12232
rect 41788 12189 41797 12223
rect 41797 12189 41831 12223
rect 41831 12189 41840 12223
rect 41788 12180 41840 12189
rect 57520 12180 57572 12232
rect 46204 12112 46256 12164
rect 58164 12155 58216 12164
rect 58164 12121 58173 12155
rect 58173 12121 58207 12155
rect 58207 12121 58216 12155
rect 58164 12112 58216 12121
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 7564 11840 7616 11892
rect 11704 11772 11756 11824
rect 12256 11840 12308 11892
rect 15292 11883 15344 11892
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 11612 11704 11664 11756
rect 14740 11772 14792 11824
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 17040 11883 17092 11892
rect 17040 11849 17049 11883
rect 17049 11849 17083 11883
rect 17083 11849 17092 11883
rect 17040 11840 17092 11849
rect 17224 11840 17276 11892
rect 15016 11772 15068 11824
rect 15476 11704 15528 11756
rect 11796 11568 11848 11620
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 13912 11636 13964 11688
rect 15384 11636 15436 11688
rect 14188 11611 14240 11620
rect 14188 11577 14197 11611
rect 14197 11577 14231 11611
rect 14231 11577 14240 11611
rect 14188 11568 14240 11577
rect 15568 11568 15620 11620
rect 18052 11772 18104 11824
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 16580 11704 16632 11756
rect 16948 11747 17000 11756
rect 16948 11713 16990 11747
rect 16990 11713 17000 11747
rect 16948 11704 17000 11713
rect 17408 11704 17460 11756
rect 17316 11636 17368 11688
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 19340 11772 19392 11824
rect 20260 11840 20312 11892
rect 20444 11840 20496 11892
rect 23112 11840 23164 11892
rect 24032 11840 24084 11892
rect 24216 11840 24268 11892
rect 26516 11840 26568 11892
rect 27436 11840 27488 11892
rect 27712 11840 27764 11892
rect 21272 11772 21324 11824
rect 21824 11772 21876 11824
rect 18788 11704 18840 11756
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 19248 11704 19300 11756
rect 21364 11704 21416 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 22284 11747 22336 11756
rect 22284 11713 22307 11747
rect 22307 11713 22336 11747
rect 22284 11704 22336 11713
rect 26148 11772 26200 11824
rect 27344 11772 27396 11824
rect 29184 11840 29236 11892
rect 30012 11840 30064 11892
rect 30932 11840 30984 11892
rect 31300 11840 31352 11892
rect 33324 11840 33376 11892
rect 33416 11840 33468 11892
rect 34520 11840 34572 11892
rect 35072 11840 35124 11892
rect 30380 11772 30432 11824
rect 32404 11815 32456 11824
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 24492 11704 24544 11756
rect 30564 11704 30616 11756
rect 32404 11781 32413 11815
rect 32413 11781 32447 11815
rect 32447 11781 32456 11815
rect 32404 11772 32456 11781
rect 36176 11772 36228 11824
rect 36820 11772 36872 11824
rect 18604 11636 18656 11688
rect 21916 11636 21968 11688
rect 23112 11636 23164 11688
rect 27620 11636 27672 11688
rect 27804 11636 27856 11688
rect 28080 11679 28132 11688
rect 16396 11568 16448 11620
rect 17868 11568 17920 11620
rect 18696 11568 18748 11620
rect 18788 11568 18840 11620
rect 20444 11568 20496 11620
rect 24308 11568 24360 11620
rect 28080 11645 28089 11679
rect 28089 11645 28123 11679
rect 28123 11645 28132 11679
rect 28080 11636 28132 11645
rect 29184 11636 29236 11688
rect 31300 11679 31352 11688
rect 31300 11645 31309 11679
rect 31309 11645 31343 11679
rect 31343 11645 31352 11679
rect 31300 11636 31352 11645
rect 31392 11679 31444 11688
rect 31392 11645 31401 11679
rect 31401 11645 31435 11679
rect 31435 11645 31444 11679
rect 31392 11636 31444 11645
rect 31576 11636 31628 11688
rect 33048 11636 33100 11688
rect 12808 11500 12860 11552
rect 15108 11500 15160 11552
rect 20076 11500 20128 11552
rect 20260 11500 20312 11552
rect 24768 11500 24820 11552
rect 27436 11543 27488 11552
rect 27436 11509 27445 11543
rect 27445 11509 27479 11543
rect 27479 11509 27488 11543
rect 27436 11500 27488 11509
rect 28540 11568 28592 11620
rect 29828 11568 29880 11620
rect 30104 11611 30156 11620
rect 30104 11577 30113 11611
rect 30113 11577 30147 11611
rect 30147 11577 30156 11611
rect 30104 11568 30156 11577
rect 32404 11568 32456 11620
rect 34336 11704 34388 11756
rect 34888 11636 34940 11688
rect 35348 11747 35400 11756
rect 35348 11713 35357 11747
rect 35357 11713 35391 11747
rect 35391 11713 35400 11747
rect 35348 11704 35400 11713
rect 36268 11704 36320 11756
rect 36084 11636 36136 11688
rect 33416 11568 33468 11620
rect 34060 11568 34112 11620
rect 36268 11568 36320 11620
rect 30656 11500 30708 11552
rect 30840 11543 30892 11552
rect 30840 11509 30849 11543
rect 30849 11509 30883 11543
rect 30883 11509 30892 11543
rect 30840 11500 30892 11509
rect 30932 11500 30984 11552
rect 33324 11500 33376 11552
rect 33600 11500 33652 11552
rect 35348 11500 35400 11552
rect 35440 11500 35492 11552
rect 37280 11704 37332 11756
rect 38568 11704 38620 11756
rect 39672 11840 39724 11892
rect 41880 11840 41932 11892
rect 42340 11840 42392 11892
rect 42984 11840 43036 11892
rect 43076 11840 43128 11892
rect 37372 11636 37424 11688
rect 39580 11704 39632 11756
rect 40132 11747 40184 11756
rect 40132 11713 40141 11747
rect 40141 11713 40175 11747
rect 40175 11713 40184 11747
rect 40132 11704 40184 11713
rect 40684 11772 40736 11824
rect 41420 11772 41472 11824
rect 42892 11815 42944 11824
rect 42892 11781 42926 11815
rect 42926 11781 42944 11815
rect 42892 11772 42944 11781
rect 43168 11772 43220 11824
rect 50896 11772 50948 11824
rect 40316 11704 40368 11756
rect 40500 11747 40552 11756
rect 40500 11713 40509 11747
rect 40509 11713 40543 11747
rect 40543 11713 40552 11747
rect 40500 11704 40552 11713
rect 40592 11636 40644 11688
rect 41144 11747 41196 11756
rect 41144 11713 41153 11747
rect 41153 11713 41187 11747
rect 41187 11713 41196 11747
rect 41144 11704 41196 11713
rect 40776 11636 40828 11688
rect 42340 11704 42392 11756
rect 42708 11704 42760 11756
rect 43444 11704 43496 11756
rect 43720 11704 43772 11756
rect 58072 11747 58124 11756
rect 58072 11713 58081 11747
rect 58081 11713 58115 11747
rect 58115 11713 58124 11747
rect 58072 11704 58124 11713
rect 38568 11568 38620 11620
rect 42340 11568 42392 11620
rect 38752 11500 38804 11552
rect 38844 11543 38896 11552
rect 38844 11509 38853 11543
rect 38853 11509 38887 11543
rect 38887 11509 38896 11543
rect 38844 11500 38896 11509
rect 42616 11500 42668 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12808 11296 12860 11348
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 16764 11296 16816 11348
rect 17500 11296 17552 11348
rect 18880 11339 18932 11348
rect 18880 11305 18889 11339
rect 18889 11305 18923 11339
rect 18923 11305 18932 11339
rect 18880 11296 18932 11305
rect 12256 11160 12308 11212
rect 27252 11296 27304 11348
rect 27436 11296 27488 11348
rect 37188 11296 37240 11348
rect 37372 11339 37424 11348
rect 37372 11305 37381 11339
rect 37381 11305 37415 11339
rect 37415 11305 37424 11339
rect 37372 11296 37424 11305
rect 37740 11296 37792 11348
rect 39396 11296 39448 11348
rect 7564 11092 7616 11144
rect 12072 11092 12124 11144
rect 12624 11092 12676 11144
rect 13544 11160 13596 11212
rect 14556 11160 14608 11212
rect 16304 11160 16356 11212
rect 18328 11160 18380 11212
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 14832 11024 14884 11076
rect 15292 11092 15344 11144
rect 16212 11092 16264 11144
rect 20260 11160 20312 11212
rect 18880 11092 18932 11144
rect 19432 11092 19484 11144
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 21732 11228 21784 11280
rect 24492 11228 24544 11280
rect 27620 11271 27672 11280
rect 27620 11237 27629 11271
rect 27629 11237 27663 11271
rect 27663 11237 27672 11271
rect 27620 11228 27672 11237
rect 21088 11092 21140 11144
rect 22100 11160 22152 11212
rect 25596 11160 25648 11212
rect 27528 11160 27580 11212
rect 30012 11228 30064 11280
rect 33324 11228 33376 11280
rect 33508 11228 33560 11280
rect 33876 11228 33928 11280
rect 36728 11228 36780 11280
rect 28264 11160 28316 11212
rect 28724 11160 28776 11212
rect 33784 11160 33836 11212
rect 34796 11160 34848 11212
rect 21548 11092 21600 11144
rect 15384 11024 15436 11076
rect 17224 11024 17276 11076
rect 21916 11024 21968 11076
rect 22192 11092 22244 11144
rect 24492 11092 24544 11144
rect 25228 11092 25280 11144
rect 28908 11092 28960 11144
rect 30104 11092 30156 11144
rect 31024 11092 31076 11144
rect 32312 11092 32364 11144
rect 33324 11092 33376 11144
rect 34428 11092 34480 11144
rect 14740 10956 14792 11008
rect 17040 10956 17092 11008
rect 24952 11024 25004 11076
rect 29092 11024 29144 11076
rect 35808 11160 35860 11212
rect 37096 11228 37148 11280
rect 37280 11228 37332 11280
rect 38016 11228 38068 11280
rect 38844 11228 38896 11280
rect 36912 11092 36964 11144
rect 26608 10956 26660 11008
rect 29368 10956 29420 11008
rect 30656 10956 30708 11008
rect 31116 10956 31168 11008
rect 32680 10956 32732 11008
rect 32956 10956 33008 11008
rect 33324 10956 33376 11008
rect 34520 10956 34572 11008
rect 36728 11024 36780 11076
rect 35992 10956 36044 11008
rect 38292 11160 38344 11212
rect 37188 11135 37240 11144
rect 37188 11101 37197 11135
rect 37197 11101 37231 11135
rect 37231 11101 37240 11135
rect 37188 11092 37240 11101
rect 38016 11135 38068 11144
rect 38016 11101 38025 11135
rect 38025 11101 38059 11135
rect 38059 11101 38068 11135
rect 38016 11092 38068 11101
rect 38752 11092 38804 11144
rect 40684 11228 40736 11280
rect 43628 11228 43680 11280
rect 38936 11024 38988 11076
rect 41144 11160 41196 11212
rect 40776 11135 40828 11144
rect 40776 11101 40785 11135
rect 40785 11101 40819 11135
rect 40819 11101 40828 11135
rect 40776 11092 40828 11101
rect 52460 11160 52512 11212
rect 43168 11092 43220 11144
rect 43260 11092 43312 11144
rect 44088 11135 44140 11144
rect 44088 11101 44097 11135
rect 44097 11101 44131 11135
rect 44131 11101 44140 11135
rect 44088 11092 44140 11101
rect 54208 11228 54260 11280
rect 52736 11160 52788 11212
rect 54484 11160 54536 11212
rect 43444 11067 43496 11076
rect 43444 11033 43453 11067
rect 43453 11033 43487 11067
rect 43487 11033 43496 11067
rect 43444 11024 43496 11033
rect 43628 11024 43680 11076
rect 52828 11135 52880 11144
rect 52828 11101 52837 11135
rect 52837 11101 52871 11135
rect 52871 11101 52880 11135
rect 52828 11092 52880 11101
rect 53012 11135 53064 11144
rect 53012 11101 53021 11135
rect 53021 11101 53055 11135
rect 53055 11101 53064 11135
rect 53012 11092 53064 11101
rect 46204 11024 46256 11076
rect 50620 11024 50672 11076
rect 53104 11024 53156 11076
rect 37188 10956 37240 11008
rect 37372 10956 37424 11008
rect 57888 10956 57940 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 7564 10752 7616 10804
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 14096 10727 14148 10736
rect 14096 10693 14121 10727
rect 14121 10693 14148 10727
rect 14096 10684 14148 10693
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 13084 10616 13136 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 14832 10752 14884 10804
rect 15016 10752 15068 10804
rect 15384 10752 15436 10804
rect 15476 10752 15528 10804
rect 19156 10752 19208 10804
rect 22376 10752 22428 10804
rect 22836 10752 22888 10804
rect 29092 10795 29144 10804
rect 29092 10761 29101 10795
rect 29101 10761 29135 10795
rect 29135 10761 29144 10795
rect 29092 10752 29144 10761
rect 29368 10752 29420 10804
rect 30564 10752 30616 10804
rect 14280 10616 14332 10668
rect 14832 10616 14884 10668
rect 15200 10616 15252 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15752 10659 15804 10668
rect 15292 10616 15344 10625
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 15844 10616 15896 10668
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16856 10659 16908 10668
rect 16120 10616 16172 10625
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 16212 10548 16264 10600
rect 17040 10548 17092 10600
rect 20076 10684 20128 10736
rect 20904 10684 20956 10736
rect 21272 10684 21324 10736
rect 18328 10616 18380 10668
rect 18972 10616 19024 10668
rect 19524 10616 19576 10668
rect 20812 10616 20864 10668
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 22652 10616 22704 10668
rect 18420 10548 18472 10600
rect 19708 10548 19760 10600
rect 20076 10548 20128 10600
rect 22284 10548 22336 10600
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 15200 10412 15252 10464
rect 16212 10412 16264 10464
rect 17316 10412 17368 10464
rect 17592 10455 17644 10464
rect 17592 10421 17601 10455
rect 17601 10421 17635 10455
rect 17635 10421 17644 10455
rect 17592 10412 17644 10421
rect 23480 10480 23532 10532
rect 24032 10684 24084 10736
rect 31116 10752 31168 10804
rect 31300 10795 31352 10804
rect 31300 10761 31309 10795
rect 31309 10761 31343 10795
rect 31343 10761 31352 10795
rect 31300 10752 31352 10761
rect 32404 10752 32456 10804
rect 33968 10752 34020 10804
rect 34336 10752 34388 10804
rect 25044 10616 25096 10668
rect 27620 10616 27672 10668
rect 28172 10616 28224 10668
rect 32864 10684 32916 10736
rect 33140 10727 33192 10736
rect 33140 10693 33149 10727
rect 33149 10693 33183 10727
rect 33183 10693 33192 10727
rect 33140 10684 33192 10693
rect 30564 10616 30616 10668
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 32588 10616 32640 10625
rect 33784 10616 33836 10668
rect 33968 10659 34020 10668
rect 33968 10625 33977 10659
rect 33977 10625 34011 10659
rect 34011 10625 34020 10659
rect 33968 10616 34020 10625
rect 34520 10684 34572 10736
rect 34704 10752 34756 10804
rect 36452 10752 36504 10804
rect 36728 10752 36780 10804
rect 37648 10752 37700 10804
rect 38476 10752 38528 10804
rect 40960 10752 41012 10804
rect 41144 10752 41196 10804
rect 42340 10752 42392 10804
rect 46296 10752 46348 10804
rect 49700 10752 49752 10804
rect 56876 10752 56928 10804
rect 24952 10548 25004 10600
rect 26332 10548 26384 10600
rect 31576 10548 31628 10600
rect 30104 10480 30156 10532
rect 30656 10480 30708 10532
rect 31760 10480 31812 10532
rect 32588 10480 32640 10532
rect 34520 10548 34572 10600
rect 34060 10480 34112 10532
rect 20352 10455 20404 10464
rect 20352 10421 20361 10455
rect 20361 10421 20395 10455
rect 20395 10421 20404 10455
rect 20352 10412 20404 10421
rect 20720 10412 20772 10464
rect 22284 10412 22336 10464
rect 24768 10412 24820 10464
rect 27160 10412 27212 10464
rect 28724 10412 28776 10464
rect 35532 10616 35584 10668
rect 35624 10616 35676 10668
rect 36268 10659 36320 10668
rect 36268 10625 36277 10659
rect 36277 10625 36311 10659
rect 36311 10625 36320 10659
rect 36268 10616 36320 10625
rect 38660 10659 38712 10668
rect 35808 10548 35860 10600
rect 35900 10548 35952 10600
rect 36176 10548 36228 10600
rect 35624 10480 35676 10532
rect 37372 10548 37424 10600
rect 35808 10412 35860 10464
rect 36912 10480 36964 10532
rect 38660 10625 38669 10659
rect 38669 10625 38703 10659
rect 38703 10625 38712 10659
rect 38660 10616 38712 10625
rect 38752 10616 38804 10668
rect 39580 10616 39632 10668
rect 37924 10591 37976 10600
rect 37924 10557 37933 10591
rect 37933 10557 37967 10591
rect 37967 10557 37976 10591
rect 37924 10548 37976 10557
rect 40592 10659 40644 10668
rect 40592 10625 40601 10659
rect 40601 10625 40635 10659
rect 40635 10625 40644 10659
rect 40592 10616 40644 10625
rect 40868 10659 40920 10668
rect 38936 10523 38988 10532
rect 36452 10455 36504 10464
rect 36452 10421 36461 10455
rect 36461 10421 36495 10455
rect 36495 10421 36504 10455
rect 36452 10412 36504 10421
rect 37372 10412 37424 10464
rect 38936 10489 38945 10523
rect 38945 10489 38979 10523
rect 38979 10489 38988 10523
rect 38936 10480 38988 10489
rect 40868 10625 40877 10659
rect 40877 10625 40911 10659
rect 40911 10625 40920 10659
rect 40868 10616 40920 10625
rect 40960 10659 41012 10668
rect 40960 10625 40969 10659
rect 40969 10625 41003 10659
rect 41003 10625 41012 10659
rect 41604 10684 41656 10736
rect 43260 10684 43312 10736
rect 43444 10684 43496 10736
rect 47216 10684 47268 10736
rect 49516 10684 49568 10736
rect 53288 10684 53340 10736
rect 40960 10616 41012 10625
rect 42800 10616 42852 10668
rect 57244 10659 57296 10668
rect 43352 10548 43404 10600
rect 57244 10625 57253 10659
rect 57253 10625 57287 10659
rect 57287 10625 57296 10659
rect 57244 10616 57296 10625
rect 57520 10616 57572 10668
rect 52000 10548 52052 10600
rect 40316 10412 40368 10464
rect 40500 10412 40552 10464
rect 40776 10412 40828 10464
rect 41328 10412 41380 10464
rect 41788 10455 41840 10464
rect 41788 10421 41797 10455
rect 41797 10421 41831 10455
rect 41831 10421 41840 10455
rect 41788 10412 41840 10421
rect 42064 10412 42116 10464
rect 42892 10412 42944 10464
rect 45468 10455 45520 10464
rect 45468 10421 45477 10455
rect 45477 10421 45511 10455
rect 45511 10421 45520 10455
rect 45468 10412 45520 10421
rect 46296 10480 46348 10532
rect 58256 10480 58308 10532
rect 51724 10412 51776 10464
rect 57336 10455 57388 10464
rect 57336 10421 57345 10455
rect 57345 10421 57379 10455
rect 57379 10421 57388 10455
rect 57336 10412 57388 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1952 10208 2004 10260
rect 7564 10208 7616 10260
rect 11888 10208 11940 10260
rect 16028 10208 16080 10260
rect 16120 10208 16172 10260
rect 24032 10208 24084 10260
rect 24400 10208 24452 10260
rect 24676 10251 24728 10260
rect 24676 10217 24685 10251
rect 24685 10217 24719 10251
rect 24719 10217 24728 10251
rect 24676 10208 24728 10217
rect 24952 10208 25004 10260
rect 25320 10208 25372 10260
rect 25504 10208 25556 10260
rect 7656 10140 7708 10192
rect 12348 10140 12400 10192
rect 14740 10140 14792 10192
rect 11796 10072 11848 10124
rect 12532 10072 12584 10124
rect 13820 10004 13872 10056
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 20352 10140 20404 10192
rect 20812 10140 20864 10192
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16948 10047 17000 10056
rect 13728 9936 13780 9988
rect 16028 9936 16080 9988
rect 16488 9979 16540 9988
rect 16488 9945 16497 9979
rect 16497 9945 16531 9979
rect 16531 9945 16540 9979
rect 16488 9936 16540 9945
rect 14096 9868 14148 9920
rect 16672 9868 16724 9920
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 17776 10072 17828 10124
rect 17868 10072 17920 10124
rect 17684 9936 17736 9988
rect 18512 10072 18564 10124
rect 18696 10072 18748 10124
rect 20720 10072 20772 10124
rect 21548 10072 21600 10124
rect 21916 10072 21968 10124
rect 23388 10072 23440 10124
rect 24676 10072 24728 10124
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 28632 10072 28684 10124
rect 33140 10140 33192 10192
rect 35808 10208 35860 10260
rect 34336 10140 34388 10192
rect 35900 10140 35952 10192
rect 18328 10004 18380 10056
rect 19524 10004 19576 10056
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 19800 10004 19852 10056
rect 20536 10004 20588 10056
rect 20904 10004 20956 10056
rect 20444 9936 20496 9988
rect 21272 10004 21324 10056
rect 22100 10047 22152 10056
rect 22100 10013 22109 10047
rect 22109 10013 22143 10047
rect 22143 10013 22152 10047
rect 22100 10004 22152 10013
rect 23112 10004 23164 10056
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 25320 10004 25372 10056
rect 22284 9936 22336 9988
rect 23756 9936 23808 9988
rect 29000 10004 29052 10056
rect 29092 10004 29144 10056
rect 30288 10115 30340 10124
rect 30288 10081 30297 10115
rect 30297 10081 30331 10115
rect 30331 10081 30340 10115
rect 30288 10072 30340 10081
rect 31208 10072 31260 10124
rect 31852 10072 31904 10124
rect 32404 10072 32456 10124
rect 32772 10072 32824 10124
rect 33048 10072 33100 10124
rect 33968 10004 34020 10056
rect 19432 9868 19484 9920
rect 20996 9868 21048 9920
rect 21088 9868 21140 9920
rect 21272 9868 21324 9920
rect 21364 9868 21416 9920
rect 22192 9868 22244 9920
rect 24952 9868 25004 9920
rect 25044 9868 25096 9920
rect 27620 9868 27672 9920
rect 33784 9936 33836 9988
rect 34520 10004 34572 10056
rect 34796 10072 34848 10124
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 35072 10047 35124 10056
rect 35072 10013 35081 10047
rect 35081 10013 35115 10047
rect 35115 10013 35124 10047
rect 35072 10004 35124 10013
rect 35256 10047 35308 10056
rect 35256 10013 35265 10047
rect 35265 10013 35299 10047
rect 35299 10013 35308 10047
rect 49516 10208 49568 10260
rect 57520 10208 57572 10260
rect 36268 10140 36320 10192
rect 38108 10140 38160 10192
rect 39212 10140 39264 10192
rect 40408 10140 40460 10192
rect 35256 10004 35308 10013
rect 36176 10047 36228 10056
rect 36176 10013 36185 10047
rect 36185 10013 36219 10047
rect 36219 10013 36228 10047
rect 36176 10004 36228 10013
rect 36636 10072 36688 10124
rect 37096 10047 37148 10056
rect 37096 10013 37105 10047
rect 37105 10013 37139 10047
rect 37139 10013 37148 10047
rect 37096 10004 37148 10013
rect 37372 10047 37424 10056
rect 37372 10013 37406 10047
rect 37406 10013 37424 10047
rect 37372 10004 37424 10013
rect 38660 10004 38712 10056
rect 39948 10004 40000 10056
rect 40040 10004 40092 10056
rect 40684 10047 40736 10056
rect 40684 10013 40693 10047
rect 40693 10013 40727 10047
rect 40727 10013 40736 10047
rect 40684 10004 40736 10013
rect 40776 10047 40828 10056
rect 40776 10013 40790 10047
rect 40790 10013 40824 10047
rect 40824 10013 40828 10047
rect 40776 10004 40828 10013
rect 36452 9936 36504 9988
rect 39120 9979 39172 9988
rect 39120 9945 39129 9979
rect 39129 9945 39163 9979
rect 39163 9945 39172 9979
rect 39120 9936 39172 9945
rect 39212 9936 39264 9988
rect 32680 9868 32732 9920
rect 34796 9868 34848 9920
rect 37924 9868 37976 9920
rect 38660 9868 38712 9920
rect 41052 9936 41104 9988
rect 42708 10072 42760 10124
rect 43168 10072 43220 10124
rect 43352 10072 43404 10124
rect 56876 10115 56928 10124
rect 56876 10081 56885 10115
rect 56885 10081 56919 10115
rect 56919 10081 56928 10115
rect 56876 10072 56928 10081
rect 43628 10004 43680 10056
rect 41420 9868 41472 9920
rect 42800 9936 42852 9988
rect 45100 9936 45152 9988
rect 56784 9936 56836 9988
rect 45192 9868 45244 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 16948 9664 17000 9716
rect 17776 9664 17828 9716
rect 14372 9596 14424 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 11980 9528 12032 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 17224 9596 17276 9648
rect 16396 9528 16448 9580
rect 17132 9528 17184 9580
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 16304 9503 16356 9512
rect 15844 9460 15896 9469
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 17592 9460 17644 9512
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 22560 9664 22612 9716
rect 18880 9596 18932 9648
rect 20812 9596 20864 9648
rect 20904 9596 20956 9648
rect 24952 9664 25004 9716
rect 26608 9664 26660 9716
rect 26700 9664 26752 9716
rect 28632 9664 28684 9716
rect 29000 9707 29052 9716
rect 29000 9673 29009 9707
rect 29009 9673 29043 9707
rect 29043 9673 29052 9707
rect 29000 9664 29052 9673
rect 29736 9664 29788 9716
rect 30288 9664 30340 9716
rect 30472 9664 30524 9716
rect 30932 9664 30984 9716
rect 32404 9664 32456 9716
rect 32680 9707 32732 9716
rect 32680 9673 32689 9707
rect 32689 9673 32723 9707
rect 32723 9673 32732 9707
rect 32680 9664 32732 9673
rect 32956 9664 33008 9716
rect 34796 9664 34848 9716
rect 34888 9664 34940 9716
rect 25044 9596 25096 9648
rect 25872 9596 25924 9648
rect 27620 9596 27672 9648
rect 29460 9639 29512 9648
rect 29460 9605 29469 9639
rect 29469 9605 29503 9639
rect 29503 9605 29512 9639
rect 29460 9596 29512 9605
rect 29644 9596 29696 9648
rect 31116 9596 31168 9648
rect 18144 9528 18196 9537
rect 18972 9528 19024 9580
rect 19708 9528 19760 9580
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 20628 9571 20680 9580
rect 18328 9460 18380 9512
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 21364 9528 21416 9580
rect 21916 9528 21968 9580
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 24216 9528 24268 9580
rect 25596 9571 25648 9580
rect 20904 9460 20956 9512
rect 22100 9460 22152 9512
rect 22744 9460 22796 9512
rect 23388 9460 23440 9512
rect 25596 9537 25605 9571
rect 25605 9537 25639 9571
rect 25639 9537 25648 9571
rect 25596 9528 25648 9537
rect 5816 9392 5868 9444
rect 12072 9392 12124 9444
rect 16396 9392 16448 9444
rect 20720 9392 20772 9444
rect 20812 9392 20864 9444
rect 23664 9392 23716 9444
rect 25044 9460 25096 9512
rect 25136 9460 25188 9512
rect 25872 9460 25924 9512
rect 26056 9528 26108 9580
rect 27436 9528 27488 9580
rect 26424 9503 26476 9512
rect 26424 9469 26433 9503
rect 26433 9469 26467 9503
rect 26467 9469 26476 9503
rect 26424 9460 26476 9469
rect 26148 9392 26200 9444
rect 26976 9460 27028 9512
rect 28264 9460 28316 9512
rect 27436 9392 27488 9444
rect 10876 9324 10928 9376
rect 14924 9324 14976 9376
rect 16764 9324 16816 9376
rect 16856 9324 16908 9376
rect 18880 9324 18932 9376
rect 18972 9324 19024 9376
rect 19892 9324 19944 9376
rect 21364 9324 21416 9376
rect 24492 9324 24544 9376
rect 25136 9324 25188 9376
rect 25780 9324 25832 9376
rect 29000 9528 29052 9580
rect 30288 9528 30340 9580
rect 31024 9528 31076 9580
rect 31208 9571 31260 9580
rect 31208 9537 31217 9571
rect 31217 9537 31251 9571
rect 31251 9537 31260 9571
rect 31208 9528 31260 9537
rect 31576 9528 31628 9580
rect 31760 9571 31812 9580
rect 31760 9537 31767 9571
rect 31767 9537 31801 9571
rect 31801 9537 31812 9571
rect 33784 9596 33836 9648
rect 34244 9596 34296 9648
rect 35072 9596 35124 9648
rect 31760 9528 31812 9537
rect 32772 9571 32824 9580
rect 32772 9537 32781 9571
rect 32781 9537 32815 9571
rect 32815 9537 32824 9571
rect 32772 9528 32824 9537
rect 33416 9528 33468 9580
rect 33876 9571 33928 9580
rect 33876 9537 33885 9571
rect 33885 9537 33919 9571
rect 33919 9537 33928 9571
rect 33876 9528 33928 9537
rect 34060 9571 34112 9580
rect 34060 9537 34069 9571
rect 34069 9537 34103 9571
rect 34103 9537 34112 9571
rect 34060 9528 34112 9537
rect 34612 9528 34664 9580
rect 34888 9528 34940 9580
rect 35440 9528 35492 9580
rect 28540 9460 28592 9512
rect 29828 9392 29880 9444
rect 33968 9460 34020 9512
rect 34336 9460 34388 9512
rect 35808 9528 35860 9580
rect 36084 9571 36136 9580
rect 36084 9537 36093 9571
rect 36093 9537 36127 9571
rect 36127 9537 36136 9571
rect 36084 9528 36136 9537
rect 36544 9528 36596 9580
rect 36636 9528 36688 9580
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 39304 9596 39356 9648
rect 39856 9596 39908 9648
rect 40960 9664 41012 9716
rect 41880 9664 41932 9716
rect 43352 9664 43404 9716
rect 57336 9664 57388 9716
rect 58256 9707 58308 9716
rect 58256 9673 58265 9707
rect 58265 9673 58299 9707
rect 58299 9673 58308 9707
rect 58256 9664 58308 9673
rect 42892 9639 42944 9648
rect 42892 9605 42926 9639
rect 42926 9605 42944 9639
rect 44916 9639 44968 9648
rect 42892 9596 42944 9605
rect 44916 9605 44925 9639
rect 44925 9605 44959 9639
rect 44959 9605 44968 9639
rect 44916 9596 44968 9605
rect 37832 9571 37884 9580
rect 37832 9537 37841 9571
rect 37841 9537 37875 9571
rect 37875 9537 37884 9571
rect 37832 9528 37884 9537
rect 38660 9528 38712 9580
rect 38936 9571 38988 9580
rect 38936 9537 38945 9571
rect 38945 9537 38979 9571
rect 38979 9537 38988 9571
rect 38936 9528 38988 9537
rect 31300 9392 31352 9444
rect 31576 9392 31628 9444
rect 32956 9392 33008 9444
rect 31944 9324 31996 9376
rect 32128 9324 32180 9376
rect 33692 9324 33744 9376
rect 34980 9367 35032 9376
rect 34980 9333 34989 9367
rect 34989 9333 35023 9367
rect 35023 9333 35032 9367
rect 34980 9324 35032 9333
rect 35440 9392 35492 9444
rect 35992 9392 36044 9444
rect 35624 9324 35676 9376
rect 35808 9324 35860 9376
rect 38660 9324 38712 9376
rect 39764 9571 39816 9580
rect 39764 9537 39774 9571
rect 39774 9537 39808 9571
rect 39808 9537 39816 9571
rect 39764 9528 39816 9537
rect 39672 9392 39724 9444
rect 39856 9460 39908 9512
rect 40500 9528 40552 9580
rect 40776 9528 40828 9580
rect 41420 9571 41472 9580
rect 41420 9537 41429 9571
rect 41429 9537 41463 9571
rect 41463 9537 41472 9571
rect 41420 9528 41472 9537
rect 40316 9460 40368 9512
rect 40040 9392 40092 9444
rect 41604 9460 41656 9512
rect 42248 9392 42300 9444
rect 40776 9324 40828 9376
rect 40960 9324 41012 9376
rect 41236 9324 41288 9376
rect 42708 9528 42760 9580
rect 56692 9528 56744 9580
rect 58072 9571 58124 9580
rect 43996 9460 44048 9512
rect 45100 9503 45152 9512
rect 45100 9469 45109 9503
rect 45109 9469 45143 9503
rect 45143 9469 45152 9503
rect 45100 9460 45152 9469
rect 55404 9460 55456 9512
rect 58072 9537 58081 9571
rect 58081 9537 58115 9571
rect 58115 9537 58124 9571
rect 58072 9528 58124 9537
rect 44732 9392 44784 9444
rect 56784 9435 56836 9444
rect 56784 9401 56793 9435
rect 56793 9401 56827 9435
rect 56827 9401 56836 9435
rect 56784 9392 56836 9401
rect 44548 9367 44600 9376
rect 44548 9333 44557 9367
rect 44557 9333 44591 9367
rect 44591 9333 44600 9367
rect 44548 9324 44600 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 14832 9120 14884 9172
rect 16856 9120 16908 9172
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 18696 9120 18748 9172
rect 18972 9120 19024 9172
rect 19340 9120 19392 9172
rect 21548 9120 21600 9172
rect 15016 9052 15068 9104
rect 15844 9052 15896 9104
rect 17960 9052 18012 9104
rect 19064 9052 19116 9104
rect 13728 8916 13780 8968
rect 18052 8984 18104 9036
rect 16396 8916 16448 8968
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 16212 8848 16264 8900
rect 17592 8916 17644 8968
rect 17408 8848 17460 8900
rect 17684 8848 17736 8900
rect 18328 8916 18380 8968
rect 18972 8984 19024 9036
rect 18604 8925 18609 8946
rect 18609 8925 18643 8946
rect 18643 8925 18656 8946
rect 13728 8780 13780 8832
rect 13912 8780 13964 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 16396 8780 16448 8832
rect 18236 8848 18288 8900
rect 18604 8894 18656 8925
rect 19340 8916 19392 8968
rect 20352 8984 20404 9036
rect 19800 8959 19852 8968
rect 19800 8925 19809 8959
rect 19809 8925 19843 8959
rect 19843 8925 19852 8959
rect 19800 8916 19852 8925
rect 20628 8984 20680 9036
rect 21916 8984 21968 9036
rect 22100 8916 22152 8968
rect 22468 8916 22520 8968
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 18788 8848 18840 8900
rect 19708 8891 19760 8900
rect 19708 8857 19717 8891
rect 19717 8857 19751 8891
rect 19751 8857 19760 8891
rect 19708 8848 19760 8857
rect 19064 8780 19116 8832
rect 20444 8848 20496 8900
rect 20904 8848 20956 8900
rect 20352 8823 20404 8832
rect 20352 8789 20361 8823
rect 20361 8789 20395 8823
rect 20395 8789 20404 8823
rect 20352 8780 20404 8789
rect 20812 8780 20864 8832
rect 22100 8780 22152 8832
rect 22284 8780 22336 8832
rect 23940 9120 23992 9172
rect 24952 9120 25004 9172
rect 26608 9163 26660 9172
rect 26608 9129 26617 9163
rect 26617 9129 26651 9163
rect 26651 9129 26660 9163
rect 26608 9120 26660 9129
rect 27436 9120 27488 9172
rect 32772 9120 32824 9172
rect 32956 9120 33008 9172
rect 33600 9120 33652 9172
rect 33876 9120 33928 9172
rect 37832 9120 37884 9172
rect 39120 9120 39172 9172
rect 26976 9052 27028 9104
rect 28172 9052 28224 9104
rect 30748 9052 30800 9104
rect 31760 9052 31812 9104
rect 32680 9052 32732 9104
rect 25228 9027 25280 9036
rect 25228 8993 25237 9027
rect 25237 8993 25271 9027
rect 25271 8993 25280 9027
rect 25228 8984 25280 8993
rect 26424 8984 26476 9036
rect 32956 9027 33008 9036
rect 23940 8916 23992 8968
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 27160 8916 27212 8968
rect 32956 8993 32965 9027
rect 32965 8993 32999 9027
rect 32999 8993 33008 9027
rect 32956 8984 33008 8993
rect 33416 9052 33468 9104
rect 35808 9052 35860 9104
rect 37188 9052 37240 9104
rect 41420 9052 41472 9104
rect 43996 9095 44048 9104
rect 43996 9061 44005 9095
rect 44005 9061 44039 9095
rect 44039 9061 44048 9095
rect 43996 9052 44048 9061
rect 28724 8916 28776 8968
rect 29092 8916 29144 8968
rect 26700 8780 26752 8832
rect 28356 8848 28408 8900
rect 28908 8848 28960 8900
rect 29644 8916 29696 8968
rect 29828 8959 29880 8968
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 30748 8959 30800 8968
rect 29828 8916 29880 8925
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 31392 8916 31444 8968
rect 33508 8916 33560 8968
rect 33784 8916 33836 8968
rect 29368 8848 29420 8900
rect 29552 8848 29604 8900
rect 37096 8984 37148 9036
rect 37832 8984 37884 9036
rect 39580 8984 39632 9036
rect 40592 8984 40644 9036
rect 41328 8984 41380 9036
rect 41604 8984 41656 9036
rect 34704 8916 34756 8968
rect 34796 8916 34848 8968
rect 34980 8916 35032 8968
rect 35440 8916 35492 8968
rect 35624 8916 35676 8968
rect 35992 8916 36044 8968
rect 38016 8959 38068 8968
rect 37556 8891 37608 8900
rect 30840 8780 30892 8832
rect 31760 8780 31812 8832
rect 34060 8780 34112 8832
rect 37556 8857 37565 8891
rect 37565 8857 37599 8891
rect 37599 8857 37608 8891
rect 37556 8848 37608 8857
rect 35164 8780 35216 8832
rect 35440 8780 35492 8832
rect 37648 8780 37700 8832
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 38108 8959 38160 8968
rect 38108 8925 38118 8959
rect 38118 8925 38152 8959
rect 38152 8925 38160 8959
rect 38384 8959 38436 8968
rect 38108 8916 38160 8925
rect 38384 8925 38393 8959
rect 38393 8925 38427 8959
rect 38427 8925 38436 8959
rect 38384 8916 38436 8925
rect 38476 8959 38528 8968
rect 38476 8925 38490 8959
rect 38490 8925 38524 8959
rect 38524 8925 38528 8959
rect 38476 8916 38528 8925
rect 38936 8916 38988 8968
rect 39764 8916 39816 8968
rect 40408 8916 40460 8968
rect 40684 8916 40736 8968
rect 41144 8916 41196 8968
rect 42708 8916 42760 8968
rect 44548 8916 44600 8968
rect 57152 8916 57204 8968
rect 58256 8916 58308 8968
rect 37924 8848 37976 8900
rect 39120 8891 39172 8900
rect 38844 8780 38896 8832
rect 39120 8857 39129 8891
rect 39129 8857 39163 8891
rect 39163 8857 39172 8891
rect 39120 8848 39172 8857
rect 39580 8848 39632 8900
rect 39856 8848 39908 8900
rect 42984 8848 43036 8900
rect 44088 8848 44140 8900
rect 58164 8891 58216 8900
rect 58164 8857 58173 8891
rect 58173 8857 58207 8891
rect 58207 8857 58216 8891
rect 58164 8848 58216 8857
rect 40684 8780 40736 8832
rect 56600 8780 56652 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 15200 8576 15252 8628
rect 16396 8576 16448 8628
rect 2504 8508 2556 8560
rect 8668 8508 8720 8560
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 13636 8440 13688 8492
rect 17408 8508 17460 8560
rect 10324 8415 10376 8424
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 11244 8372 11296 8424
rect 12072 8372 12124 8424
rect 17132 8440 17184 8492
rect 18604 8576 18656 8628
rect 19248 8576 19300 8628
rect 19340 8576 19392 8628
rect 21456 8619 21508 8628
rect 18788 8508 18840 8560
rect 18328 8440 18380 8492
rect 19340 8440 19392 8492
rect 21456 8585 21465 8619
rect 21465 8585 21499 8619
rect 21499 8585 21508 8619
rect 21456 8576 21508 8585
rect 20076 8508 20128 8560
rect 16672 8372 16724 8424
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 20260 8483 20312 8492
rect 19984 8440 20036 8449
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20812 8508 20864 8560
rect 24952 8576 25004 8628
rect 25412 8576 25464 8628
rect 26976 8576 27028 8628
rect 27068 8576 27120 8628
rect 28356 8619 28408 8628
rect 28356 8585 28365 8619
rect 28365 8585 28399 8619
rect 28399 8585 28408 8619
rect 28356 8576 28408 8585
rect 28448 8576 28500 8628
rect 29092 8576 29144 8628
rect 31300 8576 31352 8628
rect 33232 8619 33284 8628
rect 33232 8585 33241 8619
rect 33241 8585 33275 8619
rect 33275 8585 33284 8619
rect 33232 8576 33284 8585
rect 21824 8440 21876 8492
rect 23756 8483 23808 8492
rect 19800 8372 19852 8424
rect 20996 8372 21048 8424
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 25780 8440 25832 8492
rect 27160 8508 27212 8560
rect 27252 8508 27304 8560
rect 26148 8440 26200 8492
rect 27436 8440 27488 8492
rect 22836 8415 22888 8424
rect 22836 8381 22845 8415
rect 22845 8381 22879 8415
rect 22879 8381 22888 8415
rect 22836 8372 22888 8381
rect 24032 8372 24084 8424
rect 24952 8372 25004 8424
rect 25044 8372 25096 8424
rect 25872 8372 25924 8424
rect 16764 8304 16816 8356
rect 26332 8304 26384 8356
rect 27988 8372 28040 8424
rect 28724 8372 28776 8424
rect 29736 8440 29788 8492
rect 32312 8508 32364 8560
rect 32588 8551 32640 8560
rect 32588 8517 32597 8551
rect 32597 8517 32631 8551
rect 32631 8517 32640 8551
rect 32588 8508 32640 8517
rect 32956 8508 33008 8560
rect 37648 8576 37700 8628
rect 39396 8619 39448 8628
rect 33416 8508 33468 8560
rect 30104 8483 30156 8492
rect 30104 8449 30138 8483
rect 30138 8449 30156 8483
rect 30104 8440 30156 8449
rect 31484 8440 31536 8492
rect 33692 8483 33744 8492
rect 33692 8449 33701 8483
rect 33701 8449 33735 8483
rect 33735 8449 33744 8483
rect 33692 8440 33744 8449
rect 35072 8508 35124 8560
rect 36084 8508 36136 8560
rect 31024 8372 31076 8424
rect 32404 8372 32456 8424
rect 33324 8372 33376 8424
rect 29460 8304 29512 8356
rect 35164 8440 35216 8492
rect 36268 8483 36320 8492
rect 36268 8449 36277 8483
rect 36277 8449 36311 8483
rect 36311 8449 36320 8483
rect 36268 8440 36320 8449
rect 36452 8483 36504 8492
rect 36452 8449 36459 8483
rect 36459 8449 36504 8483
rect 36452 8440 36504 8449
rect 34888 8415 34940 8424
rect 34888 8381 34897 8415
rect 34897 8381 34931 8415
rect 34931 8381 34940 8415
rect 34888 8372 34940 8381
rect 35716 8372 35768 8424
rect 36912 8508 36964 8560
rect 37464 8508 37516 8560
rect 37096 8440 37148 8492
rect 39396 8585 39405 8619
rect 39405 8585 39439 8619
rect 39439 8585 39448 8619
rect 39396 8576 39448 8585
rect 39580 8576 39632 8628
rect 40592 8576 40644 8628
rect 41236 8619 41288 8628
rect 41236 8585 41245 8619
rect 41245 8585 41279 8619
rect 41279 8585 41288 8619
rect 41236 8576 41288 8585
rect 38476 8508 38528 8560
rect 39672 8508 39724 8560
rect 40868 8508 40920 8560
rect 40040 8483 40092 8492
rect 40040 8449 40049 8483
rect 40049 8449 40083 8483
rect 40083 8449 40092 8483
rect 40040 8440 40092 8449
rect 40316 8483 40368 8492
rect 34980 8304 35032 8356
rect 35072 8304 35124 8356
rect 37188 8304 37240 8356
rect 40040 8304 40092 8356
rect 40316 8449 40325 8483
rect 40325 8449 40359 8483
rect 40359 8449 40368 8483
rect 40316 8440 40368 8449
rect 40505 8483 40557 8492
rect 40505 8449 40514 8483
rect 40514 8449 40548 8483
rect 40548 8449 40557 8483
rect 40505 8440 40557 8449
rect 41328 8440 41380 8492
rect 52644 8576 52696 8628
rect 41696 8483 41748 8492
rect 41696 8449 41705 8483
rect 41705 8449 41739 8483
rect 41739 8449 41748 8483
rect 41696 8440 41748 8449
rect 43628 8483 43680 8492
rect 42984 8415 43036 8424
rect 42984 8381 42993 8415
rect 42993 8381 43027 8415
rect 43027 8381 43036 8415
rect 42984 8372 43036 8381
rect 43628 8449 43637 8483
rect 43637 8449 43671 8483
rect 43671 8449 43680 8483
rect 43628 8440 43680 8449
rect 44088 8440 44140 8492
rect 57152 8483 57204 8492
rect 57152 8449 57161 8483
rect 57161 8449 57195 8483
rect 57195 8449 57204 8483
rect 57152 8440 57204 8449
rect 43812 8415 43864 8424
rect 43812 8381 43821 8415
rect 43821 8381 43855 8415
rect 43855 8381 43864 8415
rect 43812 8372 43864 8381
rect 44180 8372 44232 8424
rect 42616 8304 42668 8356
rect 18236 8236 18288 8288
rect 19248 8279 19300 8288
rect 19248 8245 19257 8279
rect 19257 8245 19291 8279
rect 19291 8245 19300 8279
rect 19248 8236 19300 8245
rect 19708 8236 19760 8288
rect 27528 8236 27580 8288
rect 28632 8236 28684 8288
rect 29092 8236 29144 8288
rect 31208 8279 31260 8288
rect 31208 8245 31217 8279
rect 31217 8245 31251 8279
rect 31251 8245 31260 8279
rect 31208 8236 31260 8245
rect 33232 8236 33284 8288
rect 35808 8236 35860 8288
rect 36176 8236 36228 8288
rect 36268 8236 36320 8288
rect 37832 8236 37884 8288
rect 39120 8236 39172 8288
rect 40132 8236 40184 8288
rect 41696 8236 41748 8288
rect 44180 8236 44232 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 10600 8032 10652 8084
rect 16672 8032 16724 8084
rect 20720 8032 20772 8084
rect 11152 7964 11204 8016
rect 15752 7964 15804 8016
rect 10140 7828 10192 7880
rect 12992 7828 13044 7880
rect 17132 7896 17184 7948
rect 17224 7896 17276 7948
rect 18788 7964 18840 8016
rect 20536 7964 20588 8016
rect 21088 8032 21140 8084
rect 21824 8032 21876 8084
rect 22468 8032 22520 8084
rect 25596 8032 25648 8084
rect 25780 8032 25832 8084
rect 26056 8032 26108 8084
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 19708 7939 19760 7948
rect 17592 7896 17644 7905
rect 19708 7905 19717 7939
rect 19717 7905 19751 7939
rect 19751 7905 19760 7939
rect 19708 7896 19760 7905
rect 20260 7896 20312 7948
rect 20904 7896 20956 7948
rect 23756 7964 23808 8016
rect 32036 8032 32088 8084
rect 16672 7828 16724 7880
rect 17960 7828 18012 7880
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18604 7828 18656 7880
rect 18696 7828 18748 7880
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 9680 7760 9732 7812
rect 10508 7760 10560 7812
rect 17132 7692 17184 7744
rect 18788 7760 18840 7812
rect 18972 7828 19024 7880
rect 20812 7828 20864 7880
rect 21732 7896 21784 7948
rect 22100 7896 22152 7948
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 22560 7896 22612 7948
rect 25136 7939 25188 7948
rect 25136 7905 25145 7939
rect 25145 7905 25179 7939
rect 25179 7905 25188 7939
rect 25136 7896 25188 7905
rect 25228 7896 25280 7948
rect 25596 7896 25648 7948
rect 21456 7828 21508 7837
rect 19984 7760 20036 7812
rect 21272 7760 21324 7812
rect 22284 7760 22336 7812
rect 24676 7871 24728 7880
rect 24676 7837 24685 7871
rect 24685 7837 24719 7871
rect 24719 7837 24728 7871
rect 24676 7828 24728 7837
rect 30288 7964 30340 8016
rect 32956 8032 33008 8084
rect 33692 8032 33744 8084
rect 34336 8032 34388 8084
rect 35072 8032 35124 8084
rect 32772 7964 32824 8016
rect 28632 7896 28684 7948
rect 28816 7896 28868 7948
rect 21732 7692 21784 7744
rect 24216 7692 24268 7744
rect 24584 7760 24636 7812
rect 26976 7828 27028 7880
rect 29092 7896 29144 7948
rect 30104 7871 30156 7880
rect 30104 7837 30113 7871
rect 30113 7837 30147 7871
rect 30147 7837 30156 7871
rect 30288 7871 30340 7880
rect 30104 7828 30156 7837
rect 30288 7837 30297 7871
rect 30297 7837 30331 7871
rect 30331 7837 30340 7871
rect 30288 7828 30340 7837
rect 31024 7828 31076 7880
rect 25872 7760 25924 7812
rect 25136 7692 25188 7744
rect 25504 7692 25556 7744
rect 27252 7735 27304 7744
rect 27252 7701 27261 7735
rect 27261 7701 27295 7735
rect 27295 7701 27304 7735
rect 27252 7692 27304 7701
rect 32312 7896 32364 7948
rect 34244 7964 34296 8016
rect 35256 7964 35308 8016
rect 35348 7964 35400 8016
rect 33876 7871 33928 7880
rect 33048 7760 33100 7812
rect 27988 7692 28040 7744
rect 28908 7692 28960 7744
rect 29092 7735 29144 7744
rect 29092 7701 29101 7735
rect 29101 7701 29135 7735
rect 29135 7701 29144 7735
rect 29092 7692 29144 7701
rect 30104 7692 30156 7744
rect 30380 7692 30432 7744
rect 30840 7692 30892 7744
rect 32772 7692 32824 7744
rect 33876 7837 33885 7871
rect 33885 7837 33919 7871
rect 33919 7837 33928 7871
rect 33876 7828 33928 7837
rect 34428 7896 34480 7948
rect 34704 7828 34756 7880
rect 35072 7871 35124 7880
rect 35072 7837 35081 7871
rect 35081 7837 35115 7871
rect 35115 7837 35124 7871
rect 35072 7828 35124 7837
rect 36084 8032 36136 8084
rect 37004 8032 37056 8084
rect 37280 8032 37332 8084
rect 37556 8032 37608 8084
rect 38016 8032 38068 8084
rect 40776 8075 40828 8084
rect 40776 8041 40785 8075
rect 40785 8041 40819 8075
rect 40819 8041 40828 8075
rect 40776 8032 40828 8041
rect 41788 8032 41840 8084
rect 36912 7964 36964 8016
rect 36728 7896 36780 7948
rect 37372 7964 37424 8016
rect 37648 7964 37700 8016
rect 34152 7760 34204 7812
rect 34520 7692 34572 7744
rect 36176 7828 36228 7880
rect 39856 7896 39908 7948
rect 35348 7803 35400 7812
rect 35348 7769 35357 7803
rect 35357 7769 35391 7803
rect 35391 7769 35400 7803
rect 37740 7828 37792 7880
rect 38384 7828 38436 7880
rect 38476 7828 38528 7880
rect 38752 7871 38804 7880
rect 38752 7837 38761 7871
rect 38761 7837 38795 7871
rect 38795 7837 38804 7871
rect 38752 7828 38804 7837
rect 39120 7828 39172 7880
rect 39396 7828 39448 7880
rect 35348 7760 35400 7769
rect 37280 7760 37332 7812
rect 37372 7760 37424 7812
rect 39764 7760 39816 7812
rect 40132 7828 40184 7880
rect 41696 7828 41748 7880
rect 42248 7896 42300 7948
rect 42156 7871 42208 7880
rect 44916 8032 44968 8084
rect 58256 8075 58308 8084
rect 58256 8041 58265 8075
rect 58265 8041 58299 8075
rect 58299 8041 58308 8075
rect 58256 8032 58308 8041
rect 56876 7939 56928 7948
rect 42156 7837 42170 7871
rect 42170 7837 42204 7871
rect 42204 7837 42208 7871
rect 42156 7828 42208 7837
rect 42708 7828 42760 7880
rect 45468 7828 45520 7880
rect 49700 7828 49752 7880
rect 56876 7905 56885 7939
rect 56885 7905 56919 7939
rect 56919 7905 56928 7939
rect 56876 7896 56928 7905
rect 37004 7692 37056 7744
rect 37556 7692 37608 7744
rect 44272 7760 44324 7812
rect 56140 7803 56192 7812
rect 56140 7769 56149 7803
rect 56149 7769 56183 7803
rect 56183 7769 56192 7803
rect 56140 7760 56192 7769
rect 56600 7760 56652 7812
rect 44180 7735 44232 7744
rect 44180 7701 44189 7735
rect 44189 7701 44223 7735
rect 44223 7701 44232 7735
rect 44180 7692 44232 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 18696 7488 18748 7540
rect 19340 7488 19392 7540
rect 20904 7488 20956 7540
rect 21088 7488 21140 7540
rect 21548 7488 21600 7540
rect 22284 7488 22336 7540
rect 22744 7488 22796 7540
rect 23112 7488 23164 7540
rect 25872 7531 25924 7540
rect 25872 7497 25881 7531
rect 25881 7497 25915 7531
rect 25915 7497 25924 7531
rect 25872 7488 25924 7497
rect 26516 7488 26568 7540
rect 26700 7488 26752 7540
rect 31116 7531 31168 7540
rect 7012 7284 7064 7336
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 10324 7395 10376 7404
rect 9404 7352 9456 7361
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 27252 7420 27304 7472
rect 30104 7420 30156 7472
rect 31116 7497 31125 7531
rect 31125 7497 31159 7531
rect 31159 7497 31168 7531
rect 31116 7488 31168 7497
rect 32680 7531 32732 7540
rect 32680 7497 32689 7531
rect 32689 7497 32723 7531
rect 32723 7497 32732 7531
rect 32680 7488 32732 7497
rect 33784 7488 33836 7540
rect 35900 7488 35952 7540
rect 36084 7488 36136 7540
rect 36912 7488 36964 7540
rect 9680 7284 9732 7336
rect 10140 7327 10192 7336
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 17132 7327 17184 7336
rect 10600 7284 10652 7293
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 19340 7352 19392 7404
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 18052 7284 18104 7336
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 19800 7352 19852 7404
rect 20260 7352 20312 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 22008 7395 22060 7404
rect 20904 7352 20956 7361
rect 8852 7148 8904 7200
rect 18328 7216 18380 7268
rect 18604 7216 18656 7268
rect 19064 7216 19116 7268
rect 19892 7284 19944 7336
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 21364 7327 21416 7336
rect 21364 7293 21373 7327
rect 21373 7293 21407 7327
rect 21407 7293 21416 7327
rect 21364 7284 21416 7293
rect 21548 7284 21600 7336
rect 24584 7284 24636 7336
rect 15476 7148 15528 7200
rect 19524 7148 19576 7200
rect 20260 7216 20312 7268
rect 20720 7216 20772 7268
rect 21456 7216 21508 7268
rect 22192 7148 22244 7200
rect 24216 7148 24268 7200
rect 24952 7284 25004 7336
rect 25780 7284 25832 7336
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 33140 7420 33192 7472
rect 34704 7420 34756 7472
rect 35440 7463 35492 7472
rect 32036 7352 32088 7404
rect 34244 7352 34296 7404
rect 35440 7429 35449 7463
rect 35449 7429 35483 7463
rect 35483 7429 35492 7463
rect 35440 7420 35492 7429
rect 35256 7352 35308 7404
rect 28632 7284 28684 7336
rect 32588 7284 32640 7336
rect 34336 7327 34388 7336
rect 25228 7216 25280 7268
rect 27620 7216 27672 7268
rect 29276 7216 29328 7268
rect 31024 7216 31076 7268
rect 25044 7148 25096 7200
rect 28264 7148 28316 7200
rect 28816 7148 28868 7200
rect 29552 7148 29604 7200
rect 30748 7148 30800 7200
rect 31208 7148 31260 7200
rect 31484 7148 31536 7200
rect 31760 7148 31812 7200
rect 32680 7216 32732 7268
rect 33140 7216 33192 7268
rect 33600 7216 33652 7268
rect 34336 7293 34345 7327
rect 34345 7293 34379 7327
rect 34379 7293 34388 7327
rect 34336 7284 34388 7293
rect 34428 7327 34480 7336
rect 34428 7293 34437 7327
rect 34437 7293 34471 7327
rect 34471 7293 34480 7327
rect 35808 7352 35860 7404
rect 37004 7420 37056 7472
rect 37280 7352 37332 7404
rect 37464 7395 37516 7404
rect 37464 7361 37473 7395
rect 37473 7361 37507 7395
rect 37507 7361 37516 7395
rect 37464 7352 37516 7361
rect 37740 7352 37792 7404
rect 34428 7284 34480 7293
rect 35992 7284 36044 7336
rect 37188 7284 37240 7336
rect 37832 7327 37884 7336
rect 37832 7293 37841 7327
rect 37841 7293 37875 7327
rect 37875 7293 37884 7327
rect 37832 7284 37884 7293
rect 36084 7216 36136 7268
rect 36268 7259 36320 7268
rect 36268 7225 36277 7259
rect 36277 7225 36311 7259
rect 36311 7225 36320 7259
rect 36268 7216 36320 7225
rect 37004 7216 37056 7268
rect 38200 7352 38252 7404
rect 42616 7488 42668 7540
rect 43628 7488 43680 7540
rect 39120 7420 39172 7472
rect 42156 7420 42208 7472
rect 55220 7488 55272 7540
rect 55404 7488 55456 7540
rect 57244 7488 57296 7540
rect 43904 7420 43956 7472
rect 44180 7420 44232 7472
rect 38292 7284 38344 7336
rect 40132 7352 40184 7404
rect 41604 7395 41656 7404
rect 41604 7361 41613 7395
rect 41613 7361 41647 7395
rect 41647 7361 41656 7395
rect 41604 7352 41656 7361
rect 41788 7395 41840 7404
rect 41788 7361 41797 7395
rect 41797 7361 41831 7395
rect 41831 7361 41840 7395
rect 41788 7352 41840 7361
rect 38384 7216 38436 7268
rect 40408 7216 40460 7268
rect 42064 7216 42116 7268
rect 42708 7352 42760 7404
rect 42892 7352 42944 7404
rect 51080 7420 51132 7472
rect 56140 7420 56192 7472
rect 44824 7395 44876 7404
rect 44824 7361 44833 7395
rect 44833 7361 44867 7395
rect 44867 7361 44876 7395
rect 44824 7352 44876 7361
rect 43260 7284 43312 7336
rect 42800 7216 42852 7268
rect 53932 7284 53984 7336
rect 57336 7327 57388 7336
rect 57336 7293 57345 7327
rect 57345 7293 57379 7327
rect 57379 7293 57388 7327
rect 57336 7284 57388 7293
rect 58256 7395 58308 7404
rect 58256 7361 58265 7395
rect 58265 7361 58299 7395
rect 58299 7361 58308 7395
rect 58256 7352 58308 7361
rect 39212 7148 39264 7200
rect 42892 7148 42944 7200
rect 44824 7148 44876 7200
rect 56784 7148 56836 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10508 6944 10560 6996
rect 17592 6987 17644 6996
rect 17592 6953 17601 6987
rect 17601 6953 17635 6987
rect 17635 6953 17644 6987
rect 17592 6944 17644 6953
rect 14556 6876 14608 6928
rect 19294 6944 19346 6996
rect 19432 6944 19484 6996
rect 19524 6944 19576 6996
rect 22928 6944 22980 6996
rect 17224 6808 17276 6860
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11336 6740 11388 6792
rect 11704 6740 11756 6792
rect 16396 6740 16448 6792
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 18052 6808 18104 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 22100 6876 22152 6928
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 18696 6808 18748 6860
rect 22836 6808 22888 6860
rect 24216 6944 24268 6996
rect 25228 6944 25280 6996
rect 23756 6876 23808 6928
rect 24952 6876 25004 6928
rect 18144 6740 18196 6792
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20076 6740 20128 6792
rect 10508 6672 10560 6724
rect 13452 6672 13504 6724
rect 18972 6672 19024 6724
rect 19616 6672 19668 6724
rect 20260 6740 20312 6792
rect 20628 6740 20680 6792
rect 21088 6740 21140 6792
rect 22192 6740 22244 6792
rect 22304 6783 22356 6792
rect 22304 6749 22327 6783
rect 22327 6749 22356 6783
rect 22304 6740 22356 6749
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 21272 6672 21324 6724
rect 23112 6740 23164 6792
rect 23756 6740 23808 6792
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 24124 6740 24176 6792
rect 23388 6672 23440 6724
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 25596 6851 25648 6860
rect 25596 6817 25605 6851
rect 25605 6817 25639 6851
rect 25639 6817 25648 6851
rect 25596 6808 25648 6817
rect 24860 6740 24912 6749
rect 27068 6740 27120 6792
rect 29552 6944 29604 6996
rect 30288 6944 30340 6996
rect 29460 6808 29512 6860
rect 30196 6808 30248 6860
rect 30472 6851 30524 6860
rect 30472 6817 30481 6851
rect 30481 6817 30515 6851
rect 30515 6817 30524 6851
rect 33140 6876 33192 6928
rect 30472 6808 30524 6817
rect 27528 6740 27580 6792
rect 29276 6740 29328 6792
rect 32772 6808 32824 6860
rect 33324 6944 33376 6996
rect 34152 6944 34204 6996
rect 35256 6944 35308 6996
rect 35716 6944 35768 6996
rect 33600 6876 33652 6928
rect 34888 6876 34940 6928
rect 35992 6944 36044 6996
rect 36084 6944 36136 6996
rect 31116 6783 31168 6792
rect 14832 6604 14884 6656
rect 17500 6604 17552 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 20352 6604 20404 6656
rect 23020 6604 23072 6656
rect 25688 6672 25740 6724
rect 26056 6672 26108 6724
rect 27988 6672 28040 6724
rect 23756 6604 23808 6656
rect 26976 6647 27028 6656
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 26976 6604 27028 6613
rect 27344 6604 27396 6656
rect 27528 6604 27580 6656
rect 27896 6604 27948 6656
rect 28724 6672 28776 6724
rect 28816 6647 28868 6656
rect 28816 6613 28825 6647
rect 28825 6613 28859 6647
rect 28859 6613 28868 6647
rect 28816 6604 28868 6613
rect 31116 6749 31125 6783
rect 31125 6749 31159 6783
rect 31159 6749 31168 6783
rect 31116 6740 31168 6749
rect 31208 6740 31260 6792
rect 31024 6672 31076 6724
rect 31576 6672 31628 6724
rect 32680 6783 32732 6792
rect 32680 6749 32689 6783
rect 32689 6749 32723 6783
rect 32723 6749 32732 6783
rect 32680 6740 32732 6749
rect 33140 6740 33192 6792
rect 33692 6808 33744 6860
rect 34244 6808 34296 6860
rect 33784 6783 33836 6792
rect 33048 6672 33100 6724
rect 33784 6749 33793 6783
rect 33793 6749 33827 6783
rect 33827 6749 33836 6783
rect 33784 6740 33836 6749
rect 33968 6740 34020 6792
rect 30380 6604 30432 6656
rect 31484 6604 31536 6656
rect 31668 6647 31720 6656
rect 31668 6613 31677 6647
rect 31677 6613 31711 6647
rect 31711 6613 31720 6647
rect 31668 6604 31720 6613
rect 32220 6604 32272 6656
rect 33232 6604 33284 6656
rect 33692 6715 33744 6724
rect 33692 6681 33701 6715
rect 33701 6681 33735 6715
rect 33735 6681 33744 6715
rect 34796 6808 34848 6860
rect 33692 6672 33744 6681
rect 34612 6672 34664 6724
rect 36912 6876 36964 6928
rect 37832 6876 37884 6928
rect 38384 6944 38436 6996
rect 42800 6987 42852 6996
rect 42800 6953 42809 6987
rect 42809 6953 42843 6987
rect 42843 6953 42852 6987
rect 42800 6944 42852 6953
rect 58256 6987 58308 6996
rect 58256 6953 58265 6987
rect 58265 6953 58299 6987
rect 58299 6953 58308 6987
rect 58256 6944 58308 6953
rect 35624 6808 35676 6860
rect 35348 6783 35400 6792
rect 35348 6749 35375 6783
rect 35375 6749 35400 6783
rect 35348 6740 35400 6749
rect 35716 6740 35768 6792
rect 36084 6740 36136 6792
rect 36360 6740 36412 6792
rect 37004 6740 37056 6792
rect 37648 6808 37700 6860
rect 38292 6808 38344 6860
rect 41604 6876 41656 6928
rect 42064 6851 42116 6860
rect 35992 6672 36044 6724
rect 36084 6604 36136 6656
rect 36268 6604 36320 6656
rect 36544 6604 36596 6656
rect 37004 6647 37056 6656
rect 37004 6613 37013 6647
rect 37013 6613 37047 6647
rect 37047 6613 37056 6647
rect 37004 6604 37056 6613
rect 37832 6672 37884 6724
rect 38476 6740 38528 6792
rect 40040 6783 40092 6792
rect 40040 6749 40049 6783
rect 40049 6749 40083 6783
rect 40083 6749 40092 6783
rect 40040 6740 40092 6749
rect 38200 6672 38252 6724
rect 40592 6740 40644 6792
rect 40868 6740 40920 6792
rect 37924 6604 37976 6656
rect 41696 6672 41748 6724
rect 42064 6817 42073 6851
rect 42073 6817 42107 6851
rect 42107 6817 42116 6851
rect 42064 6808 42116 6817
rect 47676 6876 47728 6928
rect 56876 6851 56928 6860
rect 56876 6817 56885 6851
rect 56885 6817 56919 6851
rect 56919 6817 56928 6851
rect 56876 6808 56928 6817
rect 43260 6783 43312 6792
rect 43260 6749 43269 6783
rect 43269 6749 43303 6783
rect 43303 6749 43312 6783
rect 43260 6740 43312 6749
rect 43444 6740 43496 6792
rect 43812 6783 43864 6792
rect 43812 6749 43821 6783
rect 43821 6749 43855 6783
rect 43855 6749 43864 6783
rect 43812 6740 43864 6749
rect 56784 6740 56836 6792
rect 45284 6672 45336 6724
rect 56048 6672 56100 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 10600 6400 10652 6452
rect 15292 6400 15344 6452
rect 18052 6400 18104 6452
rect 19340 6400 19392 6452
rect 19984 6400 20036 6452
rect 21088 6400 21140 6452
rect 22652 6400 22704 6452
rect 22836 6400 22888 6452
rect 23296 6400 23348 6452
rect 26792 6400 26844 6452
rect 27988 6443 28040 6452
rect 27988 6409 27997 6443
rect 27997 6409 28031 6443
rect 28031 6409 28040 6443
rect 27988 6400 28040 6409
rect 29460 6400 29512 6452
rect 9680 6375 9732 6384
rect 9680 6341 9689 6375
rect 9689 6341 9723 6375
rect 9723 6341 9732 6375
rect 9680 6332 9732 6341
rect 9588 6264 9640 6316
rect 11612 6264 11664 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 8944 6196 8996 6248
rect 20536 6332 20588 6384
rect 21732 6332 21784 6384
rect 22100 6332 22152 6384
rect 28816 6332 28868 6384
rect 29184 6332 29236 6384
rect 15844 6264 15896 6316
rect 18696 6264 18748 6316
rect 19248 6264 19300 6316
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 20076 6264 20128 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 21272 6264 21324 6316
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 18972 6196 19024 6248
rect 19892 6196 19944 6248
rect 21732 6196 21784 6248
rect 21916 6196 21968 6248
rect 22468 6264 22520 6316
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 23296 6264 23348 6316
rect 24952 6307 25004 6316
rect 24952 6273 24961 6307
rect 24961 6273 24995 6307
rect 24995 6273 25004 6307
rect 24952 6264 25004 6273
rect 24216 6196 24268 6248
rect 27160 6239 27212 6248
rect 5080 6128 5132 6180
rect 11060 6171 11112 6180
rect 11060 6137 11069 6171
rect 11069 6137 11103 6171
rect 11103 6137 11112 6171
rect 11060 6128 11112 6137
rect 17132 6171 17184 6180
rect 17132 6137 17141 6171
rect 17141 6137 17175 6171
rect 17175 6137 17184 6171
rect 17132 6128 17184 6137
rect 17776 6128 17828 6180
rect 10324 6060 10376 6112
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 21916 6060 21968 6112
rect 22192 6128 22244 6180
rect 25044 6128 25096 6180
rect 25504 6128 25556 6180
rect 27160 6205 27169 6239
rect 27169 6205 27203 6239
rect 27203 6205 27212 6239
rect 27160 6196 27212 6205
rect 27528 6264 27580 6316
rect 29368 6264 29420 6316
rect 36176 6400 36228 6452
rect 36544 6400 36596 6452
rect 29736 6307 29788 6316
rect 28632 6239 28684 6248
rect 28632 6205 28641 6239
rect 28641 6205 28675 6239
rect 28675 6205 28684 6239
rect 28632 6196 28684 6205
rect 29736 6273 29745 6307
rect 29745 6273 29779 6307
rect 29779 6273 29788 6307
rect 29736 6264 29788 6273
rect 31668 6332 31720 6384
rect 32496 6332 32548 6384
rect 34244 6375 34296 6384
rect 30288 6307 30340 6316
rect 30288 6273 30297 6307
rect 30297 6273 30331 6307
rect 30331 6273 30340 6307
rect 30288 6264 30340 6273
rect 29920 6196 29972 6248
rect 26608 6128 26660 6180
rect 32312 6307 32364 6316
rect 32312 6273 32321 6307
rect 32321 6273 32355 6307
rect 32355 6273 32364 6307
rect 32312 6264 32364 6273
rect 34244 6341 34253 6375
rect 34253 6341 34287 6375
rect 34287 6341 34296 6375
rect 34244 6332 34296 6341
rect 34796 6332 34848 6384
rect 35256 6375 35308 6384
rect 35256 6341 35265 6375
rect 35265 6341 35299 6375
rect 35299 6341 35308 6375
rect 35256 6332 35308 6341
rect 36268 6332 36320 6384
rect 34520 6307 34572 6316
rect 34520 6273 34529 6307
rect 34529 6273 34563 6307
rect 34563 6273 34572 6307
rect 34520 6264 34572 6273
rect 22284 6060 22336 6112
rect 23756 6060 23808 6112
rect 29000 6060 29052 6112
rect 29184 6060 29236 6112
rect 31116 6060 31168 6112
rect 31484 6103 31536 6112
rect 31484 6069 31493 6103
rect 31493 6069 31527 6103
rect 31527 6069 31536 6103
rect 31484 6060 31536 6069
rect 31852 6060 31904 6112
rect 34152 6196 34204 6248
rect 33600 6128 33652 6180
rect 34060 6128 34112 6180
rect 34612 6196 34664 6248
rect 35164 6264 35216 6316
rect 35532 6264 35584 6316
rect 35808 6264 35860 6316
rect 36360 6307 36412 6316
rect 36360 6273 36369 6307
rect 36369 6273 36403 6307
rect 36403 6273 36412 6307
rect 36360 6264 36412 6273
rect 37004 6264 37056 6316
rect 37096 6264 37148 6316
rect 38200 6400 38252 6452
rect 38292 6332 38344 6384
rect 39028 6400 39080 6452
rect 40040 6400 40092 6452
rect 43260 6400 43312 6452
rect 35624 6196 35676 6248
rect 34428 6128 34480 6180
rect 37188 6196 37240 6248
rect 41788 6264 41840 6316
rect 45100 6332 45152 6384
rect 56140 6400 56192 6452
rect 57244 6332 57296 6384
rect 56048 6307 56100 6316
rect 56048 6273 56057 6307
rect 56057 6273 56091 6307
rect 56091 6273 56100 6307
rect 56048 6264 56100 6273
rect 56692 6264 56744 6316
rect 58072 6307 58124 6316
rect 58072 6273 58081 6307
rect 58081 6273 58115 6307
rect 58115 6273 58124 6307
rect 58072 6264 58124 6273
rect 35992 6128 36044 6180
rect 34704 6060 34756 6112
rect 36176 6060 36228 6112
rect 41696 6128 41748 6180
rect 45008 6196 45060 6248
rect 56140 6196 56192 6248
rect 48596 6128 48648 6180
rect 55220 6128 55272 6180
rect 38476 6060 38528 6112
rect 55772 6103 55824 6112
rect 55772 6069 55781 6103
rect 55781 6069 55815 6103
rect 55815 6069 55824 6103
rect 55772 6060 55824 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 10968 5856 11020 5908
rect 16488 5856 16540 5908
rect 18972 5856 19024 5908
rect 20260 5856 20312 5908
rect 20996 5856 21048 5908
rect 23572 5856 23624 5908
rect 5540 5788 5592 5840
rect 17132 5788 17184 5840
rect 16120 5720 16172 5772
rect 9220 5652 9272 5704
rect 17316 5720 17368 5772
rect 18696 5720 18748 5772
rect 19340 5720 19392 5772
rect 19892 5763 19944 5772
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 23204 5788 23256 5840
rect 23848 5788 23900 5840
rect 16488 5652 16540 5704
rect 16856 5652 16908 5704
rect 17592 5652 17644 5704
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 18788 5652 18840 5704
rect 20260 5652 20312 5704
rect 21088 5720 21140 5772
rect 22836 5763 22888 5772
rect 22836 5729 22845 5763
rect 22845 5729 22879 5763
rect 22879 5729 22888 5763
rect 22836 5720 22888 5729
rect 25136 5720 25188 5772
rect 25596 5856 25648 5908
rect 27068 5856 27120 5908
rect 26608 5831 26660 5840
rect 26608 5797 26617 5831
rect 26617 5797 26651 5831
rect 26651 5797 26660 5831
rect 26608 5788 26660 5797
rect 27344 5856 27396 5908
rect 21824 5695 21876 5704
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 10508 5584 10560 5636
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 12256 5584 12308 5636
rect 12532 5627 12584 5636
rect 12532 5593 12541 5627
rect 12541 5593 12575 5627
rect 12575 5593 12584 5627
rect 12532 5584 12584 5593
rect 13084 5584 13136 5636
rect 14648 5584 14700 5636
rect 17776 5627 17828 5636
rect 17776 5593 17785 5627
rect 17785 5593 17819 5627
rect 17819 5593 17828 5627
rect 17776 5584 17828 5593
rect 12624 5516 12676 5568
rect 19984 5584 20036 5636
rect 20260 5516 20312 5568
rect 21272 5584 21324 5636
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 24308 5652 24360 5704
rect 24400 5652 24452 5704
rect 24676 5652 24728 5704
rect 29368 5788 29420 5840
rect 31484 5788 31536 5840
rect 28448 5720 28500 5772
rect 29000 5695 29052 5704
rect 23480 5584 23532 5636
rect 24860 5584 24912 5636
rect 25596 5584 25648 5636
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 29184 5695 29236 5704
rect 29184 5661 29193 5695
rect 29193 5661 29227 5695
rect 29227 5661 29236 5695
rect 29184 5652 29236 5661
rect 29736 5720 29788 5772
rect 30472 5720 30524 5772
rect 33232 5788 33284 5840
rect 33324 5788 33376 5840
rect 34980 5788 35032 5840
rect 35624 5788 35676 5840
rect 35532 5720 35584 5772
rect 35900 5720 35952 5772
rect 27712 5584 27764 5636
rect 27804 5584 27856 5636
rect 28080 5584 28132 5636
rect 31024 5652 31076 5704
rect 33416 5652 33468 5704
rect 34980 5652 35032 5704
rect 37648 5856 37700 5908
rect 37832 5856 37884 5908
rect 38752 5856 38804 5908
rect 39120 5856 39172 5908
rect 41696 5899 41748 5908
rect 41696 5865 41705 5899
rect 41705 5865 41739 5899
rect 41739 5865 41748 5899
rect 41696 5856 41748 5865
rect 43720 5856 43772 5908
rect 45284 5899 45336 5908
rect 45284 5865 45293 5899
rect 45293 5865 45327 5899
rect 45327 5865 45336 5899
rect 45284 5856 45336 5865
rect 31668 5584 31720 5636
rect 31852 5584 31904 5636
rect 34520 5584 34572 5636
rect 36268 5652 36320 5704
rect 53932 5788 53984 5840
rect 37096 5720 37148 5772
rect 37372 5720 37424 5772
rect 38384 5763 38436 5772
rect 38384 5729 38393 5763
rect 38393 5729 38427 5763
rect 38427 5729 38436 5763
rect 38384 5720 38436 5729
rect 40408 5652 40460 5704
rect 40868 5652 40920 5704
rect 20904 5516 20956 5568
rect 22100 5516 22152 5568
rect 26148 5516 26200 5568
rect 28172 5516 28224 5568
rect 28724 5516 28776 5568
rect 30656 5559 30708 5568
rect 30656 5525 30665 5559
rect 30665 5525 30699 5559
rect 30699 5525 30708 5559
rect 30656 5516 30708 5525
rect 31484 5516 31536 5568
rect 32220 5516 32272 5568
rect 32404 5559 32456 5568
rect 32404 5525 32413 5559
rect 32413 5525 32447 5559
rect 32447 5525 32456 5559
rect 32404 5516 32456 5525
rect 32588 5516 32640 5568
rect 33416 5516 33468 5568
rect 34612 5516 34664 5568
rect 37188 5559 37240 5568
rect 37188 5525 37197 5559
rect 37197 5525 37231 5559
rect 37231 5525 37240 5559
rect 37188 5516 37240 5525
rect 37832 5516 37884 5568
rect 38476 5584 38528 5636
rect 38936 5584 38988 5636
rect 41604 5627 41656 5636
rect 41604 5593 41613 5627
rect 41613 5593 41647 5627
rect 41647 5593 41656 5627
rect 41604 5584 41656 5593
rect 38200 5516 38252 5568
rect 42800 5652 42852 5704
rect 42892 5652 42944 5704
rect 43720 5720 43772 5772
rect 56876 5763 56928 5772
rect 56876 5729 56885 5763
rect 56885 5729 56919 5763
rect 56919 5729 56928 5763
rect 56876 5720 56928 5729
rect 43720 5627 43772 5636
rect 43720 5593 43729 5627
rect 43729 5593 43763 5627
rect 43763 5593 43772 5627
rect 43720 5584 43772 5593
rect 44364 5584 44416 5636
rect 55772 5652 55824 5704
rect 58348 5584 58400 5636
rect 43444 5516 43496 5568
rect 43812 5559 43864 5568
rect 43812 5525 43821 5559
rect 43821 5525 43855 5559
rect 43855 5525 43864 5559
rect 43812 5516 43864 5525
rect 57336 5516 57388 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 9588 5355 9640 5364
rect 9588 5321 9597 5355
rect 9597 5321 9631 5355
rect 9631 5321 9640 5355
rect 9588 5312 9640 5321
rect 8392 5176 8444 5228
rect 8576 5176 8628 5228
rect 9036 5176 9088 5228
rect 9864 5312 9916 5364
rect 23756 5312 23808 5364
rect 24860 5312 24912 5364
rect 27712 5355 27764 5364
rect 27712 5321 27721 5355
rect 27721 5321 27755 5355
rect 27755 5321 27764 5355
rect 27712 5312 27764 5321
rect 28080 5355 28132 5364
rect 28080 5321 28089 5355
rect 28089 5321 28123 5355
rect 28123 5321 28132 5355
rect 28080 5312 28132 5321
rect 31484 5312 31536 5364
rect 10600 5244 10652 5296
rect 11244 5244 11296 5296
rect 11980 5244 12032 5296
rect 15844 5287 15896 5296
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 7564 5040 7616 5092
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 10784 5176 10836 5228
rect 11796 5176 11848 5228
rect 10324 5108 10376 5160
rect 11336 5108 11388 5160
rect 13820 5176 13872 5228
rect 15844 5253 15853 5287
rect 15853 5253 15887 5287
rect 15887 5253 15896 5287
rect 15844 5244 15896 5253
rect 19340 5244 19392 5296
rect 24032 5244 24084 5296
rect 24952 5244 25004 5296
rect 28724 5244 28776 5296
rect 14096 5176 14148 5228
rect 16948 5219 17000 5228
rect 8484 4972 8536 5024
rect 10048 5040 10100 5092
rect 11428 5040 11480 5092
rect 12164 4972 12216 5024
rect 13360 4972 13412 5024
rect 16120 5083 16172 5092
rect 16120 5049 16129 5083
rect 16129 5049 16163 5083
rect 16163 5049 16172 5083
rect 16120 5040 16172 5049
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 19248 5176 19300 5228
rect 19432 5219 19484 5228
rect 19432 5185 19441 5219
rect 19441 5185 19475 5219
rect 19475 5185 19484 5219
rect 19432 5176 19484 5185
rect 19984 5176 20036 5228
rect 20628 5176 20680 5228
rect 21824 5176 21876 5228
rect 22468 5176 22520 5228
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 16764 5108 16816 5160
rect 18972 5151 19024 5160
rect 18972 5117 18981 5151
rect 18981 5117 19015 5151
rect 19015 5117 19024 5151
rect 18972 5108 19024 5117
rect 19064 5108 19116 5160
rect 20812 5108 20864 5160
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 19156 5040 19208 5092
rect 19248 5040 19300 5092
rect 20260 5040 20312 5092
rect 24492 5176 24544 5228
rect 25136 5219 25188 5228
rect 25136 5185 25145 5219
rect 25145 5185 25179 5219
rect 25179 5185 25188 5219
rect 25136 5176 25188 5185
rect 28264 5176 28316 5228
rect 28908 5219 28960 5228
rect 28908 5185 28917 5219
rect 28917 5185 28951 5219
rect 28951 5185 28960 5219
rect 28908 5176 28960 5185
rect 29184 5176 29236 5228
rect 29552 5219 29604 5228
rect 29552 5185 29561 5219
rect 29561 5185 29595 5219
rect 29595 5185 29604 5219
rect 29552 5176 29604 5185
rect 29828 5219 29880 5228
rect 29828 5185 29862 5219
rect 29862 5185 29880 5219
rect 30196 5244 30248 5296
rect 31024 5244 31076 5296
rect 35348 5312 35400 5364
rect 36084 5312 36136 5364
rect 36452 5312 36504 5364
rect 38476 5312 38528 5364
rect 38568 5312 38620 5364
rect 40776 5312 40828 5364
rect 43352 5312 43404 5364
rect 43536 5355 43588 5364
rect 43536 5321 43545 5355
rect 43545 5321 43579 5355
rect 43579 5321 43588 5355
rect 43536 5312 43588 5321
rect 45008 5355 45060 5364
rect 45008 5321 45017 5355
rect 45017 5321 45051 5355
rect 45051 5321 45060 5355
rect 45008 5312 45060 5321
rect 45376 5312 45428 5364
rect 57244 5355 57296 5364
rect 57244 5321 57253 5355
rect 57253 5321 57287 5355
rect 57287 5321 57296 5355
rect 57244 5312 57296 5321
rect 29828 5176 29880 5185
rect 31760 5176 31812 5228
rect 31852 5176 31904 5228
rect 24400 5151 24452 5160
rect 24400 5117 24409 5151
rect 24409 5117 24443 5151
rect 24443 5117 24452 5151
rect 24400 5108 24452 5117
rect 24676 5108 24728 5160
rect 28172 5151 28224 5160
rect 28172 5117 28181 5151
rect 28181 5117 28215 5151
rect 28215 5117 28224 5151
rect 28172 5108 28224 5117
rect 27896 5040 27948 5092
rect 28632 5108 28684 5160
rect 29460 5108 29512 5160
rect 31392 5151 31444 5160
rect 31392 5117 31401 5151
rect 31401 5117 31435 5151
rect 31435 5117 31444 5151
rect 31392 5108 31444 5117
rect 31944 5108 31996 5160
rect 33784 5176 33836 5228
rect 34244 5176 34296 5228
rect 38660 5244 38712 5296
rect 35072 5219 35124 5228
rect 35072 5185 35081 5219
rect 35081 5185 35115 5219
rect 35115 5185 35124 5219
rect 35072 5176 35124 5185
rect 30564 5040 30616 5092
rect 31116 5040 31168 5092
rect 31484 5040 31536 5092
rect 32036 5040 32088 5092
rect 34060 5108 34112 5160
rect 35808 5176 35860 5228
rect 36176 5219 36228 5228
rect 36176 5185 36185 5219
rect 36185 5185 36219 5219
rect 36219 5185 36228 5219
rect 36176 5176 36228 5185
rect 38292 5219 38344 5228
rect 38292 5185 38301 5219
rect 38301 5185 38335 5219
rect 38335 5185 38344 5219
rect 38292 5176 38344 5185
rect 38568 5176 38620 5228
rect 40316 5244 40368 5296
rect 41512 5244 41564 5296
rect 39580 5176 39632 5228
rect 40500 5219 40552 5228
rect 40500 5185 40509 5219
rect 40509 5185 40543 5219
rect 40543 5185 40552 5219
rect 40500 5176 40552 5185
rect 41696 5176 41748 5228
rect 35348 5151 35400 5160
rect 35348 5117 35357 5151
rect 35357 5117 35391 5151
rect 35391 5117 35400 5151
rect 35348 5108 35400 5117
rect 35900 5108 35952 5160
rect 37372 5108 37424 5160
rect 40132 5108 40184 5160
rect 43536 5176 43588 5228
rect 44824 5219 44876 5228
rect 44824 5185 44833 5219
rect 44833 5185 44867 5219
rect 44867 5185 44876 5219
rect 44824 5176 44876 5185
rect 45284 5176 45336 5228
rect 45652 5219 45704 5228
rect 45652 5185 45661 5219
rect 45661 5185 45695 5219
rect 45695 5185 45704 5219
rect 45652 5176 45704 5185
rect 45744 5176 45796 5228
rect 53196 5176 53248 5228
rect 57152 5219 57204 5228
rect 57152 5185 57161 5219
rect 57161 5185 57195 5219
rect 57195 5185 57204 5219
rect 57152 5176 57204 5185
rect 57336 5219 57388 5228
rect 57336 5185 57345 5219
rect 57345 5185 57379 5219
rect 57379 5185 57388 5219
rect 57336 5176 57388 5185
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 44916 5108 44968 5160
rect 45008 5108 45060 5160
rect 33508 5083 33560 5092
rect 33508 5049 33517 5083
rect 33517 5049 33551 5083
rect 33551 5049 33560 5083
rect 33508 5040 33560 5049
rect 35072 5040 35124 5092
rect 38752 5040 38804 5092
rect 39396 5040 39448 5092
rect 19064 4972 19116 5024
rect 21364 4972 21416 5024
rect 24032 4972 24084 5024
rect 25872 4972 25924 5024
rect 27528 4972 27580 5024
rect 30196 4972 30248 5024
rect 30288 4972 30340 5024
rect 32404 5015 32456 5024
rect 32404 4981 32413 5015
rect 32413 4981 32447 5015
rect 32447 4981 32456 5015
rect 32404 4972 32456 4981
rect 32680 5015 32732 5024
rect 32680 4981 32689 5015
rect 32689 4981 32723 5015
rect 32723 4981 32732 5015
rect 32680 4972 32732 4981
rect 34428 4972 34480 5024
rect 34796 4972 34848 5024
rect 36544 4972 36596 5024
rect 36636 4972 36688 5024
rect 38476 4972 38528 5024
rect 39212 4972 39264 5024
rect 40592 4972 40644 5024
rect 42708 4972 42760 5024
rect 43996 4972 44048 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 9404 4768 9456 4820
rect 9588 4768 9640 4820
rect 7012 4743 7064 4752
rect 7012 4709 7021 4743
rect 7021 4709 7055 4743
rect 7055 4709 7064 4743
rect 7012 4700 7064 4709
rect 8668 4700 8720 4752
rect 10140 4768 10192 4820
rect 12348 4768 12400 4820
rect 11704 4743 11756 4752
rect 11704 4709 11713 4743
rect 11713 4709 11747 4743
rect 11747 4709 11756 4743
rect 11704 4700 11756 4709
rect 12072 4700 12124 4752
rect 12532 4743 12584 4752
rect 12532 4709 12541 4743
rect 12541 4709 12575 4743
rect 12575 4709 12584 4743
rect 12532 4700 12584 4709
rect 12900 4700 12952 4752
rect 19432 4768 19484 4820
rect 28080 4768 28132 4820
rect 29828 4811 29880 4820
rect 29828 4777 29837 4811
rect 29837 4777 29871 4811
rect 29871 4777 29880 4811
rect 29828 4768 29880 4777
rect 30656 4768 30708 4820
rect 33784 4768 33836 4820
rect 37096 4768 37148 4820
rect 37924 4768 37976 4820
rect 40224 4768 40276 4820
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 9772 4632 9824 4684
rect 10324 4632 10376 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 12164 4632 12216 4684
rect 9680 4607 9732 4616
rect 6644 4496 6696 4548
rect 8024 4496 8076 4548
rect 8668 4496 8720 4548
rect 9312 4496 9364 4548
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 19064 4632 19116 4684
rect 20996 4700 21048 4752
rect 22008 4700 22060 4752
rect 21088 4632 21140 4684
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 21456 4632 21508 4684
rect 23480 4700 23532 4752
rect 28632 4700 28684 4752
rect 36084 4700 36136 4752
rect 39304 4700 39356 4752
rect 40592 4700 40644 4752
rect 44272 4768 44324 4820
rect 45744 4768 45796 4820
rect 41512 4700 41564 4752
rect 44916 4700 44968 4752
rect 48228 4768 48280 4820
rect 54208 4811 54260 4820
rect 54208 4777 54217 4811
rect 54217 4777 54251 4811
rect 54251 4777 54260 4811
rect 54208 4768 54260 4777
rect 56692 4768 56744 4820
rect 12164 4496 12216 4548
rect 13544 4496 13596 4548
rect 15844 4496 15896 4548
rect 16764 4496 16816 4548
rect 17224 4496 17276 4548
rect 9128 4428 9180 4480
rect 9496 4428 9548 4480
rect 12348 4428 12400 4480
rect 18512 4564 18564 4616
rect 19616 4564 19668 4616
rect 20720 4564 20772 4616
rect 20812 4564 20864 4616
rect 22560 4632 22612 4684
rect 23756 4632 23808 4684
rect 23940 4675 23992 4684
rect 23940 4641 23949 4675
rect 23949 4641 23983 4675
rect 23983 4641 23992 4675
rect 23940 4632 23992 4641
rect 24860 4632 24912 4684
rect 25136 4675 25188 4684
rect 25136 4641 25145 4675
rect 25145 4641 25179 4675
rect 25179 4641 25188 4675
rect 25136 4632 25188 4641
rect 22100 4564 22152 4616
rect 22192 4564 22244 4616
rect 24768 4564 24820 4616
rect 27528 4675 27580 4684
rect 27528 4641 27537 4675
rect 27537 4641 27571 4675
rect 27571 4641 27580 4675
rect 27528 4632 27580 4641
rect 28954 4632 29006 4684
rect 30288 4675 30340 4684
rect 30288 4641 30297 4675
rect 30297 4641 30331 4675
rect 30331 4641 30340 4675
rect 30288 4632 30340 4641
rect 30472 4675 30524 4684
rect 30472 4641 30481 4675
rect 30481 4641 30515 4675
rect 30515 4641 30524 4675
rect 30472 4632 30524 4641
rect 27988 4564 28040 4616
rect 28356 4564 28408 4616
rect 20628 4496 20680 4548
rect 24492 4496 24544 4548
rect 24584 4496 24636 4548
rect 22652 4428 22704 4480
rect 23572 4428 23624 4480
rect 27804 4496 27856 4548
rect 29184 4564 29236 4616
rect 30104 4564 30156 4616
rect 32312 4564 32364 4616
rect 30840 4496 30892 4548
rect 34612 4632 34664 4684
rect 35532 4675 35584 4684
rect 35532 4641 35541 4675
rect 35541 4641 35575 4675
rect 35575 4641 35584 4675
rect 35532 4632 35584 4641
rect 33600 4607 33652 4616
rect 33600 4573 33609 4607
rect 33609 4573 33643 4607
rect 33643 4573 33652 4607
rect 33600 4564 33652 4573
rect 38292 4632 38344 4684
rect 36176 4607 36228 4616
rect 32956 4539 33008 4548
rect 32956 4505 32965 4539
rect 32965 4505 32999 4539
rect 32999 4505 33008 4539
rect 32956 4496 33008 4505
rect 33140 4539 33192 4548
rect 33140 4505 33149 4539
rect 33149 4505 33183 4539
rect 33183 4505 33192 4539
rect 33140 4496 33192 4505
rect 26976 4471 27028 4480
rect 26976 4437 26985 4471
rect 26985 4437 27019 4471
rect 27019 4437 27028 4471
rect 26976 4428 27028 4437
rect 29000 4471 29052 4480
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 29184 4428 29236 4480
rect 36176 4573 36185 4607
rect 36185 4573 36219 4607
rect 36219 4573 36228 4607
rect 36176 4564 36228 4573
rect 36544 4564 36596 4616
rect 34428 4496 34480 4548
rect 34244 4428 34296 4480
rect 37004 4496 37056 4548
rect 37556 4564 37608 4616
rect 39948 4632 40000 4684
rect 40040 4632 40092 4684
rect 38568 4564 38620 4616
rect 42340 4607 42392 4616
rect 42340 4573 42349 4607
rect 42349 4573 42383 4607
rect 42383 4573 42392 4607
rect 42340 4564 42392 4573
rect 43260 4632 43312 4684
rect 42800 4607 42852 4616
rect 42800 4573 42814 4607
rect 42814 4573 42848 4607
rect 42848 4573 42852 4607
rect 43536 4607 43588 4616
rect 42800 4564 42852 4573
rect 43536 4573 43545 4607
rect 43545 4573 43579 4607
rect 43579 4573 43588 4607
rect 43536 4564 43588 4573
rect 43996 4632 44048 4684
rect 45468 4632 45520 4684
rect 58164 4675 58216 4684
rect 58164 4641 58173 4675
rect 58173 4641 58207 4675
rect 58207 4641 58216 4675
rect 58164 4632 58216 4641
rect 35900 4428 35952 4480
rect 35992 4428 36044 4480
rect 37924 4496 37976 4548
rect 38936 4496 38988 4548
rect 41328 4496 41380 4548
rect 40868 4428 40920 4480
rect 41052 4428 41104 4480
rect 43168 4496 43220 4548
rect 43720 4539 43772 4548
rect 43720 4505 43729 4539
rect 43729 4505 43763 4539
rect 43763 4505 43772 4539
rect 43720 4496 43772 4505
rect 45560 4564 45612 4616
rect 52000 4564 52052 4616
rect 57336 4564 57388 4616
rect 43260 4428 43312 4480
rect 43904 4428 43956 4480
rect 45468 4496 45520 4548
rect 53932 4496 53984 4548
rect 57244 4539 57296 4548
rect 57244 4505 57253 4539
rect 57253 4505 57287 4539
rect 57287 4505 57296 4539
rect 57244 4496 57296 4505
rect 44548 4428 44600 4480
rect 48412 4428 48464 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 5632 4224 5684 4276
rect 7012 4224 7064 4276
rect 12900 4224 12952 4276
rect 3148 4088 3200 4140
rect 3700 4088 3752 4140
rect 4620 4156 4672 4208
rect 6368 4156 6420 4208
rect 7748 4156 7800 4208
rect 7932 4156 7984 4208
rect 8116 4156 8168 4208
rect 6920 4088 6972 4140
rect 8852 4131 8904 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 2872 4020 2924 4072
rect 7932 4020 7984 4072
rect 5356 3952 5408 4004
rect 6460 3952 6512 4004
rect 6552 3952 6604 4004
rect 5540 3884 5592 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 11980 4156 12032 4208
rect 9588 4088 9640 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 8392 4020 8444 4072
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 13544 4156 13596 4208
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 15936 4156 15988 4208
rect 16948 4199 17000 4208
rect 16948 4165 16957 4199
rect 16957 4165 16991 4199
rect 16991 4165 17000 4199
rect 16948 4156 17000 4165
rect 17224 4224 17276 4276
rect 18328 4224 18380 4276
rect 19340 4224 19392 4276
rect 19248 4156 19300 4208
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 20352 4224 20404 4276
rect 20444 4199 20496 4208
rect 20444 4165 20453 4199
rect 20453 4165 20487 4199
rect 20487 4165 20496 4199
rect 20904 4224 20956 4276
rect 22100 4224 22152 4276
rect 22192 4224 22244 4276
rect 24400 4224 24452 4276
rect 20444 4156 20496 4165
rect 21732 4156 21784 4208
rect 22468 4156 22520 4208
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15660 4088 15712 4140
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 19616 4131 19668 4140
rect 19616 4097 19628 4131
rect 19628 4097 19662 4131
rect 19662 4097 19668 4131
rect 20628 4131 20680 4140
rect 19616 4088 19668 4097
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 20812 4088 20864 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 11060 3952 11112 4004
rect 12716 3952 12768 4004
rect 15384 4020 15436 4072
rect 17592 4063 17644 4072
rect 17592 4029 17601 4063
rect 17601 4029 17635 4063
rect 17635 4029 17644 4063
rect 17592 4020 17644 4029
rect 18236 4020 18288 4072
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 9404 3884 9456 3936
rect 10600 3884 10652 3936
rect 12440 3884 12492 3936
rect 12992 3884 13044 3936
rect 20996 3952 21048 4004
rect 21640 3952 21692 4004
rect 22376 4088 22428 4140
rect 24308 4199 24360 4208
rect 24308 4165 24317 4199
rect 24317 4165 24351 4199
rect 24351 4165 24360 4199
rect 24308 4156 24360 4165
rect 22744 4131 22796 4140
rect 22744 4097 22753 4131
rect 22753 4097 22787 4131
rect 22787 4097 22796 4131
rect 22744 4088 22796 4097
rect 23296 4088 23348 4140
rect 23388 4088 23440 4140
rect 29184 4224 29236 4276
rect 29368 4224 29420 4276
rect 32312 4267 32364 4276
rect 32312 4233 32321 4267
rect 32321 4233 32355 4267
rect 32355 4233 32364 4267
rect 32312 4224 32364 4233
rect 32588 4224 32640 4276
rect 35900 4224 35952 4276
rect 36728 4224 36780 4276
rect 39396 4224 39448 4276
rect 45928 4267 45980 4276
rect 24860 4156 24912 4208
rect 27436 4156 27488 4208
rect 27620 4156 27672 4208
rect 28724 4156 28776 4208
rect 28908 4156 28960 4208
rect 29000 4156 29052 4208
rect 35716 4156 35768 4208
rect 37464 4156 37516 4208
rect 38660 4199 38712 4208
rect 38660 4165 38669 4199
rect 38669 4165 38703 4199
rect 38703 4165 38712 4199
rect 45928 4233 45937 4267
rect 45937 4233 45971 4267
rect 45971 4233 45980 4267
rect 45928 4224 45980 4233
rect 53472 4224 53524 4276
rect 38660 4156 38712 4165
rect 42248 4156 42300 4208
rect 25136 4131 25188 4140
rect 25136 4097 25145 4131
rect 25145 4097 25179 4131
rect 25179 4097 25188 4131
rect 25136 4088 25188 4097
rect 25412 4131 25464 4140
rect 25412 4097 25446 4131
rect 25446 4097 25464 4131
rect 25412 4088 25464 4097
rect 25780 4088 25832 4140
rect 27252 4088 27304 4140
rect 24216 4020 24268 4072
rect 24860 4020 24912 4072
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 27896 4020 27948 4072
rect 28356 4063 28408 4072
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 19984 3884 20036 3936
rect 21824 3884 21876 3936
rect 22836 3884 22888 3936
rect 23204 3884 23256 3936
rect 25044 3952 25096 4004
rect 28632 4020 28684 4072
rect 33232 4088 33284 4140
rect 33508 4088 33560 4140
rect 33692 4088 33744 4140
rect 35348 4088 35400 4140
rect 29460 4020 29512 4072
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 29920 4020 29972 4072
rect 36268 4088 36320 4140
rect 36452 4131 36504 4140
rect 36452 4097 36461 4131
rect 36461 4097 36495 4131
rect 36495 4097 36504 4131
rect 36452 4088 36504 4097
rect 37004 4088 37056 4140
rect 38936 4088 38988 4140
rect 39304 4131 39356 4140
rect 39304 4097 39313 4131
rect 39313 4097 39347 4131
rect 39347 4097 39356 4131
rect 39304 4088 39356 4097
rect 39948 4088 40000 4140
rect 42524 4088 42576 4140
rect 43260 4131 43312 4140
rect 43260 4097 43269 4131
rect 43269 4097 43303 4131
rect 43303 4097 43312 4131
rect 43260 4088 43312 4097
rect 43720 4088 43772 4140
rect 45100 4199 45152 4208
rect 45100 4165 45109 4199
rect 45109 4165 45143 4199
rect 45143 4165 45152 4199
rect 45100 4156 45152 4165
rect 45744 4156 45796 4208
rect 48872 4156 48924 4208
rect 50620 4156 50672 4208
rect 51356 4156 51408 4208
rect 52460 4156 52512 4208
rect 53104 4156 53156 4208
rect 57888 4156 57940 4208
rect 44548 4088 44600 4140
rect 46756 4131 46808 4140
rect 46756 4097 46765 4131
rect 46765 4097 46799 4131
rect 46799 4097 46808 4131
rect 46756 4088 46808 4097
rect 48228 4131 48280 4140
rect 48228 4097 48237 4131
rect 48237 4097 48271 4131
rect 48271 4097 48280 4131
rect 48228 4088 48280 4097
rect 48412 4131 48464 4140
rect 48412 4097 48421 4131
rect 48421 4097 48455 4131
rect 48455 4097 48464 4131
rect 48412 4088 48464 4097
rect 49240 4088 49292 4140
rect 50804 4088 50856 4140
rect 51724 4131 51776 4140
rect 51724 4097 51733 4131
rect 51733 4097 51767 4131
rect 51767 4097 51776 4131
rect 51724 4088 51776 4097
rect 53196 4131 53248 4140
rect 53196 4097 53205 4131
rect 53205 4097 53239 4131
rect 53239 4097 53248 4131
rect 53196 4088 53248 4097
rect 53288 4088 53340 4140
rect 54116 4088 54168 4140
rect 31760 3952 31812 4004
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 27160 3884 27212 3893
rect 27344 3884 27396 3936
rect 28448 3884 28500 3936
rect 28540 3884 28592 3936
rect 29184 3927 29236 3936
rect 29184 3893 29193 3927
rect 29193 3893 29227 3927
rect 29227 3893 29236 3927
rect 29184 3884 29236 3893
rect 29920 3884 29972 3936
rect 35900 4020 35952 4072
rect 36360 4020 36412 4072
rect 34796 3952 34848 4004
rect 38752 4020 38804 4072
rect 40408 4020 40460 4072
rect 41512 4020 41564 4072
rect 42984 4020 43036 4072
rect 43536 4063 43588 4072
rect 35348 3884 35400 3936
rect 35624 3884 35676 3936
rect 37924 3952 37976 4004
rect 37648 3927 37700 3936
rect 37648 3893 37657 3927
rect 37657 3893 37691 3927
rect 37691 3893 37700 3927
rect 37648 3884 37700 3893
rect 37740 3884 37792 3936
rect 39120 3952 39172 4004
rect 41144 3952 41196 4004
rect 42800 3952 42852 4004
rect 43536 4029 43545 4063
rect 43545 4029 43579 4063
rect 43579 4029 43588 4063
rect 43536 4020 43588 4029
rect 43812 4020 43864 4072
rect 44456 4020 44508 4072
rect 45376 4020 45428 4072
rect 44548 3952 44600 4004
rect 44732 3952 44784 4004
rect 45652 3952 45704 4004
rect 46572 3952 46624 4004
rect 50896 3952 50948 4004
rect 54300 4020 54352 4072
rect 57980 4088 58032 4140
rect 58348 4131 58400 4140
rect 58348 4097 58357 4131
rect 58357 4097 58391 4131
rect 58391 4097 58400 4131
rect 58348 4088 58400 4097
rect 58256 4020 58308 4072
rect 55312 3995 55364 4004
rect 38752 3927 38804 3936
rect 38752 3893 38761 3927
rect 38761 3893 38795 3927
rect 38795 3893 38804 3927
rect 38752 3884 38804 3893
rect 38844 3884 38896 3936
rect 39948 3884 40000 3936
rect 41420 3884 41472 3936
rect 43536 3884 43588 3936
rect 43628 3884 43680 3936
rect 51540 3884 51592 3936
rect 55312 3961 55321 3995
rect 55321 3961 55355 3995
rect 55355 3961 55364 3995
rect 55312 3952 55364 3961
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3148 3476 3200 3528
rect 5724 3680 5776 3732
rect 7196 3680 7248 3732
rect 4160 3612 4212 3664
rect 5080 3612 5132 3664
rect 8668 3612 8720 3664
rect 9128 3612 9180 3664
rect 6000 3544 6052 3596
rect 7012 3544 7064 3596
rect 7288 3544 7340 3596
rect 14096 3680 14148 3732
rect 17592 3680 17644 3732
rect 19340 3680 19392 3732
rect 22928 3723 22980 3732
rect 10324 3612 10376 3664
rect 11520 3655 11572 3664
rect 11520 3621 11529 3655
rect 11529 3621 11563 3655
rect 11563 3621 11572 3655
rect 11520 3612 11572 3621
rect 11888 3612 11940 3664
rect 4988 3476 5040 3528
rect 7380 3476 7432 3528
rect 9956 3476 10008 3528
rect 10416 3476 10468 3528
rect 14924 3612 14976 3664
rect 16764 3612 16816 3664
rect 18144 3612 18196 3664
rect 18788 3612 18840 3664
rect 15752 3544 15804 3596
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 5908 3340 5960 3392
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 6736 3451 6788 3460
rect 6736 3417 6745 3451
rect 6745 3417 6779 3451
rect 6779 3417 6788 3451
rect 6736 3408 6788 3417
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 8116 3451 8168 3460
rect 8116 3417 8125 3451
rect 8125 3417 8159 3451
rect 8159 3417 8168 3451
rect 8116 3408 8168 3417
rect 8852 3408 8904 3460
rect 13176 3476 13228 3528
rect 13636 3476 13688 3528
rect 14464 3476 14516 3528
rect 12164 3408 12216 3460
rect 13452 3408 13504 3460
rect 8668 3340 8720 3392
rect 14556 3340 14608 3392
rect 15844 3408 15896 3460
rect 16212 3408 16264 3460
rect 17684 3544 17736 3596
rect 19248 3544 19300 3596
rect 22928 3689 22937 3723
rect 22937 3689 22971 3723
rect 22971 3689 22980 3723
rect 22928 3680 22980 3689
rect 24400 3680 24452 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 24860 3680 24912 3732
rect 29184 3680 29236 3732
rect 19708 3612 19760 3664
rect 18052 3476 18104 3528
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 19340 3476 19392 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 16764 3408 16816 3460
rect 18972 3408 19024 3460
rect 19984 3544 20036 3596
rect 23388 3612 23440 3664
rect 28356 3612 28408 3664
rect 31392 3680 31444 3732
rect 20628 3519 20680 3528
rect 20628 3485 20637 3519
rect 20637 3485 20671 3519
rect 20671 3485 20680 3519
rect 20628 3476 20680 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 20904 3476 20956 3528
rect 23020 3544 23072 3596
rect 24676 3544 24728 3596
rect 25780 3587 25832 3596
rect 22284 3476 22336 3528
rect 23204 3476 23256 3528
rect 24860 3476 24912 3528
rect 25780 3553 25789 3587
rect 25789 3553 25823 3587
rect 25823 3553 25832 3587
rect 25780 3544 25832 3553
rect 29460 3544 29512 3596
rect 29552 3544 29604 3596
rect 29736 3587 29788 3596
rect 29736 3553 29745 3587
rect 29745 3553 29779 3587
rect 29779 3553 29788 3587
rect 29736 3544 29788 3553
rect 25688 3476 25740 3528
rect 27160 3476 27212 3528
rect 27252 3476 27304 3528
rect 19064 3340 19116 3392
rect 19708 3383 19760 3392
rect 19708 3349 19717 3383
rect 19717 3349 19751 3383
rect 19751 3349 19760 3383
rect 19708 3340 19760 3349
rect 20720 3408 20772 3460
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 20904 3340 20956 3349
rect 21088 3408 21140 3460
rect 21640 3451 21692 3460
rect 21640 3417 21649 3451
rect 21649 3417 21683 3451
rect 21683 3417 21692 3451
rect 21640 3408 21692 3417
rect 22192 3451 22244 3460
rect 22192 3417 22201 3451
rect 22201 3417 22235 3451
rect 22235 3417 22244 3451
rect 22192 3408 22244 3417
rect 26976 3408 27028 3460
rect 27528 3408 27580 3460
rect 30932 3476 30984 3528
rect 34244 3680 34296 3732
rect 34428 3680 34480 3732
rect 35900 3680 35952 3732
rect 36176 3680 36228 3732
rect 36452 3680 36504 3732
rect 39028 3680 39080 3732
rect 41972 3723 42024 3732
rect 33232 3612 33284 3664
rect 36084 3612 36136 3664
rect 37188 3612 37240 3664
rect 37280 3612 37332 3664
rect 37556 3612 37608 3664
rect 40500 3612 40552 3664
rect 40684 3612 40736 3664
rect 41972 3689 41981 3723
rect 41981 3689 42015 3723
rect 42015 3689 42024 3723
rect 41972 3680 42024 3689
rect 43076 3680 43128 3732
rect 45100 3680 45152 3732
rect 45192 3680 45244 3732
rect 46020 3680 46072 3732
rect 48596 3723 48648 3732
rect 48596 3689 48605 3723
rect 48605 3689 48639 3723
rect 48639 3689 48648 3723
rect 48596 3680 48648 3689
rect 49332 3723 49384 3732
rect 49332 3689 49341 3723
rect 49341 3689 49375 3723
rect 49375 3689 49384 3723
rect 49332 3680 49384 3689
rect 50068 3680 50120 3732
rect 52000 3723 52052 3732
rect 52000 3689 52009 3723
rect 52009 3689 52043 3723
rect 52043 3689 52052 3723
rect 52000 3680 52052 3689
rect 52644 3680 52696 3732
rect 47032 3655 47084 3664
rect 34888 3587 34940 3596
rect 34888 3553 34897 3587
rect 34897 3553 34931 3587
rect 34931 3553 34940 3587
rect 34888 3544 34940 3553
rect 35900 3544 35952 3596
rect 37004 3544 37056 3596
rect 28264 3408 28316 3460
rect 28540 3408 28592 3460
rect 29552 3408 29604 3460
rect 29828 3408 29880 3460
rect 32312 3451 32364 3460
rect 32312 3417 32346 3451
rect 32346 3417 32364 3451
rect 32312 3408 32364 3417
rect 32404 3408 32456 3460
rect 32864 3408 32916 3460
rect 36084 3476 36136 3528
rect 36728 3519 36780 3528
rect 36728 3485 36737 3519
rect 36737 3485 36771 3519
rect 36771 3485 36780 3519
rect 36728 3476 36780 3485
rect 36912 3519 36964 3528
rect 36912 3485 36919 3519
rect 36919 3485 36964 3519
rect 36912 3476 36964 3485
rect 37740 3476 37792 3528
rect 38660 3544 38712 3596
rect 42616 3544 42668 3596
rect 43168 3544 43220 3596
rect 47032 3621 47041 3655
rect 47041 3621 47075 3655
rect 47075 3621 47084 3655
rect 47032 3612 47084 3621
rect 49700 3612 49752 3664
rect 44548 3544 44600 3596
rect 51540 3544 51592 3596
rect 56876 3587 56928 3596
rect 36636 3408 36688 3460
rect 37004 3451 37056 3460
rect 37004 3417 37013 3451
rect 37013 3417 37047 3451
rect 37047 3417 37056 3451
rect 37004 3408 37056 3417
rect 22468 3340 22520 3392
rect 23112 3383 23164 3392
rect 23112 3349 23121 3383
rect 23121 3349 23155 3383
rect 23155 3349 23164 3383
rect 23112 3340 23164 3349
rect 23204 3340 23256 3392
rect 23940 3340 23992 3392
rect 25228 3340 25280 3392
rect 26332 3340 26384 3392
rect 27620 3340 27672 3392
rect 28632 3340 28684 3392
rect 29000 3340 29052 3392
rect 30196 3340 30248 3392
rect 35256 3340 35308 3392
rect 38384 3408 38436 3460
rect 38568 3408 38620 3460
rect 38660 3408 38712 3460
rect 38936 3408 38988 3460
rect 40132 3408 40184 3460
rect 38292 3340 38344 3392
rect 39580 3340 39632 3392
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 41144 3519 41196 3528
rect 41144 3485 41153 3519
rect 41153 3485 41187 3519
rect 41187 3485 41196 3519
rect 42156 3519 42208 3528
rect 41144 3476 41196 3485
rect 42156 3485 42165 3519
rect 42165 3485 42199 3519
rect 42199 3485 42208 3519
rect 42156 3476 42208 3485
rect 42708 3519 42760 3528
rect 41328 3408 41380 3460
rect 42708 3485 42717 3519
rect 42717 3485 42751 3519
rect 42751 3485 42760 3519
rect 42708 3476 42760 3485
rect 42800 3519 42852 3528
rect 42800 3485 42809 3519
rect 42809 3485 42843 3519
rect 42843 3485 42852 3519
rect 42800 3476 42852 3485
rect 43352 3519 43404 3528
rect 43352 3485 43361 3519
rect 43361 3485 43395 3519
rect 43395 3485 43404 3519
rect 43536 3519 43588 3528
rect 43352 3476 43404 3485
rect 43536 3485 43543 3519
rect 43543 3485 43588 3519
rect 43536 3476 43588 3485
rect 43812 3519 43864 3528
rect 43812 3485 43826 3519
rect 43826 3485 43860 3519
rect 43860 3485 43864 3519
rect 43812 3476 43864 3485
rect 43260 3408 43312 3460
rect 45008 3476 45060 3528
rect 46020 3519 46072 3528
rect 46020 3485 46029 3519
rect 46029 3485 46063 3519
rect 46063 3485 46072 3519
rect 46020 3476 46072 3485
rect 44548 3408 44600 3460
rect 45468 3408 45520 3460
rect 49148 3476 49200 3528
rect 46664 3408 46716 3460
rect 47124 3408 47176 3460
rect 48136 3408 48188 3460
rect 45192 3340 45244 3392
rect 50712 3476 50764 3528
rect 49516 3408 49568 3460
rect 50804 3408 50856 3460
rect 52000 3476 52052 3528
rect 51632 3408 51684 3460
rect 52736 3408 52788 3460
rect 53932 3408 53984 3460
rect 51816 3340 51868 3392
rect 53472 3383 53524 3392
rect 53472 3349 53481 3383
rect 53481 3349 53515 3383
rect 53515 3349 53524 3383
rect 53472 3340 53524 3349
rect 53656 3340 53708 3392
rect 56876 3553 56885 3587
rect 56885 3553 56919 3587
rect 56919 3553 56928 3587
rect 56876 3544 56928 3553
rect 56232 3451 56284 3460
rect 56232 3417 56241 3451
rect 56241 3417 56275 3451
rect 56275 3417 56284 3451
rect 56232 3408 56284 3417
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4160 3136 4212 3188
rect 6552 3136 6604 3188
rect 9036 3136 9088 3188
rect 4804 3068 4856 3120
rect 7288 3111 7340 3120
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4712 3000 4764 3052
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 8116 3068 8168 3120
rect 17684 3136 17736 3188
rect 17776 3136 17828 3188
rect 18788 3136 18840 3188
rect 19248 3136 19300 3188
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 9220 3000 9272 3052
rect 10232 3000 10284 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 12532 3000 12584 3052
rect 13728 3000 13780 3052
rect 13912 3000 13964 3052
rect 14740 3043 14792 3052
rect 6092 2864 6144 2916
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 5816 2796 5868 2848
rect 10140 2932 10192 2984
rect 9864 2864 9916 2916
rect 12072 2864 12124 2916
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 16580 3068 16632 3120
rect 16764 3068 16816 3120
rect 15200 3000 15252 3052
rect 17132 3043 17184 3052
rect 15292 2932 15344 2984
rect 15476 2864 15528 2916
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 16948 2864 17000 2916
rect 18052 2932 18104 2984
rect 18880 3000 18932 3052
rect 20444 3068 20496 3120
rect 20996 3136 21048 3188
rect 21364 3068 21416 3120
rect 21456 3068 21508 3120
rect 22560 3068 22612 3120
rect 19524 3000 19576 3052
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 19800 3000 19852 3052
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 11060 2796 11112 2848
rect 14556 2796 14608 2848
rect 15016 2796 15068 2848
rect 15384 2796 15436 2848
rect 19432 2796 19484 2848
rect 20352 2864 20404 2916
rect 20536 3000 20588 3052
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 20720 2932 20772 2984
rect 21364 2932 21416 2984
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 23572 3136 23624 3188
rect 25412 3136 25464 3188
rect 25504 3179 25556 3188
rect 25504 3145 25513 3179
rect 25513 3145 25547 3179
rect 25547 3145 25556 3179
rect 25504 3136 25556 3145
rect 27436 3136 27488 3188
rect 26332 3068 26384 3120
rect 27620 3068 27672 3120
rect 29184 3136 29236 3188
rect 29552 3136 29604 3188
rect 29828 3136 29880 3188
rect 30012 3136 30064 3188
rect 28264 3068 28316 3120
rect 32036 3136 32088 3188
rect 33232 3136 33284 3188
rect 36084 3136 36136 3188
rect 36268 3179 36320 3188
rect 36268 3145 36277 3179
rect 36277 3145 36311 3179
rect 36311 3145 36320 3179
rect 36268 3136 36320 3145
rect 36452 3136 36504 3188
rect 39488 3179 39540 3188
rect 30472 3068 30524 3120
rect 30748 3068 30800 3120
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 23296 3043 23348 3052
rect 22928 3000 22980 3009
rect 23296 3009 23305 3043
rect 23305 3009 23339 3043
rect 23339 3009 23348 3043
rect 23296 3000 23348 3009
rect 24032 3000 24084 3052
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 23756 2932 23808 2984
rect 25596 2975 25648 2984
rect 20812 2864 20864 2916
rect 22468 2864 22520 2916
rect 22744 2907 22796 2916
rect 22744 2873 22753 2907
rect 22753 2873 22787 2907
rect 22787 2873 22796 2907
rect 22744 2864 22796 2873
rect 24400 2864 24452 2916
rect 25596 2941 25605 2975
rect 25605 2941 25639 2975
rect 25639 2941 25648 2975
rect 25596 2932 25648 2941
rect 25688 2932 25740 2984
rect 28356 3000 28408 3052
rect 29920 3000 29972 3052
rect 30288 3000 30340 3052
rect 30196 2932 30248 2984
rect 31300 3043 31352 3052
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31300 3000 31352 3009
rect 32312 3043 32364 3052
rect 32312 3009 32321 3043
rect 32321 3009 32355 3043
rect 32355 3009 32364 3043
rect 32312 3000 32364 3009
rect 32496 3068 32548 3120
rect 33968 3068 34020 3120
rect 34152 3000 34204 3052
rect 34428 3043 34480 3052
rect 31208 2932 31260 2984
rect 31760 2932 31812 2984
rect 28356 2907 28408 2916
rect 22376 2796 22428 2848
rect 25136 2796 25188 2848
rect 28356 2873 28365 2907
rect 28365 2873 28399 2907
rect 28399 2873 28408 2907
rect 28356 2864 28408 2873
rect 28632 2864 28684 2916
rect 34428 3009 34437 3043
rect 34437 3009 34471 3043
rect 34471 3009 34480 3043
rect 34428 3000 34480 3009
rect 34888 3043 34940 3052
rect 34888 3009 34897 3043
rect 34897 3009 34931 3043
rect 34931 3009 34940 3043
rect 34888 3000 34940 3009
rect 35348 3068 35400 3120
rect 35440 3068 35492 3120
rect 39488 3145 39497 3179
rect 39497 3145 39531 3179
rect 39531 3145 39540 3179
rect 39488 3136 39540 3145
rect 40592 3179 40644 3188
rect 40592 3145 40601 3179
rect 40601 3145 40635 3179
rect 40635 3145 40644 3179
rect 40592 3136 40644 3145
rect 41144 3136 41196 3188
rect 41880 3068 41932 3120
rect 42432 3068 42484 3120
rect 38200 3000 38252 3052
rect 38844 3000 38896 3052
rect 39120 3000 39172 3052
rect 39764 3000 39816 3052
rect 36544 2864 36596 2916
rect 38292 2932 38344 2984
rect 37832 2864 37884 2916
rect 43260 3043 43312 3052
rect 43260 3009 43269 3043
rect 43269 3009 43303 3043
rect 43303 3009 43312 3043
rect 43628 3043 43680 3052
rect 43260 3000 43312 3009
rect 43628 3009 43637 3043
rect 43637 3009 43671 3043
rect 43671 3009 43680 3043
rect 43628 3000 43680 3009
rect 43812 3043 43864 3052
rect 43812 3009 43821 3043
rect 43821 3009 43855 3043
rect 43855 3009 43864 3043
rect 44640 3136 44692 3188
rect 45192 3179 45244 3188
rect 45192 3145 45201 3179
rect 45201 3145 45235 3179
rect 45235 3145 45244 3179
rect 45192 3136 45244 3145
rect 46388 3179 46440 3188
rect 46388 3145 46397 3179
rect 46397 3145 46431 3179
rect 46431 3145 46440 3179
rect 46388 3136 46440 3145
rect 47400 3136 47452 3188
rect 48044 3136 48096 3188
rect 50252 3136 50304 3188
rect 50712 3136 50764 3188
rect 51264 3179 51316 3188
rect 51264 3145 51273 3179
rect 51273 3145 51307 3179
rect 51307 3145 51316 3179
rect 51264 3136 51316 3145
rect 51816 3136 51868 3188
rect 53840 3179 53892 3188
rect 45468 3068 45520 3120
rect 47492 3068 47544 3120
rect 49884 3068 49936 3120
rect 53840 3145 53849 3179
rect 53849 3145 53883 3179
rect 53883 3145 53892 3179
rect 53840 3136 53892 3145
rect 54760 3179 54812 3188
rect 54760 3145 54769 3179
rect 54769 3145 54803 3179
rect 54803 3145 54812 3179
rect 54760 3136 54812 3145
rect 58256 3179 58308 3188
rect 58256 3145 58265 3179
rect 58265 3145 58299 3179
rect 58299 3145 58308 3179
rect 58256 3136 58308 3145
rect 43812 3000 43864 3009
rect 44456 3000 44508 3052
rect 46112 3000 46164 3052
rect 47032 3000 47084 3052
rect 45284 2932 45336 2984
rect 48136 3000 48188 3052
rect 48596 3000 48648 3052
rect 48964 3000 49016 3052
rect 48044 2932 48096 2984
rect 51172 3000 51224 3052
rect 53656 3068 53708 3120
rect 55680 3068 55732 3120
rect 58164 3111 58216 3120
rect 58164 3077 58173 3111
rect 58173 3077 58207 3111
rect 58207 3077 58216 3111
rect 58164 3068 58216 3077
rect 53564 3000 53616 3052
rect 53840 3000 53892 3052
rect 54944 3000 54996 3052
rect 50896 2932 50948 2984
rect 53380 2932 53432 2984
rect 55772 2932 55824 2984
rect 26792 2796 26844 2848
rect 31668 2796 31720 2848
rect 32036 2796 32088 2848
rect 33416 2796 33468 2848
rect 37004 2796 37056 2848
rect 40132 2796 40184 2848
rect 40868 2796 40920 2848
rect 41604 2796 41656 2848
rect 45284 2796 45336 2848
rect 48964 2796 49016 2848
rect 49056 2839 49108 2848
rect 49056 2805 49065 2839
rect 49065 2805 49099 2839
rect 49099 2805 49108 2839
rect 49056 2796 49108 2805
rect 49700 2796 49752 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 9588 2592 9640 2644
rect 7564 2524 7616 2576
rect 7840 2524 7892 2576
rect 8484 2567 8536 2576
rect 8484 2533 8493 2567
rect 8493 2533 8527 2567
rect 8527 2533 8536 2567
rect 8484 2524 8536 2533
rect 12716 2592 12768 2644
rect 14740 2592 14792 2644
rect 18052 2592 18104 2644
rect 18972 2592 19024 2644
rect 19708 2592 19760 2644
rect 21456 2592 21508 2644
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 9312 2431 9364 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 4896 2320 4948 2372
rect 5080 2363 5132 2372
rect 5080 2329 5089 2363
rect 5089 2329 5123 2363
rect 5123 2329 5132 2363
rect 5080 2320 5132 2329
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6736 2363 6788 2372
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 7012 2320 7064 2372
rect 8116 2363 8168 2372
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 8116 2329 8125 2363
rect 8125 2329 8159 2363
rect 8159 2329 8168 2363
rect 8116 2320 8168 2329
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10876 2524 10928 2576
rect 14556 2524 14608 2576
rect 15016 2524 15068 2576
rect 23296 2592 23348 2644
rect 24768 2592 24820 2644
rect 25044 2592 25096 2644
rect 25504 2592 25556 2644
rect 22008 2567 22060 2576
rect 22008 2533 22017 2567
rect 22017 2533 22051 2567
rect 22051 2533 22060 2567
rect 22008 2524 22060 2533
rect 23020 2567 23072 2576
rect 23020 2533 23029 2567
rect 23029 2533 23063 2567
rect 23063 2533 23072 2567
rect 23020 2524 23072 2533
rect 23112 2524 23164 2576
rect 12716 2456 12768 2508
rect 18052 2456 18104 2508
rect 19156 2456 19208 2508
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14740 2388 14792 2440
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 16028 2388 16080 2440
rect 16396 2388 16448 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18512 2388 18564 2440
rect 18604 2388 18656 2440
rect 19984 2431 20036 2440
rect 9680 2320 9732 2372
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 13360 2320 13412 2372
rect 13544 2363 13596 2372
rect 13544 2329 13553 2363
rect 13553 2329 13587 2363
rect 13587 2329 13596 2363
rect 13544 2320 13596 2329
rect 15936 2320 15988 2372
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 17776 2363 17828 2372
rect 17776 2329 17785 2363
rect 17785 2329 17819 2363
rect 17819 2329 17828 2363
rect 17776 2320 17828 2329
rect 18696 2363 18748 2372
rect 18696 2329 18705 2363
rect 18705 2329 18739 2363
rect 18739 2329 18748 2363
rect 18696 2320 18748 2329
rect 14372 2252 14424 2304
rect 19248 2252 19300 2304
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 19524 2320 19576 2372
rect 20076 2320 20128 2372
rect 20260 2363 20312 2372
rect 20260 2329 20269 2363
rect 20269 2329 20303 2363
rect 20303 2329 20312 2363
rect 20260 2320 20312 2329
rect 22284 2431 22336 2440
rect 22284 2397 22313 2431
rect 22313 2397 22336 2431
rect 22468 2456 22520 2508
rect 25596 2524 25648 2576
rect 29368 2592 29420 2644
rect 31668 2592 31720 2644
rect 33600 2592 33652 2644
rect 34336 2592 34388 2644
rect 22284 2388 22336 2397
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 26332 2456 26384 2508
rect 26884 2456 26936 2508
rect 23572 2363 23624 2372
rect 23572 2329 23581 2363
rect 23581 2329 23615 2363
rect 23615 2329 23624 2363
rect 23572 2320 23624 2329
rect 26332 2320 26384 2372
rect 27804 2388 27856 2440
rect 28356 2388 28408 2440
rect 33048 2524 33100 2576
rect 30380 2456 30432 2508
rect 37648 2592 37700 2644
rect 40224 2635 40276 2644
rect 40224 2601 40233 2635
rect 40233 2601 40267 2635
rect 40267 2601 40276 2635
rect 40224 2592 40276 2601
rect 41328 2635 41380 2644
rect 41328 2601 41337 2635
rect 41337 2601 41371 2635
rect 41371 2601 41380 2635
rect 41328 2592 41380 2601
rect 42800 2635 42852 2644
rect 42800 2601 42809 2635
rect 42809 2601 42843 2635
rect 42843 2601 42852 2635
rect 42800 2592 42852 2601
rect 45836 2635 45888 2644
rect 45836 2601 45845 2635
rect 45845 2601 45879 2635
rect 45879 2601 45888 2635
rect 45836 2592 45888 2601
rect 46940 2635 46992 2644
rect 46940 2601 46949 2635
rect 46949 2601 46983 2635
rect 46983 2601 46992 2635
rect 46940 2592 46992 2601
rect 47952 2635 48004 2644
rect 47952 2601 47961 2635
rect 47961 2601 47995 2635
rect 47995 2601 48004 2635
rect 47952 2592 48004 2601
rect 49424 2592 49476 2644
rect 50160 2592 50212 2644
rect 54024 2635 54076 2644
rect 54024 2601 54033 2635
rect 54033 2601 54067 2635
rect 54067 2601 54076 2635
rect 54024 2592 54076 2601
rect 57980 2592 58032 2644
rect 29276 2388 29328 2440
rect 31944 2388 31996 2440
rect 32772 2388 32824 2440
rect 34060 2388 34112 2440
rect 34244 2388 34296 2440
rect 37280 2524 37332 2576
rect 36084 2499 36136 2508
rect 36084 2465 36093 2499
rect 36093 2465 36127 2499
rect 36127 2465 36136 2499
rect 36084 2456 36136 2465
rect 38476 2524 38528 2576
rect 38568 2524 38620 2576
rect 38752 2456 38804 2508
rect 40132 2456 40184 2508
rect 41420 2388 41472 2440
rect 44364 2456 44416 2508
rect 55404 2456 55456 2508
rect 29828 2320 29880 2372
rect 30656 2320 30708 2372
rect 30932 2320 30984 2372
rect 31484 2320 31536 2372
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 21364 2252 21416 2304
rect 23480 2252 23532 2304
rect 25596 2295 25648 2304
rect 25596 2261 25605 2295
rect 25605 2261 25639 2295
rect 25639 2261 25648 2295
rect 26516 2295 26568 2304
rect 25596 2252 25648 2261
rect 26516 2261 26525 2295
rect 26525 2261 26559 2295
rect 26559 2261 26568 2295
rect 26516 2252 26568 2261
rect 32036 2252 32088 2304
rect 33784 2320 33836 2372
rect 35256 2320 35308 2372
rect 38660 2363 38712 2372
rect 38660 2329 38669 2363
rect 38669 2329 38703 2363
rect 38703 2329 38712 2363
rect 38660 2320 38712 2329
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 41236 2320 41288 2372
rect 43444 2363 43496 2372
rect 43444 2329 43453 2363
rect 43453 2329 43487 2363
rect 43487 2329 43496 2363
rect 43444 2320 43496 2329
rect 46388 2388 46440 2440
rect 45560 2320 45612 2372
rect 45836 2320 45888 2372
rect 47216 2320 47268 2372
rect 48044 2320 48096 2372
rect 49976 2320 50028 2372
rect 54668 2388 54720 2440
rect 56416 2431 56468 2440
rect 56416 2397 56425 2431
rect 56425 2397 56459 2431
rect 56459 2397 56468 2431
rect 56416 2388 56468 2397
rect 57888 2388 57940 2440
rect 33600 2252 33652 2304
rect 43536 2295 43588 2304
rect 43536 2261 43545 2295
rect 43545 2261 43579 2295
rect 43579 2261 43588 2295
rect 43536 2252 43588 2261
rect 48320 2252 48372 2304
rect 52184 2320 52236 2372
rect 53288 2320 53340 2372
rect 51264 2295 51316 2304
rect 51264 2261 51273 2295
rect 51273 2261 51307 2295
rect 51307 2261 51316 2295
rect 51264 2252 51316 2261
rect 53104 2295 53156 2304
rect 53104 2261 53113 2295
rect 53113 2261 53147 2295
rect 53147 2261 53156 2295
rect 53104 2252 53156 2261
rect 55496 2252 55548 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 9312 2048 9364 2100
rect 17224 2048 17276 2100
rect 18696 2048 18748 2100
rect 29000 2048 29052 2100
rect 29368 2048 29420 2100
rect 5816 1980 5868 2032
rect 13268 1980 13320 2032
rect 5080 1912 5132 1964
rect 11888 1912 11940 1964
rect 12348 1912 12400 1964
rect 15568 1980 15620 2032
rect 17776 1980 17828 2032
rect 28448 1980 28500 2032
rect 33416 2048 33468 2100
rect 35256 2048 35308 2100
rect 36728 2048 36780 2100
rect 43444 2048 43496 2100
rect 43904 2048 43956 2100
rect 45744 2048 45796 2100
rect 34152 1980 34204 2032
rect 34244 1980 34296 2032
rect 38660 1980 38712 2032
rect 13544 1912 13596 1964
rect 22928 1912 22980 1964
rect 31576 1912 31628 1964
rect 51264 1912 51316 1964
rect 7012 1844 7064 1896
rect 12808 1844 12860 1896
rect 18420 1844 18472 1896
rect 19892 1844 19944 1896
rect 20260 1844 20312 1896
rect 29276 1844 29328 1896
rect 29644 1844 29696 1896
rect 53104 1844 53156 1896
rect 6736 1776 6788 1828
rect 13544 1776 13596 1828
rect 15936 1776 15988 1828
rect 24584 1776 24636 1828
rect 26516 1776 26568 1828
rect 56416 1776 56468 1828
rect 4896 1708 4948 1760
rect 11336 1708 11388 1760
rect 12716 1708 12768 1760
rect 20444 1708 20496 1760
rect 20628 1708 20680 1760
rect 23480 1708 23532 1760
rect 24216 1708 24268 1760
rect 53472 1708 53524 1760
rect 5172 1572 5224 1624
rect 11428 1640 11480 1692
rect 16120 1640 16172 1692
rect 28172 1640 28224 1692
rect 39488 1640 39540 1692
rect 46020 1640 46072 1692
rect 10968 1572 11020 1624
rect 17960 1572 18012 1624
rect 19248 1572 19300 1624
rect 27896 1572 27948 1624
rect 1584 1504 1636 1556
rect 15108 1504 15160 1556
rect 15844 1504 15896 1556
rect 28264 1504 28316 1556
rect 4712 1436 4764 1488
rect 8300 1436 8352 1488
rect 10600 1436 10652 1488
rect 17408 1436 17460 1488
rect 20352 1436 20404 1488
rect 23204 1436 23256 1488
rect 3332 1368 3384 1420
rect 11152 1368 11204 1420
rect 13360 1368 13412 1420
rect 19248 1368 19300 1420
rect 20076 1368 20128 1420
rect 20996 1368 21048 1420
rect 22284 1368 22336 1420
rect 40776 1436 40828 1488
rect 43352 1436 43404 1488
rect 47124 1436 47176 1488
rect 32588 1368 32640 1420
rect 33784 1368 33836 1420
rect 37280 1368 37332 1420
rect 38568 1368 38620 1420
rect 16948 1300 17000 1352
rect 40960 1300 41012 1352
rect 13452 1232 13504 1284
rect 23572 1232 23624 1284
rect 10692 1164 10744 1216
rect 33508 1164 33560 1216
rect 42524 1164 42576 1216
rect 44548 1164 44600 1216
rect 3608 1096 3660 1148
rect 7196 1096 7248 1148
rect 8668 1096 8720 1148
rect 29184 1096 29236 1148
rect 4988 1028 5040 1080
rect 24768 1028 24820 1080
rect 6460 960 6512 1012
rect 24400 960 24452 1012
rect 5356 892 5408 944
rect 23388 892 23440 944
rect 3148 824 3200 876
rect 22744 824 22796 876
rect 6184 756 6236 808
rect 24492 756 24544 808
rect 4804 688 4856 740
rect 28632 688 28684 740
rect 2320 620 2372 672
rect 21640 620 21692 672
rect 18972 552 19024 604
rect 25780 552 25832 604
rect 18880 484 18932 536
rect 24216 484 24268 536
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63322 2374 64000
rect 3054 63322 3110 64000
rect 3790 63322 3846 64000
rect 4526 63322 4582 64000
rect 5262 63322 5318 64000
rect 2318 63294 2636 63322
rect 2318 63200 2374 63294
rect 860 59022 888 63200
rect 1596 61962 1624 63200
rect 1596 61934 1808 61962
rect 1674 61840 1730 61849
rect 1674 61775 1730 61784
rect 1688 61198 1716 61775
rect 1676 61192 1728 61198
rect 1676 61134 1728 61140
rect 1584 60716 1636 60722
rect 1584 60658 1636 60664
rect 1596 60489 1624 60658
rect 1582 60480 1638 60489
rect 1582 60415 1638 60424
rect 1676 60036 1728 60042
rect 1676 59978 1728 59984
rect 1688 59809 1716 59978
rect 1674 59800 1730 59809
rect 1674 59735 1730 59744
rect 1780 59702 1808 61934
rect 2608 60110 2636 63294
rect 3054 63294 3188 63322
rect 3054 63200 3110 63294
rect 2780 61192 2832 61198
rect 2778 61160 2780 61169
rect 2832 61160 2834 61169
rect 2778 61095 2834 61104
rect 3160 60722 3188 63294
rect 3790 63294 4016 63322
rect 3790 63200 3846 63294
rect 3988 60790 4016 63294
rect 4526 63294 4752 63322
rect 4526 63200 4582 63294
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4724 61198 4752 63294
rect 5262 63294 5488 63322
rect 5262 63200 5318 63294
rect 4712 61192 4764 61198
rect 4712 61134 4764 61140
rect 5460 60790 5488 63294
rect 5998 63200 6054 64000
rect 6734 63322 6790 64000
rect 6656 63294 6790 63322
rect 6012 61198 6040 63200
rect 6276 61328 6328 61334
rect 6276 61270 6328 61276
rect 6000 61192 6052 61198
rect 6000 61134 6052 61140
rect 5540 61124 5592 61130
rect 5540 61066 5592 61072
rect 3976 60784 4028 60790
rect 3976 60726 4028 60732
rect 5448 60784 5500 60790
rect 5448 60726 5500 60732
rect 3148 60716 3200 60722
rect 3148 60658 3200 60664
rect 4804 60648 4856 60654
rect 4804 60590 4856 60596
rect 4620 60580 4672 60586
rect 4620 60522 4672 60528
rect 3332 60512 3384 60518
rect 3332 60454 3384 60460
rect 2596 60104 2648 60110
rect 2596 60046 2648 60052
rect 2044 60036 2096 60042
rect 2044 59978 2096 59984
rect 1768 59696 1820 59702
rect 1768 59638 1820 59644
rect 1584 59628 1636 59634
rect 1584 59570 1636 59576
rect 1596 59129 1624 59570
rect 1768 59424 1820 59430
rect 1768 59366 1820 59372
rect 1780 59226 1808 59366
rect 1768 59220 1820 59226
rect 1768 59162 1820 59168
rect 1582 59120 1638 59129
rect 1582 59055 1638 59064
rect 848 59016 900 59022
rect 848 58958 900 58964
rect 1584 58540 1636 58546
rect 1584 58482 1636 58488
rect 1596 58449 1624 58482
rect 2056 58478 2084 59978
rect 2504 59968 2556 59974
rect 2504 59910 2556 59916
rect 2320 59424 2372 59430
rect 2320 59366 2372 59372
rect 1768 58472 1820 58478
rect 1582 58440 1638 58449
rect 1768 58414 1820 58420
rect 2044 58472 2096 58478
rect 2044 58414 2096 58420
rect 1582 58375 1638 58384
rect 1584 57928 1636 57934
rect 1584 57870 1636 57876
rect 1596 57769 1624 57870
rect 1582 57760 1638 57769
rect 1582 57695 1638 57704
rect 1584 57452 1636 57458
rect 1584 57394 1636 57400
rect 1596 57089 1624 57394
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1584 56840 1636 56846
rect 1584 56782 1636 56788
rect 1596 56409 1624 56782
rect 1582 56400 1638 56409
rect 1582 56335 1638 56344
rect 1674 55720 1730 55729
rect 1674 55655 1676 55664
rect 1728 55655 1730 55664
rect 1676 55626 1728 55632
rect 1584 55276 1636 55282
rect 1584 55218 1636 55224
rect 1596 55049 1624 55218
rect 1582 55040 1638 55049
rect 1582 54975 1638 54984
rect 1676 54596 1728 54602
rect 1676 54538 1728 54544
rect 1688 54369 1716 54538
rect 1674 54360 1730 54369
rect 1674 54295 1730 54304
rect 1584 54188 1636 54194
rect 1584 54130 1636 54136
rect 1596 53689 1624 54130
rect 1582 53680 1638 53689
rect 1582 53615 1638 53624
rect 1676 53100 1728 53106
rect 1676 53042 1728 53048
rect 1688 53009 1716 53042
rect 1674 53000 1730 53009
rect 1674 52935 1730 52944
rect 1584 52488 1636 52494
rect 1584 52430 1636 52436
rect 1596 52329 1624 52430
rect 1582 52320 1638 52329
rect 1582 52255 1638 52264
rect 1676 52012 1728 52018
rect 1676 51954 1728 51960
rect 1688 51649 1716 51954
rect 1674 51640 1730 51649
rect 1674 51575 1730 51584
rect 1676 51332 1728 51338
rect 1676 51274 1728 51280
rect 1688 50969 1716 51274
rect 1674 50960 1730 50969
rect 1674 50895 1730 50904
rect 1674 50280 1730 50289
rect 1674 50215 1676 50224
rect 1728 50215 1730 50224
rect 1676 50186 1728 50192
rect 1584 49836 1636 49842
rect 1584 49778 1636 49784
rect 1596 49609 1624 49778
rect 1582 49600 1638 49609
rect 1582 49535 1638 49544
rect 1676 49156 1728 49162
rect 1676 49098 1728 49104
rect 1688 48929 1716 49098
rect 1674 48920 1730 48929
rect 1674 48855 1730 48864
rect 1676 48748 1728 48754
rect 1676 48690 1728 48696
rect 1688 48249 1716 48690
rect 1674 48240 1730 48249
rect 1674 48175 1730 48184
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1688 47569 1716 47602
rect 1674 47560 1730 47569
rect 1780 47546 1808 58414
rect 1858 52592 1914 52601
rect 1858 52527 1860 52536
rect 1912 52527 1914 52536
rect 1860 52498 1912 52504
rect 2044 50244 2096 50250
rect 2044 50186 2096 50192
rect 1952 48612 2004 48618
rect 1952 48554 2004 48560
rect 1858 47560 1914 47569
rect 1780 47518 1858 47546
rect 1674 47495 1730 47504
rect 1858 47495 1914 47504
rect 1584 47048 1636 47054
rect 1584 46990 1636 46996
rect 1596 46889 1624 46990
rect 1582 46880 1638 46889
rect 1582 46815 1638 46824
rect 1584 46572 1636 46578
rect 1584 46514 1636 46520
rect 1596 46209 1624 46514
rect 1582 46200 1638 46209
rect 1582 46135 1638 46144
rect 1676 45892 1728 45898
rect 1676 45834 1728 45840
rect 1688 45529 1716 45834
rect 1674 45520 1730 45529
rect 1674 45455 1730 45464
rect 1584 44872 1636 44878
rect 1582 44840 1584 44849
rect 1636 44840 1638 44849
rect 1582 44775 1638 44784
rect 1676 44396 1728 44402
rect 1676 44338 1728 44344
rect 1688 44169 1716 44338
rect 1674 44160 1730 44169
rect 1674 44095 1730 44104
rect 1676 43716 1728 43722
rect 1676 43658 1728 43664
rect 1688 43489 1716 43658
rect 1674 43480 1730 43489
rect 1674 43415 1730 43424
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1596 42809 1624 43250
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1582 42800 1638 42809
rect 1582 42735 1638 42744
rect 1780 42702 1808 43046
rect 1768 42696 1820 42702
rect 1768 42638 1820 42644
rect 1676 42220 1728 42226
rect 1676 42162 1728 42168
rect 1688 42129 1716 42162
rect 1674 42120 1730 42129
rect 1674 42055 1730 42064
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41449 1716 41482
rect 1860 41472 1912 41478
rect 1674 41440 1730 41449
rect 1860 41414 1912 41420
rect 1674 41375 1730 41384
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 1688 40769 1716 41074
rect 1674 40760 1730 40769
rect 1674 40695 1730 40704
rect 1676 40452 1728 40458
rect 1676 40394 1728 40400
rect 1688 40089 1716 40394
rect 1674 40080 1730 40089
rect 1674 40015 1730 40024
rect 1674 39400 1730 39409
rect 1674 39335 1676 39344
rect 1728 39335 1730 39344
rect 1676 39306 1728 39312
rect 1676 38956 1728 38962
rect 1676 38898 1728 38904
rect 1688 38729 1716 38898
rect 1674 38720 1730 38729
rect 1674 38655 1730 38664
rect 1676 38276 1728 38282
rect 1676 38218 1728 38224
rect 1688 38049 1716 38218
rect 1674 38040 1730 38049
rect 1674 37975 1730 37984
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 1688 37369 1716 37810
rect 1674 37360 1730 37369
rect 1674 37295 1730 37304
rect 1676 36100 1728 36106
rect 1676 36042 1728 36048
rect 1688 36009 1716 36042
rect 1674 36000 1730 36009
rect 1674 35935 1730 35944
rect 1872 35894 1900 41414
rect 1964 36786 1992 48554
rect 2056 37262 2084 50186
rect 2332 39438 2360 59366
rect 2320 39432 2372 39438
rect 2320 39374 2372 39380
rect 2044 37256 2096 37262
rect 2044 37198 2096 37204
rect 2228 37188 2280 37194
rect 2228 37130 2280 37136
rect 2320 37188 2372 37194
rect 2320 37130 2372 37136
rect 2136 36848 2188 36854
rect 2136 36790 2188 36796
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 1872 35866 1992 35894
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1688 35329 1716 35634
rect 1674 35320 1730 35329
rect 1674 35255 1730 35264
rect 1676 35012 1728 35018
rect 1676 34954 1728 34960
rect 1688 34649 1716 34954
rect 1674 34640 1730 34649
rect 1674 34575 1730 34584
rect 1674 33960 1730 33969
rect 1674 33895 1676 33904
rect 1728 33895 1730 33904
rect 1676 33866 1728 33872
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1688 33289 1716 33458
rect 1674 33280 1730 33289
rect 1674 33215 1730 33224
rect 1676 32836 1728 32842
rect 1676 32778 1728 32784
rect 1688 32609 1716 32778
rect 1674 32600 1730 32609
rect 1674 32535 1730 32544
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 31929 1716 32370
rect 1674 31920 1730 31929
rect 1674 31855 1730 31864
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1688 31249 1716 31282
rect 1674 31240 1730 31249
rect 1674 31175 1730 31184
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1780 30938 1808 31078
rect 1768 30932 1820 30938
rect 1768 30874 1820 30880
rect 1676 30660 1728 30666
rect 1676 30602 1728 30608
rect 1688 30569 1716 30602
rect 1674 30560 1730 30569
rect 1674 30495 1730 30504
rect 1768 30184 1820 30190
rect 1768 30126 1820 30132
rect 1780 29889 1808 30126
rect 1766 29880 1822 29889
rect 1766 29815 1822 29824
rect 1860 29572 1912 29578
rect 1860 29514 1912 29520
rect 1872 29209 1900 29514
rect 1858 29200 1914 29209
rect 1858 29135 1914 29144
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1858 28520 1914 28529
rect 1596 28218 1624 28494
rect 1858 28455 1860 28464
rect 1912 28455 1914 28464
rect 1860 28426 1912 28432
rect 1584 28212 1636 28218
rect 1584 28154 1636 28160
rect 1768 28008 1820 28014
rect 1768 27950 1820 27956
rect 1780 27849 1808 27950
rect 1766 27840 1822 27849
rect 1766 27775 1822 27784
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 27130 1624 27406
rect 1860 27396 1912 27402
rect 1860 27338 1912 27344
rect 1872 27169 1900 27338
rect 1858 27160 1914 27169
rect 1584 27124 1636 27130
rect 1858 27095 1914 27104
rect 1584 27066 1636 27072
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 1780 26489 1808 26862
rect 1766 26480 1822 26489
rect 1766 26415 1822 26424
rect 1768 25832 1820 25838
rect 1766 25800 1768 25809
rect 1820 25800 1822 25809
rect 1766 25735 1822 25744
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1872 25129 1900 25162
rect 1858 25120 1914 25129
rect 1858 25055 1914 25064
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24410 1624 24754
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 1780 24449 1808 24686
rect 1766 24440 1822 24449
rect 1584 24404 1636 24410
rect 1766 24375 1822 24384
rect 1584 24346 1636 24352
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1872 23769 1900 24074
rect 1858 23760 1914 23769
rect 1858 23695 1914 23704
rect 1858 23080 1914 23089
rect 1858 23015 1860 23024
rect 1912 23015 1914 23024
rect 1860 22986 1912 22992
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1780 22409 1808 22510
rect 1766 22400 1822 22409
rect 1766 22335 1822 22344
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1872 21729 1900 21898
rect 1858 21720 1914 21729
rect 1858 21655 1914 21664
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21049 1808 21286
rect 1766 21040 1822 21049
rect 1766 20975 1822 20984
rect 1768 20392 1820 20398
rect 1766 20360 1768 20369
rect 1820 20360 1822 20369
rect 1766 20295 1822 20304
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1872 19689 1900 19722
rect 1858 19680 1914 19689
rect 1858 19615 1914 19624
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 19009 1900 19314
rect 1858 19000 1914 19009
rect 1858 18935 1914 18944
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18329 1900 18634
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1858 17640 1914 17649
rect 1858 17575 1860 17584
rect 1912 17575 1914 17584
rect 1860 17546 1912 17552
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1780 16969 1808 17070
rect 1766 16960 1822 16969
rect 1766 16895 1822 16904
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16250 1624 16526
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1872 16289 1900 16458
rect 1858 16280 1914 16289
rect 1584 16244 1636 16250
rect 1858 16215 1914 16224
rect 1584 16186 1636 16192
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1780 15609 1808 15982
rect 1766 15600 1822 15609
rect 1766 15535 1822 15544
rect 1768 14952 1820 14958
rect 1766 14920 1768 14929
rect 1820 14920 1822 14929
rect 1766 14855 1822 14864
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1872 14249 1900 14282
rect 1858 14240 1914 14249
rect 1858 14175 1914 14184
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13569 1808 13806
rect 1766 13560 1822 13569
rect 1766 13495 1822 13504
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1872 12889 1900 13194
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1860 12232 1912 12238
rect 1858 12200 1860 12209
rect 1912 12200 1914 12209
rect 1858 12135 1914 12144
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1780 11529 1808 11630
rect 1766 11520 1822 11529
rect 1766 11455 1822 11464
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10849 1900 11018
rect 1858 10840 1914 10849
rect 1858 10775 1914 10784
rect 1582 10704 1638 10713
rect 1582 10639 1584 10648
rect 1636 10639 1638 10648
rect 1584 10610 1636 10616
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1780 10169 1808 10542
rect 1964 10266 1992 35866
rect 2148 33590 2176 36790
rect 2240 36786 2268 37130
rect 2228 36780 2280 36786
rect 2228 36722 2280 36728
rect 2332 35766 2360 37130
rect 2516 36174 2544 59910
rect 2596 50856 2648 50862
rect 2596 50798 2648 50804
rect 2608 39302 2636 50798
rect 3344 47598 3372 60454
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 3884 60036 3936 60042
rect 3884 59978 3936 59984
rect 3896 50930 3924 59978
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 3976 51332 4028 51338
rect 3976 51274 4028 51280
rect 3988 50998 4016 51274
rect 4632 51066 4660 60522
rect 4816 51785 4844 60590
rect 5552 59634 5580 61066
rect 5724 61056 5776 61062
rect 5724 60998 5776 61004
rect 5540 59628 5592 59634
rect 5540 59570 5592 59576
rect 4802 51776 4858 51785
rect 4802 51711 4858 51720
rect 4620 51060 4672 51066
rect 4620 51002 4672 51008
rect 3976 50992 4028 50998
rect 3976 50934 4028 50940
rect 3884 50924 3936 50930
rect 3884 50866 3936 50872
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 3332 47592 3384 47598
rect 3332 47534 3384 47540
rect 5448 47524 5500 47530
rect 5448 47466 5500 47472
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 5460 42158 5488 47466
rect 5448 42152 5500 42158
rect 5448 42094 5500 42100
rect 5540 42084 5592 42090
rect 5540 42026 5592 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 5552 41002 5580 42026
rect 5632 42016 5684 42022
rect 5632 41958 5684 41964
rect 5540 40996 5592 41002
rect 5540 40938 5592 40944
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 2596 39296 2648 39302
rect 2596 39238 2648 39244
rect 2608 36854 2636 39238
rect 4804 38820 4856 38826
rect 4804 38762 4856 38768
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4816 37874 4844 38762
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4988 37868 5040 37874
rect 4988 37810 5040 37816
rect 4068 37732 4120 37738
rect 4068 37674 4120 37680
rect 2596 36848 2648 36854
rect 2596 36790 2648 36796
rect 2504 36168 2556 36174
rect 2504 36110 2556 36116
rect 2608 36106 2636 36790
rect 2688 36780 2740 36786
rect 2688 36722 2740 36728
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 2700 36242 2728 36722
rect 3068 36689 3096 36722
rect 3054 36680 3110 36689
rect 3054 36615 3110 36624
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 2688 36236 2740 36242
rect 2688 36178 2740 36184
rect 2596 36100 2648 36106
rect 2596 36042 2648 36048
rect 2320 35760 2372 35766
rect 2320 35702 2372 35708
rect 2136 33584 2188 33590
rect 2136 33526 2188 33532
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2516 26994 2544 28018
rect 2700 26994 2728 36178
rect 2780 36100 2832 36106
rect 2780 36042 2832 36048
rect 2792 35222 2820 36042
rect 2780 35216 2832 35222
rect 2780 35158 2832 35164
rect 3252 27402 3280 36518
rect 4080 30190 4108 37674
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5000 28082 5028 37810
rect 5644 36174 5672 41958
rect 5632 36168 5684 36174
rect 5632 36110 5684 36116
rect 5172 36032 5224 36038
rect 5172 35974 5224 35980
rect 4988 28076 5040 28082
rect 4988 28018 5040 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3240 27396 3292 27402
rect 3240 27338 3292 27344
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2688 26988 2740 26994
rect 2688 26930 2740 26936
rect 2516 25294 2544 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5184 25702 5212 35974
rect 5736 30326 5764 60998
rect 6288 60110 6316 61270
rect 6656 61198 6684 63294
rect 6734 63200 6790 63294
rect 7470 63322 7526 64000
rect 7470 63294 7604 63322
rect 7470 63200 7526 63294
rect 7576 61198 7604 63294
rect 8206 63200 8262 64000
rect 8942 63322 8998 64000
rect 9678 63322 9734 64000
rect 10414 63322 10470 64000
rect 8942 63294 9260 63322
rect 8942 63200 8998 63294
rect 7656 61396 7708 61402
rect 7656 61338 7708 61344
rect 6644 61192 6696 61198
rect 6644 61134 6696 61140
rect 7564 61192 7616 61198
rect 7564 61134 7616 61140
rect 6644 60240 6696 60246
rect 6644 60182 6696 60188
rect 6000 60104 6052 60110
rect 6000 60046 6052 60052
rect 6276 60104 6328 60110
rect 6276 60046 6328 60052
rect 6012 59158 6040 60046
rect 6000 59152 6052 59158
rect 6000 59094 6052 59100
rect 5908 50720 5960 50726
rect 5908 50662 5960 50668
rect 5920 36174 5948 50662
rect 6184 37256 6236 37262
rect 6184 37198 6236 37204
rect 6196 36174 6224 37198
rect 6656 36854 6684 60182
rect 7012 60104 7064 60110
rect 7012 60046 7064 60052
rect 6736 60036 6788 60042
rect 6736 59978 6788 59984
rect 6748 59702 6776 59978
rect 6736 59696 6788 59702
rect 6736 59638 6788 59644
rect 6826 59664 6882 59673
rect 7024 59634 7052 60046
rect 6826 59599 6828 59608
rect 6880 59599 6882 59608
rect 7012 59628 7064 59634
rect 6828 59570 6880 59576
rect 7012 59570 7064 59576
rect 6828 59424 6880 59430
rect 6828 59366 6880 59372
rect 6840 52018 6868 59366
rect 6828 52012 6880 52018
rect 6828 51954 6880 51960
rect 6736 51808 6788 51814
rect 6736 51750 6788 51756
rect 6748 43450 6776 51750
rect 6736 43444 6788 43450
rect 6736 43386 6788 43392
rect 6736 37664 6788 37670
rect 6736 37606 6788 37612
rect 6644 36848 6696 36854
rect 6644 36790 6696 36796
rect 6748 36718 6776 37606
rect 7024 36854 7052 59570
rect 7104 52012 7156 52018
rect 7104 51954 7156 51960
rect 7116 50930 7144 51954
rect 7104 50924 7156 50930
rect 7104 50866 7156 50872
rect 7564 50924 7616 50930
rect 7564 50866 7616 50872
rect 7576 45490 7604 50866
rect 7564 45484 7616 45490
rect 7564 45426 7616 45432
rect 7576 37194 7604 45426
rect 7564 37188 7616 37194
rect 7564 37130 7616 37136
rect 7012 36848 7064 36854
rect 7012 36790 7064 36796
rect 6736 36712 6788 36718
rect 6736 36654 6788 36660
rect 5908 36168 5960 36174
rect 5908 36110 5960 36116
rect 6184 36168 6236 36174
rect 6184 36110 6236 36116
rect 5724 30320 5776 30326
rect 5724 30262 5776 30268
rect 6196 26926 6224 36110
rect 7024 36106 7052 36790
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7208 36174 7236 36314
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 7012 36100 7064 36106
rect 7012 36042 7064 36048
rect 7668 28422 7696 61338
rect 7840 61124 7892 61130
rect 7840 61066 7892 61072
rect 7852 49162 7880 61066
rect 8220 60874 8248 63200
rect 9232 61198 9260 63294
rect 9678 63294 9904 63322
rect 9678 63200 9734 63294
rect 9220 61192 9272 61198
rect 9220 61134 9272 61140
rect 9312 61056 9364 61062
rect 9312 60998 9364 61004
rect 8220 60846 8340 60874
rect 8312 60790 8340 60846
rect 8300 60784 8352 60790
rect 8300 60726 8352 60732
rect 7840 49156 7892 49162
rect 7840 49098 7892 49104
rect 9324 39030 9352 60998
rect 9876 60790 9904 63294
rect 10244 63294 10470 63322
rect 10244 61198 10272 63294
rect 10414 63200 10470 63294
rect 11150 63200 11206 64000
rect 11886 63322 11942 64000
rect 12622 63322 12678 64000
rect 13358 63322 13414 64000
rect 14094 63322 14150 64000
rect 14830 63322 14886 64000
rect 15566 63322 15622 64000
rect 16302 63322 16358 64000
rect 11886 63294 12112 63322
rect 11886 63200 11942 63294
rect 11164 61198 11192 63200
rect 12084 61198 12112 63294
rect 12622 63294 12848 63322
rect 12622 63200 12678 63294
rect 12820 61198 12848 63294
rect 13358 63294 13584 63322
rect 13358 63200 13414 63294
rect 10232 61192 10284 61198
rect 10232 61134 10284 61140
rect 11152 61192 11204 61198
rect 11152 61134 11204 61140
rect 12072 61192 12124 61198
rect 12072 61134 12124 61140
rect 12808 61192 12860 61198
rect 12808 61134 12860 61140
rect 10508 61124 10560 61130
rect 10508 61066 10560 61072
rect 10324 61056 10376 61062
rect 10324 60998 10376 61004
rect 10336 60858 10364 60998
rect 10324 60852 10376 60858
rect 10324 60794 10376 60800
rect 9864 60784 9916 60790
rect 9864 60726 9916 60732
rect 9956 60512 10008 60518
rect 9956 60454 10008 60460
rect 9968 60314 9996 60454
rect 9956 60308 10008 60314
rect 9956 60250 10008 60256
rect 9312 39024 9364 39030
rect 9312 38966 9364 38972
rect 7840 36712 7892 36718
rect 7840 36654 7892 36660
rect 7852 36378 7880 36654
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15570 2452 15846
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2412 14952 2464 14958
rect 2410 14920 2412 14929
rect 2464 14920 2466 14929
rect 2410 14855 2466 14864
rect 2410 14376 2466 14385
rect 2410 14311 2466 14320
rect 2424 14074 2452 14311
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1766 10160 1822 10169
rect 1766 10095 1822 10104
rect 1582 9616 1638 9625
rect 1582 9551 1584 9560
rect 1636 9551 1638 9560
rect 1584 9522 1636 9528
rect 1768 9512 1820 9518
rect 1766 9480 1768 9489
rect 1820 9480 1822 9489
rect 1766 9415 1822 9424
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8809 1900 8842
rect 1858 8800 1914 8809
rect 1858 8735 1914 8744
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8129 1808 8366
rect 1766 8120 1822 8129
rect 1766 8055 1822 8064
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7449 1900 7754
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 1858 6760 1914 6769
rect 1858 6695 1860 6704
rect 1912 6695 1914 6704
rect 1860 6666 1912 6672
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1780 6089 1808 6190
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5409 1900 5578
rect 1858 5400 1914 5409
rect 1858 5335 1914 5344
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4729 1808 5102
rect 1766 4720 1822 4729
rect 1766 4655 1822 4664
rect 1768 4072 1820 4078
rect 1766 4040 1768 4049
rect 1820 4040 1822 4049
rect 1766 3975 1822 3984
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1872 3369 1900 3402
rect 1858 3360 1914 3369
rect 1858 3295 1914 3304
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2689 1808 2926
rect 1766 2680 1822 2689
rect 1766 2615 1822 2624
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1596 1562 1624 2382
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 2009 1900 2314
rect 1858 2000 1914 2009
rect 1858 1935 1914 1944
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 2332 678 2360 13126
rect 2516 8566 2544 25230
rect 2700 24750 2728 25230
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 6932 24206 6960 24278
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 3146 5128 3202 5137
rect 3146 5063 3202 5072
rect 3160 4146 3188 5063
rect 3712 4146 3740 17206
rect 4080 16046 4108 19790
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 7576 18426 7604 19110
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 8220 14958 8248 21490
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 7576 11150 7604 11834
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7576 10266 7604 10746
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2884 3058 2912 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3160 882 3188 3470
rect 4172 3194 4200 3606
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 1426 3372 2246
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3620 1154 3648 2994
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3608 1148 3660 1154
rect 3608 1090 3660 1096
rect 3712 921 3740 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2122 4660 4150
rect 5092 3670 5120 6122
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4172 2094 4660 2122
rect 3698 912 3754 921
rect 3148 876 3200 882
rect 3698 847 3754 856
rect 3148 818 3200 824
rect 4172 800 4200 2094
rect 4724 1494 4752 2994
rect 4712 1488 4764 1494
rect 4712 1430 4764 1436
rect 2320 672 2372 678
rect 2320 614 2372 620
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4816 746 4844 3062
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 4908 1766 4936 2314
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 5000 1086 5028 3470
rect 5170 3224 5226 3233
rect 5170 3159 5226 3168
rect 5184 2854 5212 3159
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 5092 1970 5120 2314
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 5184 1630 5212 2246
rect 5172 1624 5224 1630
rect 5172 1566 5224 1572
rect 4988 1080 5040 1086
rect 4988 1022 5040 1028
rect 5368 950 5396 3946
rect 5552 3942 5580 5782
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5644 2122 5672 4218
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5552 2094 5672 2122
rect 5356 944 5408 950
rect 5356 886 5408 892
rect 5552 800 5580 2094
rect 5736 1714 5764 3674
rect 5828 2854 5856 9386
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 4758 7052 7278
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5828 2038 5856 2314
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 5920 1714 5948 3334
rect 6012 1850 6040 3538
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 2922 6132 3334
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 6012 1822 6224 1850
rect 5736 1686 5856 1714
rect 5920 1686 6132 1714
rect 5828 800 5856 1686
rect 6104 800 6132 1686
rect 6196 814 6224 1822
rect 6184 808 6236 814
rect 4804 740 4856 746
rect 4804 682 4856 688
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6090 0 6146 800
rect 6380 800 6408 4150
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6472 1018 6500 3946
rect 6564 3194 6592 3946
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6460 1012 6512 1018
rect 6460 954 6512 960
rect 6656 800 6684 4490
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6748 2961 6776 3402
rect 6734 2952 6790 2961
rect 6734 2887 6790 2896
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 1834 6776 2314
rect 6736 1828 6788 1834
rect 6736 1770 6788 1776
rect 6932 800 6960 4082
rect 7024 3602 7052 4218
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3738 7236 3878
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7300 3126 7328 3538
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7392 2774 7420 3470
rect 7576 3398 7604 5034
rect 7564 3392 7616 3398
rect 7470 3360 7526 3369
rect 7564 3334 7616 3340
rect 7470 3295 7526 3304
rect 7484 3126 7512 3295
rect 7668 3210 7696 10134
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7576 3182 7696 3210
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7392 2746 7512 2774
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 7024 1902 7052 2314
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 7196 1148 7248 1154
rect 7196 1090 7248 1096
rect 7208 800 7236 1090
rect 7484 800 7512 2746
rect 7576 2582 7604 3182
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7760 800 7788 4150
rect 7852 2582 7880 13738
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 7478 8708 8502
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 4078 7972 4150
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8036 800 8064 4490
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8128 3466 8156 4150
rect 8404 4078 8432 5170
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8128 3126 8156 3402
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8128 2378 8156 3062
rect 8496 2582 8524 4966
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8300 1488 8352 1494
rect 8300 1430 8352 1436
rect 8312 800 8340 1430
rect 8588 800 8616 5170
rect 8666 4856 8722 4865
rect 8666 4791 8722 4800
rect 8680 4758 8708 4791
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 3670 8708 4490
rect 8864 4146 8892 7142
rect 8956 6254 8984 14350
rect 9600 7546 9628 27338
rect 10520 26897 10548 61066
rect 12164 61056 12216 61062
rect 12164 60998 12216 61004
rect 12900 61056 12952 61062
rect 12900 60998 12952 61004
rect 10968 53984 11020 53990
rect 10968 53926 11020 53932
rect 10980 53650 11008 53926
rect 10968 53644 11020 53650
rect 10968 53586 11020 53592
rect 11060 40384 11112 40390
rect 11060 40326 11112 40332
rect 11072 38282 11100 40326
rect 11060 38276 11112 38282
rect 11060 38218 11112 38224
rect 12176 35018 12204 60998
rect 12912 60761 12940 60998
rect 13556 60790 13584 63294
rect 14094 63294 14320 63322
rect 14094 63200 14150 63294
rect 14292 60790 14320 63294
rect 14830 63294 14964 63322
rect 14830 63200 14886 63294
rect 14936 61198 14964 63294
rect 15566 63294 15792 63322
rect 15566 63200 15622 63294
rect 15292 61396 15344 61402
rect 15292 61338 15344 61344
rect 14924 61192 14976 61198
rect 14924 61134 14976 61140
rect 15200 61124 15252 61130
rect 15200 61066 15252 61072
rect 13544 60784 13596 60790
rect 12898 60752 12954 60761
rect 13544 60726 13596 60732
rect 14280 60784 14332 60790
rect 14280 60726 14332 60732
rect 12898 60687 12954 60696
rect 13636 60648 13688 60654
rect 13636 60590 13688 60596
rect 13648 60246 13676 60590
rect 13636 60240 13688 60246
rect 13636 60182 13688 60188
rect 15212 50289 15240 61066
rect 15304 59702 15332 61338
rect 15764 60790 15792 63294
rect 16132 63294 16358 63322
rect 16132 61198 16160 63294
rect 16302 63200 16358 63294
rect 17038 63322 17094 64000
rect 17774 63322 17830 64000
rect 18510 63322 18566 64000
rect 17038 63294 17172 63322
rect 17038 63200 17094 63294
rect 17144 61198 17172 63294
rect 17774 63294 17908 63322
rect 17774 63200 17830 63294
rect 17408 61260 17460 61266
rect 17408 61202 17460 61208
rect 16120 61192 16172 61198
rect 16120 61134 16172 61140
rect 17132 61192 17184 61198
rect 17132 61134 17184 61140
rect 17316 61056 17368 61062
rect 17316 60998 17368 61004
rect 15752 60784 15804 60790
rect 15752 60726 15804 60732
rect 15844 60512 15896 60518
rect 15844 60454 15896 60460
rect 15856 60178 15884 60454
rect 15844 60172 15896 60178
rect 15844 60114 15896 60120
rect 15292 59696 15344 59702
rect 15292 59638 15344 59644
rect 17224 57860 17276 57866
rect 17224 57802 17276 57808
rect 15198 50280 15254 50289
rect 15198 50215 15254 50224
rect 15844 49088 15896 49094
rect 15844 49030 15896 49036
rect 15856 40118 15884 49030
rect 17132 44192 17184 44198
rect 17132 44134 17184 44140
rect 17144 43858 17172 44134
rect 17132 43852 17184 43858
rect 17132 43794 17184 43800
rect 15844 40112 15896 40118
rect 15844 40054 15896 40060
rect 15844 39568 15896 39574
rect 15844 39510 15896 39516
rect 15856 35494 15884 39510
rect 16396 37120 16448 37126
rect 16396 37062 16448 37068
rect 16408 36378 16436 37062
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16396 36372 16448 36378
rect 16396 36314 16448 36320
rect 15844 35488 15896 35494
rect 15844 35430 15896 35436
rect 16684 35222 16712 36518
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 12164 35012 12216 35018
rect 12164 34954 12216 34960
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 14464 27940 14516 27946
rect 14464 27882 14516 27888
rect 10506 26888 10562 26897
rect 10506 26823 10562 26832
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10230 13832 10286 13841
rect 10230 13767 10286 13776
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 12850 10088 13670
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 12442 10088 12786
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 7313 9444 7346
rect 9692 7342 9720 7754
rect 10152 7342 10180 7822
rect 9680 7336 9732 7342
rect 9402 7304 9458 7313
rect 9680 7278 9732 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9402 7239 9458 7248
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 4026 8892 4082
rect 8772 3998 8892 4026
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 1154 8708 3334
rect 8772 2553 8800 3998
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8864 800 8892 3402
rect 8956 2009 8984 4014
rect 9048 3194 9076 5170
rect 9232 4826 9260 5646
rect 9310 4992 9366 5001
rect 9310 4927 9366 4936
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9324 4554 9352 4927
rect 9416 4826 9444 7239
rect 9692 6390 9720 7278
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 5370 9628 6258
rect 9876 5370 9904 6734
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 5098 10088 5170
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9586 4856 9642 4865
rect 9404 4820 9456 4826
rect 10152 4826 10180 6734
rect 9586 4791 9588 4800
rect 9404 4762 9456 4768
rect 9640 4791 9642 4800
rect 10140 4820 10192 4826
rect 9588 4762 9640 4768
rect 10140 4762 10192 4768
rect 9600 4690 9812 4706
rect 9588 4684 9824 4690
rect 9640 4678 9772 4684
rect 9588 4626 9640 4632
rect 9772 4626 9824 4632
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9140 4185 9168 4422
rect 9218 4312 9274 4321
rect 9218 4247 9274 4256
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8942 2000 8998 2009
rect 8942 1935 8998 1944
rect 9140 800 9168 3606
rect 9232 3058 9260 4247
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9324 2106 9352 2382
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9416 800 9444 3878
rect 9508 3369 9536 4422
rect 9600 4146 9628 4626
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9494 3360 9550 3369
rect 9494 3295 9550 3304
rect 9588 2644 9640 2650
rect 9692 2632 9720 4558
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9862 2952 9918 2961
rect 9862 2887 9864 2896
rect 9916 2887 9918 2896
rect 9864 2858 9916 2864
rect 9640 2604 9720 2632
rect 9588 2586 9640 2592
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 800 9720 2314
rect 9968 800 9996 3470
rect 10244 3058 10272 13767
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10336 7857 10364 8366
rect 10322 7848 10378 7857
rect 10322 7783 10378 7792
rect 10336 7410 10364 7783
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5166 10364 6054
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10336 4690 10364 5102
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10336 3670 10364 4626
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10428 3534 10456 14826
rect 10796 14414 10824 18022
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11072 16454 11100 17614
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10980 14278 11008 14758
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10612 12889 10640 13262
rect 10598 12880 10654 12889
rect 10598 12815 10654 12824
rect 10704 12782 10732 13942
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10704 12374 10732 12718
rect 10692 12368 10744 12374
rect 10796 12345 10824 13262
rect 11072 13190 11100 14010
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11164 12986 11192 16118
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11242 15056 11298 15065
rect 11242 14991 11244 15000
rect 11296 14991 11298 15000
rect 11244 14962 11296 14968
rect 11440 14618 11468 15438
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11624 14414 11652 17478
rect 13740 17270 13768 18090
rect 14200 17678 14228 18226
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 11794 14784 11850 14793
rect 11794 14719 11850 14728
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13569 11468 13806
rect 11426 13560 11482 13569
rect 11426 13495 11482 13504
rect 11440 13326 11468 13495
rect 11624 13394 11652 14350
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11808 12730 11836 14719
rect 12176 14006 12204 15914
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12850 11928 13262
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12753 11928 12786
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11716 12702 11836 12730
rect 11886 12744 11942 12753
rect 10692 12310 10744 12316
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10690 11928 10746 11937
rect 10690 11863 10746 11872
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10520 7818 10548 8366
rect 10612 8090 10640 8366
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10520 7342 10548 7754
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10520 7002 10548 7278
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10520 6730 10548 6938
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10612 6458 10640 7278
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10152 1816 10180 2926
rect 10152 1788 10272 1816
rect 10244 800 10272 1788
rect 10520 800 10548 5578
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10612 4593 10640 5238
rect 10598 4584 10654 4593
rect 10598 4519 10654 4528
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 1494 10640 3878
rect 10704 3058 10732 11863
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10704 1222 10732 2382
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10796 800 10824 5170
rect 10888 2582 10916 9318
rect 10980 5914 11008 12650
rect 11716 12306 11744 12702
rect 11886 12679 11942 12688
rect 11992 12374 12020 13806
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11702 12200 11758 12209
rect 11624 11762 11652 12174
rect 11702 12135 11758 12144
rect 11716 11830 11744 12135
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 11393 11652 11698
rect 11808 11626 11836 12242
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11610 11384 11666 11393
rect 11610 11319 11666 11328
rect 11808 10130 11836 11562
rect 11900 10266 11928 12174
rect 12084 11150 12112 13806
rect 12268 11898 12296 13874
rect 12360 13297 12388 16458
rect 13188 16250 13216 16526
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13188 16114 13216 16186
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 14074 12480 15982
rect 13280 15978 13308 16050
rect 13556 16046 13584 16526
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14618 13492 14758
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13266 14240 13322 14249
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 13096 14006 13124 14214
rect 13266 14175 13322 14184
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12532 13864 12584 13870
rect 12452 13824 12532 13852
rect 12346 13288 12402 13297
rect 12346 13223 12402 13232
rect 12360 13190 12388 13223
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12452 12850 12480 13824
rect 12532 13806 12584 13812
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 13716 12664 13806
rect 12544 13688 12664 13716
rect 12900 13728 12952 13734
rect 12544 12866 12572 13688
rect 12900 13670 12952 13676
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12622 13016 12678 13025
rect 12622 12951 12624 12960
rect 12676 12951 12678 12960
rect 12624 12922 12676 12928
rect 12716 12912 12768 12918
rect 12544 12860 12716 12866
rect 12544 12854 12768 12860
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12544 12838 12756 12854
rect 12438 12744 12494 12753
rect 12348 12708 12400 12714
rect 12438 12679 12494 12688
rect 12348 12650 12400 12656
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9674 11836 10066
rect 11808 9646 12020 9674
rect 11992 9586 12020 9646
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11072 4010 11100 6122
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 1630 11008 2314
rect 10968 1624 11020 1630
rect 10968 1566 11020 1572
rect 11072 800 11100 2790
rect 11164 1426 11192 7958
rect 11256 5302 11284 8366
rect 11886 8256 11942 8265
rect 11886 8191 11942 8200
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11348 5166 11376 6734
rect 11716 6322 11744 6734
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11348 4690 11376 5102
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11336 1760 11388 1766
rect 11336 1702 11388 1708
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11348 800 11376 1702
rect 11440 1698 11468 5034
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3233 11560 3606
rect 11518 3224 11574 3233
rect 11518 3159 11574 3168
rect 11428 1692 11480 1698
rect 11428 1634 11480 1640
rect 11624 800 11652 6258
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 4758 11744 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11808 2417 11836 5170
rect 11900 3670 11928 8191
rect 11992 5302 12020 9522
rect 12176 9518 12204 11630
rect 12268 11218 12296 11834
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12360 10198 12388 12650
rect 12452 12170 12480 12679
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12544 10130 12572 12838
rect 12820 12730 12848 13398
rect 12912 13326 12940 13670
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12636 12702 12848 12730
rect 12636 12170 12664 12702
rect 12912 12442 12940 13262
rect 12992 13184 13044 13190
rect 12990 13152 12992 13161
rect 13176 13184 13228 13190
rect 13044 13152 13046 13161
rect 13176 13126 13228 13132
rect 12990 13087 13046 13096
rect 13188 12986 13216 13126
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13280 12866 13308 14175
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13705 13584 13874
rect 13542 13696 13598 13705
rect 13542 13631 13598 13640
rect 13556 13394 13584 13631
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13542 13152 13598 13161
rect 13542 13087 13598 13096
rect 13556 12918 13584 13087
rect 13188 12838 13308 12866
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12806 12064 12862 12073
rect 12806 11999 12862 12008
rect 12820 11558 12848 11999
rect 12900 11756 12952 11762
rect 13004 11744 13032 12106
rect 12952 11716 13032 11744
rect 12900 11698 12952 11704
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10849 12664 11086
rect 12622 10840 12678 10849
rect 12622 10775 12678 10784
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 8430 12112 9386
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 12162 5264 12218 5273
rect 11992 4214 12020 5238
rect 12162 5199 12218 5208
rect 12176 5030 12204 5199
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 12084 3233 12112 4694
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4554 12204 4626
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12176 4146 12204 4490
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12070 3224 12126 3233
rect 12070 3159 12126 3168
rect 12176 3058 12204 3402
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 12084 2689 12112 2858
rect 12268 2774 12296 5578
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12360 4486 12388 4762
rect 12544 4758 12572 5578
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12530 3904 12586 3913
rect 12452 3505 12480 3878
rect 12530 3839 12586 3848
rect 12438 3496 12494 3505
rect 12438 3431 12494 3440
rect 12544 3058 12572 3839
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12636 2774 12664 5510
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12176 2746 12296 2774
rect 12452 2746 12664 2774
rect 12070 2680 12126 2689
rect 12070 2615 12126 2624
rect 11794 2408 11850 2417
rect 11794 2343 11850 2352
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11900 800 11928 1906
rect 12176 800 12204 2746
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12360 1970 12388 2382
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12452 800 12480 2746
rect 12622 2680 12678 2689
rect 12728 2650 12756 3946
rect 12622 2615 12678 2624
rect 12716 2644 12768 2650
rect 12636 1408 12664 2615
rect 12716 2586 12768 2592
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12728 1766 12756 2450
rect 12820 1902 12848 11290
rect 13004 7886 13032 11716
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12992 7880 13044 7886
rect 13096 7857 13124 10610
rect 12992 7822 13044 7828
rect 13082 7848 13138 7857
rect 13082 7783 13138 7792
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12912 4282 12940 4694
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12990 4176 13046 4185
rect 12990 4111 13046 4120
rect 13004 3942 13032 4111
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12808 1896 12860 1902
rect 12808 1838 12860 1844
rect 12716 1760 12768 1766
rect 13096 1714 13124 5578
rect 13188 3534 13216 12838
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13358 11248 13414 11257
rect 13358 11183 13414 11192
rect 13266 11112 13322 11121
rect 13266 11047 13322 11056
rect 13280 5216 13308 11047
rect 13372 10742 13400 11183
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13464 6730 13492 12174
rect 13556 11218 13584 12718
rect 13648 11354 13676 16526
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13802 13768 14350
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12714 13768 12786
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13832 12646 13860 17138
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 15026 13952 15438
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13924 14482 13952 14962
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13924 13394 13952 13738
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12646 13952 13126
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 14016 12442 14044 14962
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 13190 14136 13262
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14200 12782 14228 17614
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11762 13860 12038
rect 14186 11792 14242 11801
rect 13820 11756 13872 11762
rect 14186 11727 14242 11736
rect 13820 11698 13872 11704
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13832 10062 13860 11698
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 10742 13952 11630
rect 14200 11626 14228 11727
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13634 9072 13690 9081
rect 13634 9007 13690 9016
rect 13648 8498 13676 9007
rect 13740 8974 13768 9930
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13924 8838 13952 10678
rect 14108 9926 14136 10678
rect 14292 10674 14320 20402
rect 14476 18057 14504 27882
rect 15200 26852 15252 26858
rect 15200 26794 15252 26800
rect 15212 23594 15240 26794
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 14462 18048 14518 18057
rect 14462 17983 14518 17992
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14844 16658 14872 17546
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15502 14596 15846
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14464 13728 14516 13734
rect 14370 13696 14426 13705
rect 14464 13670 14516 13676
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14370 13631 14426 13640
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14384 9654 14412 13631
rect 14476 13394 14504 13670
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14556 13320 14608 13326
rect 14660 13274 14688 13670
rect 14608 13268 14688 13274
rect 14556 13262 14688 13268
rect 14568 13246 14688 13262
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12442 14596 12718
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14568 12306 14596 12378
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10985 14596 11154
rect 14554 10976 14610 10985
rect 14554 10911 14610 10920
rect 14660 10062 14688 13246
rect 14752 13025 14780 13806
rect 14844 13190 14872 16594
rect 14936 15473 14964 16934
rect 14922 15464 14978 15473
rect 14922 15399 14978 15408
rect 15028 15065 15056 19790
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 17338 15240 17614
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15014 15056 15070 15065
rect 15014 14991 15070 15000
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14738 13016 14794 13025
rect 14738 12951 14794 12960
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14752 12646 14780 12854
rect 14844 12753 14872 13126
rect 14830 12744 14886 12753
rect 14830 12679 14886 12688
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14752 12306 14780 12582
rect 14844 12306 14872 12582
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14752 11354 14780 11766
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10198 14780 10950
rect 14844 10810 14872 11018
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14462 9344 14518 9353
rect 14462 9279 14518 9288
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13740 8378 13768 8774
rect 13648 8350 13768 8378
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13280 5188 13492 5216
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13372 2774 13400 4966
rect 13464 3466 13492 5188
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13556 4214 13584 4490
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13648 3534 13676 8350
rect 13726 7712 13782 7721
rect 13726 7647 13782 7656
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13740 3058 13768 7647
rect 13910 7168 13966 7177
rect 13910 7103 13966 7112
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13372 2746 13492 2774
rect 13266 2680 13322 2689
rect 13266 2615 13322 2624
rect 13280 2446 13308 2615
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 12716 1702 12768 1708
rect 13004 1686 13124 1714
rect 12636 1380 12756 1408
rect 12728 800 12756 1380
rect 13004 800 13032 1686
rect 13280 800 13308 1974
rect 13372 1426 13400 2314
rect 13360 1420 13412 1426
rect 13360 1362 13412 1368
rect 13464 1290 13492 2746
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13556 1970 13584 2314
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13452 1284 13504 1290
rect 13452 1226 13504 1232
rect 13556 800 13584 1770
rect 13832 800 13860 5170
rect 13924 3058 13952 7103
rect 14002 7032 14058 7041
rect 14002 6967 14058 6976
rect 14016 4146 14044 6967
rect 14094 5264 14150 5273
rect 14094 5199 14096 5208
rect 14148 5199 14150 5208
rect 14096 5170 14148 5176
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14108 800 14136 3674
rect 14476 3534 14504 9279
rect 14568 6934 14596 9522
rect 14844 9178 14872 10610
rect 14936 9382 14964 13330
rect 15028 13326 15056 14991
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15120 12782 15148 16050
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 14482 15240 15846
rect 15396 14890 15424 16934
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15106 12336 15162 12345
rect 15106 12271 15162 12280
rect 15120 12238 15148 12271
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15028 11937 15056 12174
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15014 11928 15070 11937
rect 15014 11863 15070 11872
rect 15028 11830 15056 11863
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15212 11778 15240 12106
rect 15304 11898 15332 13874
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12481 15516 13262
rect 15474 12472 15530 12481
rect 15474 12407 15530 12416
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15212 11750 15332 11778
rect 15198 11656 15254 11665
rect 15198 11591 15254 11600
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 15028 9110 15056 10746
rect 15120 10169 15148 11494
rect 15212 10674 15240 11591
rect 15304 11150 15332 11750
rect 15396 11694 15424 12242
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15488 11762 15516 12106
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15580 11626 15608 14758
rect 15672 13326 15700 32370
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15764 17542 15792 18226
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15658 13016 15714 13025
rect 15764 12986 15792 17478
rect 15948 16590 15976 18770
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 16040 15162 16068 17750
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15844 14272 15896 14278
rect 15842 14240 15844 14249
rect 15896 14240 15898 14249
rect 15842 14175 15898 14184
rect 15948 14074 15976 14418
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15658 12951 15660 12960
rect 15712 12951 15714 12960
rect 15752 12980 15804 12986
rect 15660 12922 15712 12928
rect 15752 12922 15804 12928
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15658 12608 15714 12617
rect 15658 12543 15714 12552
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10810 15424 11018
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15106 10160 15162 10169
rect 15106 10095 15162 10104
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 15212 8634 15240 10406
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 14738 7712 14794 7721
rect 14738 7647 14794 7656
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14292 2825 14320 2926
rect 14568 2854 14596 3334
rect 14556 2848 14608 2854
rect 14278 2816 14334 2825
rect 14556 2790 14608 2796
rect 14278 2751 14334 2760
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14384 800 14412 2246
rect 14568 1465 14596 2518
rect 14554 1456 14610 1465
rect 14554 1391 14610 1400
rect 14660 800 14688 5578
rect 14752 3058 14780 7647
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14844 2774 14872 6598
rect 14922 6488 14978 6497
rect 15304 6458 15332 10610
rect 15488 10130 15516 10746
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15672 7562 15700 12543
rect 15750 12336 15806 12345
rect 15750 12271 15806 12280
rect 15764 10826 15792 12271
rect 15856 12102 15884 12650
rect 15948 12306 15976 14010
rect 16040 13802 16068 14214
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16028 13456 16080 13462
rect 16026 13424 16028 13433
rect 16080 13424 16082 13433
rect 16026 13359 16082 13368
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 11529 15976 11698
rect 15934 11520 15990 11529
rect 15934 11455 15990 11464
rect 15764 10798 15884 10826
rect 15856 10674 15884 10798
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15764 10577 15792 10610
rect 15750 10568 15806 10577
rect 15750 10503 15806 10512
rect 15856 9761 15884 10610
rect 16040 10266 16068 13194
rect 16132 12345 16160 22034
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 13938 16252 16594
rect 16408 15570 16436 29582
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16868 23730 16896 24074
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 17678 16620 20198
rect 16684 18766 16712 20810
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16684 17882 16712 18702
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16776 17785 16804 18702
rect 16762 17776 16818 17785
rect 16762 17711 16818 17720
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16592 15502 16620 17478
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16210 13696 16266 13705
rect 16210 13631 16266 13640
rect 16224 13530 16252 13631
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16118 12336 16174 12345
rect 16118 12271 16174 12280
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 10962 16160 12038
rect 16224 11150 16252 13262
rect 16316 12306 16344 15370
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16304 12300 16356 12306
rect 16356 12260 16436 12288
rect 16304 12242 16356 12248
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 11762 16344 12106
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16316 11506 16344 11698
rect 16408 11626 16436 12260
rect 16500 12238 16528 13874
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16316 11478 16436 11506
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16132 10934 16252 10962
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16132 10266 16160 10610
rect 16224 10606 16252 10934
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 15842 9752 15898 9761
rect 15842 9687 15898 9696
rect 16040 9602 16068 9930
rect 16132 9897 16160 9998
rect 16118 9888 16174 9897
rect 16118 9823 16174 9832
rect 15948 9574 16068 9602
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15856 9110 15884 9454
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15764 8022 15792 8774
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15580 7534 15700 7562
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 14922 6423 14978 6432
rect 15292 6452 15344 6458
rect 14936 4146 14964 6423
rect 15292 6394 15344 6400
rect 15488 5681 15516 7142
rect 15474 5672 15530 5681
rect 15474 5607 15530 5616
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 15290 3632 15346 3641
rect 14752 2746 14872 2774
rect 14752 2650 14780 2746
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14752 2446 14780 2586
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14936 800 14964 3606
rect 15290 3567 15346 3576
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 2582 15056 2790
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15120 1057 15148 1498
rect 15106 1048 15162 1057
rect 15106 983 15162 992
rect 15212 800 15240 2994
rect 15304 2990 15332 3567
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15396 2854 15424 4014
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15488 800 15516 2858
rect 15580 2038 15608 7534
rect 15658 7440 15714 7449
rect 15658 7375 15714 7384
rect 15672 4622 15700 7375
rect 15856 6322 15884 9046
rect 15948 7290 15976 9574
rect 16224 9364 16252 10406
rect 16316 9518 16344 11154
rect 16408 9586 16436 11478
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16224 9336 16344 9364
rect 16210 8936 16266 8945
rect 16210 8871 16212 8880
rect 16264 8871 16266 8880
rect 16212 8842 16264 8848
rect 16316 8809 16344 9336
rect 16408 8974 16436 9386
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16396 8832 16448 8838
rect 16302 8800 16358 8809
rect 16396 8774 16448 8780
rect 16302 8735 16358 8744
rect 16408 8634 16436 8774
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 15948 7262 16252 7290
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15856 5302 15884 6258
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15856 4554 15884 5238
rect 16132 5098 16160 5714
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 4196 15884 4490
rect 15936 4208 15988 4214
rect 15856 4168 15936 4196
rect 15936 4150 15988 4156
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 15672 1193 15700 4082
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15658 1184 15714 1193
rect 15658 1119 15714 1128
rect 15764 800 15792 3538
rect 16224 3466 16252 7262
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 15856 2961 15884 3402
rect 15842 2952 15898 2961
rect 15842 2887 15898 2896
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15856 1562 15884 2382
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15948 1834 15976 2314
rect 15936 1828 15988 1834
rect 15936 1770 15988 1776
rect 15844 1556 15896 1562
rect 15844 1498 15896 1504
rect 16040 800 16068 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 1698 16160 2314
rect 16120 1692 16172 1698
rect 16120 1634 16172 1640
rect 16316 800 16344 6054
rect 16408 2446 16436 6734
rect 16500 5914 16528 9930
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 2774 16528 5646
rect 16592 4622 16620 11698
rect 16684 11121 16712 16934
rect 16776 16726 16804 17478
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16868 16046 16896 17070
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16868 14958 16896 15982
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 14482 16896 14894
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 13938 16896 14418
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12850 16896 13262
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16868 12073 16896 12174
rect 16854 12064 16910 12073
rect 16854 11999 16910 12008
rect 16960 11762 16988 32914
rect 17236 24313 17264 57802
rect 17328 51814 17356 60998
rect 17316 51808 17368 51814
rect 17316 51750 17368 51756
rect 17222 24304 17278 24313
rect 17222 24239 17278 24248
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17236 23866 17264 24142
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17328 18766 17356 19722
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17144 17921 17172 18362
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17130 17912 17186 17921
rect 17130 17847 17186 17856
rect 17236 17678 17264 18158
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17134 17264 17614
rect 17420 17241 17448 61202
rect 17880 61180 17908 63294
rect 18510 63294 18736 63322
rect 18510 63200 18566 63294
rect 18708 61198 18736 63294
rect 19246 63200 19302 64000
rect 19982 63322 20038 64000
rect 19812 63294 20038 63322
rect 17960 61192 18012 61198
rect 17880 61152 17960 61180
rect 17960 61134 18012 61140
rect 18696 61192 18748 61198
rect 18696 61134 18748 61140
rect 17500 61124 17552 61130
rect 17500 61066 17552 61072
rect 17512 48226 17540 61066
rect 18604 61056 18656 61062
rect 18604 60998 18656 61004
rect 17684 59968 17736 59974
rect 17684 59910 17736 59916
rect 17696 50425 17724 59910
rect 18512 59424 18564 59430
rect 18510 59392 18512 59401
rect 18564 59392 18566 59401
rect 18510 59327 18566 59336
rect 18052 54732 18104 54738
rect 18052 54674 18104 54680
rect 17682 50416 17738 50425
rect 17682 50351 17738 50360
rect 17512 48198 17908 48226
rect 17684 45824 17736 45830
rect 17684 45766 17736 45772
rect 17696 45490 17724 45766
rect 17880 45626 17908 48198
rect 17868 45620 17920 45626
rect 17868 45562 17920 45568
rect 17776 45552 17828 45558
rect 17776 45494 17828 45500
rect 17684 45484 17736 45490
rect 17684 45426 17736 45432
rect 17788 45082 17816 45494
rect 17776 45076 17828 45082
rect 17776 45018 17828 45024
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 17972 36689 18000 36722
rect 18064 36718 18092 54674
rect 18236 45484 18288 45490
rect 18236 45426 18288 45432
rect 18248 45370 18276 45426
rect 18248 45342 18368 45370
rect 18340 45286 18368 45342
rect 18236 45280 18288 45286
rect 18236 45222 18288 45228
rect 18328 45280 18380 45286
rect 18328 45222 18380 45228
rect 18052 36712 18104 36718
rect 17958 36680 18014 36689
rect 18052 36654 18104 36660
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 17958 36615 18014 36624
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 17972 29238 18000 30194
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17696 25906 17724 29106
rect 18064 26994 18092 36654
rect 18156 32774 18184 36654
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 18248 31278 18276 45222
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17696 23662 17724 25842
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17696 23118 17724 23598
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17696 22574 17724 23054
rect 17684 22568 17736 22574
rect 17684 22510 17736 22516
rect 17696 22030 17724 22510
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17590 19136 17646 19145
rect 17590 19071 17646 19080
rect 17604 18834 17632 19071
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17406 17232 17462 17241
rect 17406 17167 17462 17176
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17052 12782 17080 15098
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16946 11384 17002 11393
rect 16764 11348 16816 11354
rect 16946 11319 17002 11328
rect 16764 11290 16816 11296
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 8430 16712 9862
rect 16776 9382 16804 11290
rect 16960 10674 16988 11319
rect 17052 11257 17080 11834
rect 17038 11248 17094 11257
rect 17038 11183 17094 11192
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16868 10305 16896 10610
rect 17052 10606 17080 10950
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16854 10296 16910 10305
rect 16854 10231 16910 10240
rect 16946 10160 17002 10169
rect 16946 10095 17002 10104
rect 16960 10062 16988 10095
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9722 16988 9998
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 17144 9586 17172 14214
rect 17236 14074 17264 14894
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17328 12850 17356 15574
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17420 13569 17448 14010
rect 17406 13560 17462 13569
rect 17406 13495 17462 13504
rect 17512 13326 17540 18362
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12918 17448 13194
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17498 12880 17554 12889
rect 17316 12844 17368 12850
rect 17498 12815 17554 12824
rect 17316 12786 17368 12792
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17236 11898 17264 12242
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 11257 17356 11630
rect 17314 11248 17370 11257
rect 17314 11183 17370 11192
rect 17420 11121 17448 11698
rect 17512 11694 17540 12815
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17512 11354 17540 11630
rect 17590 11520 17646 11529
rect 17590 11455 17646 11464
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17406 11112 17462 11121
rect 17224 11076 17276 11082
rect 17406 11047 17462 11056
rect 17224 11018 17276 11024
rect 17236 10985 17264 11018
rect 17222 10976 17278 10985
rect 17222 10911 17278 10920
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17236 9654 17264 9998
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16946 9480 17002 9489
rect 16946 9415 17002 9424
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 9178 16896 9318
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 8090 16712 8366
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7886 16712 8026
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16776 5166 16804 8298
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16776 3670 16804 4490
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16776 3126 16804 3402
rect 16580 3120 16632 3126
rect 16578 3088 16580 3097
rect 16764 3120 16816 3126
rect 16632 3088 16634 3097
rect 16764 3062 16816 3068
rect 16578 3023 16634 3032
rect 16500 2746 16620 2774
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 16592 800 16620 2746
rect 16868 800 16896 5646
rect 16960 5234 16988 9415
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 7954 17172 8434
rect 17236 7954 17264 9590
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 7342 17172 7686
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 6769 17264 6802
rect 17222 6760 17278 6769
rect 17222 6695 17278 6704
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17144 5846 17172 6122
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17328 5778 17356 10406
rect 17420 9353 17448 11047
rect 17604 10470 17632 11455
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17498 10160 17554 10169
rect 17498 10095 17554 10104
rect 17406 9344 17462 9353
rect 17406 9279 17462 9288
rect 17406 9208 17462 9217
rect 17406 9143 17408 9152
rect 17460 9143 17462 9152
rect 17408 9114 17460 9120
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17420 8566 17448 8842
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17512 6662 17540 10095
rect 17696 9994 17724 21966
rect 18052 19848 18104 19854
rect 18050 19816 18052 19825
rect 18104 19816 18106 19825
rect 18050 19751 18106 19760
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17880 18358 17908 18770
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 18064 16590 18092 19654
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 15706 17816 16050
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15706 17908 15846
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17788 10130 17816 15506
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17866 13968 17922 13977
rect 17866 13903 17922 13912
rect 17880 11626 17908 13903
rect 17972 13326 18000 14962
rect 18050 13832 18106 13841
rect 18050 13767 18052 13776
rect 18104 13767 18106 13776
rect 18052 13738 18104 13744
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17972 12442 18000 12786
rect 18064 12646 18092 13194
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18050 12336 18106 12345
rect 18050 12271 18106 12280
rect 18064 11830 18092 12271
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8974 17632 9454
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 7954 17632 8910
rect 17696 8906 17724 9930
rect 17776 9716 17828 9722
rect 17880 9704 17908 10066
rect 17828 9676 17908 9704
rect 17776 9658 17828 9664
rect 17788 9586 17816 9658
rect 18156 9586 18184 29106
rect 18340 28490 18368 36110
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18432 24274 18460 37198
rect 18616 36174 18644 60998
rect 19260 60874 19288 63200
rect 19812 61198 19840 63294
rect 19982 63200 20038 63294
rect 20718 63200 20774 64000
rect 21454 63322 21510 64000
rect 21284 63294 21510 63322
rect 20628 61260 20680 61266
rect 20628 61202 20680 61208
rect 19800 61192 19852 61198
rect 19800 61134 19852 61140
rect 19984 61124 20036 61130
rect 19984 61066 20036 61072
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 19260 60846 19380 60874
rect 19352 60790 19380 60846
rect 19340 60784 19392 60790
rect 19340 60726 19392 60732
rect 19248 60308 19300 60314
rect 19248 60250 19300 60256
rect 19260 59702 19288 60250
rect 19996 60110 20024 61066
rect 20352 60580 20404 60586
rect 20352 60522 20404 60528
rect 19432 60104 19484 60110
rect 19432 60046 19484 60052
rect 19984 60104 20036 60110
rect 19984 60046 20036 60052
rect 19248 59696 19300 59702
rect 19248 59638 19300 59644
rect 18788 59628 18840 59634
rect 18788 59570 18840 59576
rect 19156 59628 19208 59634
rect 19156 59570 19208 59576
rect 18800 58682 18828 59570
rect 19168 59430 19196 59570
rect 19444 59566 19472 60046
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 19432 59560 19484 59566
rect 19432 59502 19484 59508
rect 19156 59424 19208 59430
rect 19156 59366 19208 59372
rect 19248 59424 19300 59430
rect 19248 59366 19300 59372
rect 18788 58676 18840 58682
rect 18788 58618 18840 58624
rect 19064 46436 19116 46442
rect 19064 46378 19116 46384
rect 18696 37188 18748 37194
rect 18696 37130 18748 37136
rect 18708 36854 18736 37130
rect 19076 36854 19104 46378
rect 19260 37874 19288 59366
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 20260 47592 20312 47598
rect 20260 47534 20312 47540
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19800 45348 19852 45354
rect 19800 45290 19852 45296
rect 19812 45082 19840 45290
rect 19800 45076 19852 45082
rect 19800 45018 19852 45024
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 20168 40724 20220 40730
rect 20168 40666 20220 40672
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19340 40112 19392 40118
rect 19340 40054 19392 40060
rect 19248 37868 19300 37874
rect 19248 37810 19300 37816
rect 19248 37188 19300 37194
rect 19248 37130 19300 37136
rect 18696 36848 18748 36854
rect 18696 36790 18748 36796
rect 19064 36848 19116 36854
rect 19064 36790 19116 36796
rect 19260 36786 19288 37130
rect 18880 36780 18932 36786
rect 18880 36722 18932 36728
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 18892 36666 18920 36722
rect 19154 36680 19210 36689
rect 18892 36638 19104 36666
rect 18880 36576 18932 36582
rect 18880 36518 18932 36524
rect 18972 36576 19024 36582
rect 18972 36518 19024 36524
rect 18892 36310 18920 36518
rect 18880 36304 18932 36310
rect 18880 36246 18932 36252
rect 18604 36168 18656 36174
rect 18604 36110 18656 36116
rect 18788 36168 18840 36174
rect 18788 36110 18840 36116
rect 18800 35986 18828 36110
rect 18984 35986 19012 36518
rect 19076 36378 19104 36638
rect 19154 36615 19156 36624
rect 19208 36615 19210 36624
rect 19156 36586 19208 36592
rect 19064 36372 19116 36378
rect 19064 36314 19116 36320
rect 18800 35958 19012 35986
rect 19352 35630 19380 40054
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38208 19484 38214
rect 19432 38150 19484 38156
rect 19444 37942 19472 38150
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 19522 37904 19578 37913
rect 19522 37839 19524 37848
rect 19576 37839 19578 37848
rect 19708 37868 19760 37874
rect 19524 37810 19576 37816
rect 19708 37810 19760 37816
rect 19720 37738 19748 37810
rect 19708 37732 19760 37738
rect 19708 37674 19760 37680
rect 20076 37664 20128 37670
rect 20076 37606 20128 37612
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20088 36786 20116 37606
rect 20180 37262 20208 40666
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20272 37194 20300 47534
rect 20260 37188 20312 37194
rect 20260 37130 20312 37136
rect 20076 36780 20128 36786
rect 20076 36722 20128 36728
rect 19432 36304 19484 36310
rect 19432 36246 19484 36252
rect 19340 35624 19392 35630
rect 19340 35566 19392 35572
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18248 16114 18276 18566
rect 18340 17218 18368 23530
rect 18432 23526 18460 24210
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18524 20074 18552 25638
rect 18708 24750 18736 29650
rect 19352 26234 19380 35022
rect 19444 34406 19472 36246
rect 19904 36230 20116 36258
rect 19904 36106 19932 36230
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19706 35048 19762 35057
rect 19706 34983 19708 34992
rect 19760 34983 19762 34992
rect 19708 34954 19760 34960
rect 19904 34932 19932 35498
rect 19996 35290 20024 36110
rect 20088 35630 20116 36230
rect 20364 36174 20392 60522
rect 20536 60240 20588 60246
rect 20536 60182 20588 60188
rect 20548 41414 20576 60182
rect 20456 41386 20576 41414
rect 20456 39250 20484 41386
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20548 39370 20576 40870
rect 20640 39438 20668 61202
rect 20732 61198 20760 63200
rect 21284 61198 21312 63294
rect 21454 63200 21510 63294
rect 22190 63322 22246 64000
rect 22926 63322 22982 64000
rect 22190 63294 22416 63322
rect 22190 63200 22246 63294
rect 22388 61198 22416 63294
rect 22926 63294 23336 63322
rect 22926 63200 22982 63294
rect 22836 61396 22888 61402
rect 22836 61338 22888 61344
rect 20720 61192 20772 61198
rect 20720 61134 20772 61140
rect 21272 61192 21324 61198
rect 21272 61134 21324 61140
rect 22376 61192 22428 61198
rect 22376 61134 22428 61140
rect 22284 61124 22336 61130
rect 22284 61066 22336 61072
rect 21456 61056 21508 61062
rect 21456 60998 21508 61004
rect 21272 60716 21324 60722
rect 21272 60658 21324 60664
rect 21284 60178 21312 60658
rect 21272 60172 21324 60178
rect 21272 60114 21324 60120
rect 21180 60104 21232 60110
rect 21178 60072 21180 60081
rect 21232 60072 21234 60081
rect 21178 60007 21234 60016
rect 21088 59492 21140 59498
rect 21088 59434 21140 59440
rect 21100 58857 21128 59434
rect 21086 58848 21142 58857
rect 21086 58783 21142 58792
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 20732 45558 20760 46310
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 21192 45286 21220 60007
rect 20812 45280 20864 45286
rect 20812 45222 20864 45228
rect 21180 45280 21232 45286
rect 21180 45222 21232 45228
rect 20824 41478 20852 45222
rect 20904 42152 20956 42158
rect 20904 42094 20956 42100
rect 20812 41472 20864 41478
rect 20812 41414 20864 41420
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20824 39370 20852 41414
rect 20536 39364 20588 39370
rect 20536 39306 20588 39312
rect 20812 39364 20864 39370
rect 20812 39306 20864 39312
rect 20456 39222 20668 39250
rect 20536 37664 20588 37670
rect 20536 37606 20588 37612
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20168 36032 20220 36038
rect 20168 35974 20220 35980
rect 20076 35624 20128 35630
rect 20076 35566 20128 35572
rect 19984 35284 20036 35290
rect 19984 35226 20036 35232
rect 20180 35057 20208 35974
rect 20260 35828 20312 35834
rect 20260 35770 20312 35776
rect 20166 35048 20222 35057
rect 20166 34983 20222 34992
rect 19904 34904 20024 34932
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34400 19484 34406
rect 19432 34342 19484 34348
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 19444 31346 19472 33050
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19524 31408 19576 31414
rect 19524 31350 19576 31356
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19444 30734 19472 31078
rect 19536 30938 19564 31350
rect 19708 31204 19760 31210
rect 19708 31146 19760 31152
rect 19720 30938 19748 31146
rect 19524 30932 19576 30938
rect 19524 30874 19576 30880
rect 19708 30932 19760 30938
rect 19708 30874 19760 30880
rect 19996 30870 20024 34904
rect 20076 31272 20128 31278
rect 20076 31214 20128 31220
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19616 30728 19668 30734
rect 20088 30705 20116 31214
rect 20168 30864 20220 30870
rect 20168 30806 20220 30812
rect 20074 30696 20130 30705
rect 19668 30676 20024 30682
rect 19616 30670 20024 30676
rect 19628 30654 20024 30670
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19352 26206 19472 26234
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18708 22094 18736 24686
rect 19444 24177 19472 26206
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24206 20024 30654
rect 20074 30631 20130 30640
rect 20180 29782 20208 30806
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 19984 24200 20036 24206
rect 19430 24168 19486 24177
rect 19984 24142 20036 24148
rect 19430 24103 19486 24112
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18984 22094 19012 23666
rect 20088 23118 20116 29446
rect 20180 29170 20208 29718
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 18708 22066 18920 22094
rect 18984 22066 19196 22094
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18524 20046 18736 20074
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18524 19394 18552 19722
rect 18432 19378 18552 19394
rect 18432 19372 18564 19378
rect 18432 19366 18512 19372
rect 18432 18766 18460 19366
rect 18512 19314 18564 19320
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18524 18834 18552 19178
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18524 18154 18552 18362
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18340 17190 18552 17218
rect 18616 17202 18644 19926
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18248 15638 18276 15846
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18340 15094 18368 16390
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 12986 18276 13670
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18234 12880 18290 12889
rect 18234 12815 18236 12824
rect 18288 12815 18290 12824
rect 18236 12786 18288 12792
rect 18340 11218 18368 15030
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18326 10976 18382 10985
rect 18326 10911 18382 10920
rect 18340 10674 18368 10911
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18432 10606 18460 17070
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18524 10130 18552 17190
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18616 16522 18644 17002
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18604 12776 18656 12782
rect 18602 12744 18604 12753
rect 18656 12744 18658 12753
rect 18602 12679 18658 12688
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18616 10849 18644 11630
rect 18708 11626 18736 20046
rect 18800 16590 18828 20402
rect 18892 17134 18920 22066
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18984 19854 19012 20266
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19145 19012 19790
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 19076 19310 19104 19654
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 18970 19136 19026 19145
rect 18970 19071 19026 19080
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18878 16960 18934 16969
rect 18878 16895 18934 16904
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 12442 18828 13194
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 11626 18828 11698
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18892 11506 18920 16895
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18800 11478 18920 11506
rect 18602 10840 18658 10849
rect 18602 10775 18658 10784
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17972 8945 18000 9046
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17958 8936 18014 8945
rect 17684 8900 17736 8906
rect 17958 8871 18014 8880
rect 17684 8842 17736 8848
rect 17682 8528 17738 8537
rect 17682 8463 17738 8472
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17604 7002 17632 7890
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17498 6216 17554 6225
rect 17498 6151 17554 6160
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17512 4622 17540 6151
rect 17604 5953 17632 6734
rect 17590 5944 17646 5953
rect 17590 5879 17646 5888
rect 17590 5808 17646 5817
rect 17590 5743 17646 5752
rect 17604 5710 17632 5743
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 4282 17264 4490
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 16948 4208 17000 4214
rect 16946 4176 16948 4185
rect 17000 4176 17002 4185
rect 16946 4111 17002 4120
rect 17592 4072 17644 4078
rect 17130 4040 17186 4049
rect 17592 4014 17644 4020
rect 17130 3975 17186 3984
rect 17144 3058 17172 3975
rect 17604 3738 17632 4014
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17696 3602 17724 8463
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6186 17816 6598
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17788 3194 17816 5578
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16960 1358 16988 2858
rect 17500 2440 17552 2446
rect 17130 2408 17186 2417
rect 17500 2382 17552 2388
rect 17130 2343 17186 2352
rect 16948 1352 17000 1358
rect 16948 1294 17000 1300
rect 17144 800 17172 2343
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 17236 1601 17264 2042
rect 17222 1592 17278 1601
rect 17222 1527 17278 1536
rect 17408 1488 17460 1494
rect 17408 1430 17460 1436
rect 17420 800 17448 1430
rect 17512 1329 17540 2382
rect 17498 1320 17554 1329
rect 17498 1255 17554 1264
rect 17696 800 17724 3130
rect 17972 2417 18000 7822
rect 18064 7342 18092 8978
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6866 18092 7278
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18156 6798 18184 9522
rect 18340 9518 18368 9998
rect 18708 9897 18736 10066
rect 18694 9888 18750 9897
rect 18694 9823 18750 9832
rect 18418 9752 18474 9761
rect 18418 9687 18474 9696
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18340 8974 18368 9454
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18248 8401 18276 8842
rect 18432 8616 18460 9687
rect 18510 9344 18566 9353
rect 18510 9279 18566 9288
rect 18340 8588 18460 8616
rect 18340 8498 18368 8588
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18234 8392 18290 8401
rect 18234 8327 18290 8336
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18248 7732 18276 8230
rect 18340 7886 18368 8434
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18432 7886 18460 7919
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18248 7704 18368 7732
rect 18340 7274 18368 7704
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18064 3534 18092 6394
rect 18156 5273 18184 6734
rect 18248 6361 18276 6802
rect 18340 6633 18368 7210
rect 18418 6896 18474 6905
rect 18418 6831 18474 6840
rect 18326 6624 18382 6633
rect 18326 6559 18382 6568
rect 18234 6352 18290 6361
rect 18234 6287 18290 6296
rect 18432 5710 18460 6831
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18142 5264 18198 5273
rect 18142 5199 18198 5208
rect 18418 4992 18474 5001
rect 18418 4927 18474 4936
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18064 2650 18092 2926
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17958 2408 18014 2417
rect 17776 2372 17828 2378
rect 17958 2343 18014 2352
rect 17776 2314 17828 2320
rect 17788 2038 17816 2314
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 18064 1737 18092 2450
rect 18050 1728 18106 1737
rect 18050 1663 18106 1672
rect 17960 1624 18012 1630
rect 17960 1566 18012 1572
rect 17972 800 18000 1566
rect 18156 1442 18184 3606
rect 18248 2774 18276 4014
rect 18340 2836 18368 4218
rect 18432 3534 18460 4927
rect 18524 4622 18552 9279
rect 18800 9217 18828 11478
rect 18878 11384 18934 11393
rect 18878 11319 18880 11328
rect 18932 11319 18934 11328
rect 18880 11290 18932 11296
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 9874 18920 11086
rect 18984 10674 19012 13398
rect 19168 12434 19196 22066
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 19260 19514 19288 21014
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19246 14240 19302 14249
rect 19246 14175 19302 14184
rect 19260 13938 19288 14175
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19076 12406 19196 12434
rect 19076 10690 19104 12406
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11762 19288 12174
rect 19352 11914 19380 23054
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19444 19854 19472 20334
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 19310 19472 19790
rect 19536 19718 19564 20402
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19720 20058 19748 20198
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 19904 19854 19932 20266
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19444 18766 19472 19246
rect 19996 19242 20024 20470
rect 20088 19242 20116 20878
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 20088 19122 20116 19178
rect 19996 19094 20116 19122
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 17678 19472 18702
rect 19996 18698 20024 19094
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19628 17134 19656 17206
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16658 19840 16934
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19444 15502 19472 16526
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 15609 20024 18294
rect 20180 17954 20208 28358
rect 20272 24138 20300 35770
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20364 30734 20392 34342
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20456 25906 20484 36654
rect 20548 36650 20576 37606
rect 20536 36644 20588 36650
rect 20536 36586 20588 36592
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20548 35630 20576 36110
rect 20536 35624 20588 35630
rect 20536 35566 20588 35572
rect 20640 33998 20668 39222
rect 20824 38654 20852 39306
rect 20732 38626 20852 38654
rect 20732 36174 20760 38626
rect 20916 38010 20944 42094
rect 21364 39296 21416 39302
rect 21364 39238 21416 39244
rect 20904 38004 20956 38010
rect 20904 37946 20956 37952
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 21100 36174 21128 37266
rect 21376 36174 21404 39238
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 21364 36168 21416 36174
rect 21364 36110 21416 36116
rect 20812 36100 20864 36106
rect 20812 36042 20864 36048
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20732 35222 20760 35974
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 20824 34474 20852 36042
rect 21364 35556 21416 35562
rect 21364 35498 21416 35504
rect 21376 35086 21404 35498
rect 21364 35080 21416 35086
rect 21364 35022 21416 35028
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 20812 34468 20864 34474
rect 20812 34410 20864 34416
rect 20628 33992 20680 33998
rect 20824 33946 20852 34410
rect 20628 33934 20680 33940
rect 20732 33930 20852 33946
rect 20720 33924 20852 33930
rect 20772 33918 20852 33924
rect 20720 33866 20772 33872
rect 21100 32978 21128 34886
rect 21272 34400 21324 34406
rect 21272 34342 21324 34348
rect 21284 33998 21312 34342
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21088 32972 21140 32978
rect 21088 32914 21140 32920
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20548 22094 20576 23462
rect 20456 22066 20576 22094
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20272 19514 20300 20402
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20364 18698 20392 21830
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20180 17926 20300 17954
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19982 15600 20038 15609
rect 19982 15535 20038 15544
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 14482 19472 15438
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 13394 19472 14418
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19444 12238 19472 13330
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19352 11886 19472 11914
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19168 10810 19196 11698
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19246 10704 19302 10713
rect 18972 10668 19024 10674
rect 19076 10662 19196 10690
rect 18972 10610 19024 10616
rect 18892 9846 19012 9874
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18892 9654 18920 9687
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18984 9586 19012 9846
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18786 9208 18842 9217
rect 18696 9172 18748 9178
rect 18616 9132 18696 9160
rect 18616 8952 18644 9132
rect 18786 9143 18842 9152
rect 18696 9114 18748 9120
rect 18604 8946 18656 8952
rect 18604 8888 18656 8894
rect 18788 8900 18840 8906
rect 18708 8860 18788 8888
rect 18604 8628 18656 8634
rect 18708 8616 18736 8860
rect 18788 8842 18840 8848
rect 18656 8588 18736 8616
rect 18604 8570 18656 8576
rect 18616 8276 18644 8570
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18616 8248 18736 8276
rect 18602 8120 18658 8129
rect 18602 8055 18658 8064
rect 18616 7886 18644 8055
rect 18708 7886 18736 8248
rect 18800 8022 18828 8502
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18800 7818 18828 7958
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18786 7712 18842 7721
rect 18786 7647 18842 7656
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18616 6866 18644 7210
rect 18708 6866 18736 7482
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18708 5778 18736 6258
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18800 5710 18828 7647
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18786 5128 18842 5137
rect 18786 5063 18842 5072
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 4049 18552 4082
rect 18696 4072 18748 4078
rect 18510 4040 18566 4049
rect 18696 4014 18748 4020
rect 18510 3975 18566 3984
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18340 2808 18460 2836
rect 18248 2746 18368 2774
rect 18156 1414 18276 1442
rect 18248 800 18276 1414
rect 18340 1034 18368 2746
rect 18432 1902 18460 2808
rect 18524 2446 18552 3703
rect 18602 3224 18658 3233
rect 18602 3159 18658 3168
rect 18616 2446 18644 3159
rect 18708 2689 18736 4014
rect 18800 3670 18828 5063
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18694 2680 18750 2689
rect 18694 2615 18750 2624
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18708 2106 18736 2314
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 18420 1896 18472 1902
rect 18420 1838 18472 1844
rect 18340 1006 18552 1034
rect 18524 800 18552 1006
rect 18800 800 18828 3130
rect 18892 3058 18920 9318
rect 18984 9178 19012 9318
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18984 8809 19012 8978
rect 19076 8945 19104 9046
rect 19062 8936 19118 8945
rect 19062 8871 19118 8880
rect 19064 8832 19116 8838
rect 18970 8800 19026 8809
rect 19064 8774 19116 8780
rect 18970 8735 19026 8744
rect 19076 8401 19104 8774
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19168 8129 19196 10662
rect 19246 10639 19302 10648
rect 19260 8634 19288 10639
rect 19352 9178 19380 11766
rect 19444 11150 19472 11886
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19536 10062 19564 10610
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10062 19748 10542
rect 19524 10056 19576 10062
rect 19430 10024 19486 10033
rect 19524 9998 19576 10004
rect 19708 10056 19760 10062
rect 19800 10056 19852 10062
rect 19708 9998 19760 10004
rect 19798 10024 19800 10033
rect 19852 10024 19854 10033
rect 19430 9959 19486 9968
rect 19798 9959 19854 9968
rect 19444 9926 19472 9959
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8634 19380 8910
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19352 8401 19380 8434
rect 19338 8392 19394 8401
rect 19338 8327 19394 8336
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19154 8120 19210 8129
rect 19154 8055 19210 8064
rect 19260 7970 19288 8230
rect 19168 7942 19288 7970
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7342 19012 7822
rect 19168 7721 19196 7942
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19444 7585 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19720 8945 19748 9522
rect 19798 9480 19854 9489
rect 19798 9415 19854 9424
rect 19812 8974 19840 9415
rect 19904 9382 19932 9522
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19800 8968 19852 8974
rect 19706 8936 19762 8945
rect 19800 8910 19852 8916
rect 19706 8871 19708 8880
rect 19760 8871 19762 8880
rect 19708 8842 19760 8848
rect 19720 8811 19748 8842
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8673 20024 15302
rect 20088 11558 20116 17818
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20088 10742 20116 11086
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19982 8664 20038 8673
rect 19982 8599 20038 8608
rect 20088 8566 20116 10542
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19800 8424 19852 8430
rect 19996 8401 20024 8434
rect 19800 8366 19852 8372
rect 19982 8392 20038 8401
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19720 7954 19748 8230
rect 19812 7993 19840 8366
rect 19982 8327 20038 8336
rect 19798 7984 19854 7993
rect 19708 7948 19760 7954
rect 19798 7919 19854 7928
rect 19708 7890 19760 7896
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19430 7576 19486 7585
rect 19574 7579 19882 7588
rect 19996 7585 20024 7754
rect 19340 7540 19392 7546
rect 19982 7576 20038 7585
rect 19430 7511 19486 7520
rect 19904 7520 19982 7528
rect 19904 7511 20038 7520
rect 19340 7482 19392 7488
rect 19904 7500 20024 7511
rect 19352 7410 19380 7482
rect 19340 7404 19392 7410
rect 19524 7404 19576 7410
rect 19340 7346 19392 7352
rect 19444 7364 19524 7392
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19076 7154 19104 7210
rect 19076 7126 19288 7154
rect 19260 7018 19288 7126
rect 19260 7002 19334 7018
rect 19444 7002 19472 7364
rect 19800 7404 19852 7410
rect 19576 7364 19656 7392
rect 19524 7346 19576 7352
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19536 7002 19564 7142
rect 19260 6996 19346 7002
rect 19260 6990 19294 6996
rect 19294 6938 19346 6944
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19628 6730 19656 7364
rect 19800 7346 19852 7352
rect 19812 6798 19840 7346
rect 19904 7342 19932 7500
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 18984 6254 19012 6666
rect 19062 6624 19118 6633
rect 19062 6559 19118 6568
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 18984 5166 19012 5850
rect 19076 5166 19104 6559
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19338 6488 19394 6497
rect 19574 6491 19882 6500
rect 19338 6423 19340 6432
rect 19392 6423 19394 6432
rect 19984 6452 20036 6458
rect 19340 6394 19392 6400
rect 19984 6394 20036 6400
rect 19246 6352 19302 6361
rect 19996 6322 20024 6394
rect 20088 6322 20116 6734
rect 19246 6287 19248 6296
rect 19300 6287 19302 6296
rect 19984 6316 20036 6322
rect 19248 6258 19300 6264
rect 19984 6258 20036 6264
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19892 6248 19944 6254
rect 20180 6202 20208 17070
rect 20272 13258 20300 17926
rect 20456 15586 20484 22066
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 18766 20576 20742
rect 20640 20602 20668 21422
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20732 20602 20760 20810
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20732 20262 20760 20538
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20548 18154 20576 18702
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 15638 20576 17138
rect 20640 16590 20668 19110
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17134 20760 17614
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20824 16998 20852 20742
rect 20916 20058 20944 21558
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20916 17066 20944 17750
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20364 15558 20484 15586
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20364 14521 20392 15558
rect 20904 15360 20956 15366
rect 20534 15328 20590 15337
rect 20904 15302 20956 15308
rect 20534 15263 20590 15272
rect 20350 14512 20406 14521
rect 20350 14447 20406 14456
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20272 12782 20300 12854
rect 20364 12782 20392 14447
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20272 11898 20300 12106
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20364 11801 20392 12582
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11898 20484 12038
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20350 11792 20406 11801
rect 20350 11727 20406 11736
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11218 20300 11494
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20350 10976 20406 10985
rect 20350 10911 20406 10920
rect 20364 10588 20392 10911
rect 20456 10849 20484 11562
rect 20442 10840 20498 10849
rect 20442 10775 20498 10784
rect 20272 10560 20392 10588
rect 20272 8498 20300 10560
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10198 20392 10406
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20456 9994 20484 10775
rect 20548 10062 20576 15263
rect 20916 15094 20944 15302
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14550 20944 14758
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20812 13184 20864 13190
rect 20810 13152 20812 13161
rect 20864 13152 20866 13161
rect 20810 13087 20866 13096
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20732 12374 20760 12650
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20824 11914 20852 12718
rect 20640 11886 20852 11914
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20442 9888 20498 9897
rect 20640 9874 20668 11886
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20824 11529 20852 11727
rect 20810 11520 20866 11529
rect 20810 11455 20866 11464
rect 20916 11336 20944 13194
rect 20824 11308 20944 11336
rect 20824 10985 20852 11308
rect 20810 10976 20866 10985
rect 20810 10911 20866 10920
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10130 20760 10406
rect 20824 10198 20852 10610
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20916 10062 20944 10678
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 21008 9926 21036 26862
rect 21468 22137 21496 60998
rect 22192 60852 22244 60858
rect 22192 60794 22244 60800
rect 22100 60716 22152 60722
rect 22100 60658 22152 60664
rect 22112 59401 22140 60658
rect 22204 59634 22232 60794
rect 22296 60110 22324 61066
rect 22848 60734 22876 61338
rect 23308 60790 23336 63294
rect 23662 63200 23718 64000
rect 24398 63322 24454 64000
rect 24398 63294 24624 63322
rect 24398 63200 24454 63294
rect 23676 61198 23704 63200
rect 23664 61192 23716 61198
rect 23664 61134 23716 61140
rect 23756 61056 23808 61062
rect 23756 60998 23808 61004
rect 23296 60784 23348 60790
rect 22848 60706 22968 60734
rect 23296 60726 23348 60732
rect 22468 60648 22520 60654
rect 22468 60590 22520 60596
rect 22652 60648 22704 60654
rect 22652 60590 22704 60596
rect 22284 60104 22336 60110
rect 22284 60046 22336 60052
rect 22192 59628 22244 59634
rect 22192 59570 22244 59576
rect 22098 59392 22154 59401
rect 22098 59327 22154 59336
rect 22480 56846 22508 60590
rect 22664 60246 22692 60590
rect 22836 60512 22888 60518
rect 22836 60454 22888 60460
rect 22652 60240 22704 60246
rect 22652 60182 22704 60188
rect 22848 60194 22876 60454
rect 22940 60314 22968 60706
rect 22928 60308 22980 60314
rect 22928 60250 22980 60256
rect 22664 60110 22692 60182
rect 22848 60166 23060 60194
rect 23032 60110 23060 60166
rect 22652 60104 22704 60110
rect 22652 60046 22704 60052
rect 23020 60104 23072 60110
rect 23020 60046 23072 60052
rect 22560 60036 22612 60042
rect 22560 59978 22612 59984
rect 22744 60036 22796 60042
rect 22744 59978 22796 59984
rect 23572 60036 23624 60042
rect 23572 59978 23624 59984
rect 22572 59537 22600 59978
rect 22650 59800 22706 59809
rect 22650 59735 22706 59744
rect 22664 59702 22692 59735
rect 22652 59696 22704 59702
rect 22652 59638 22704 59644
rect 22558 59528 22614 59537
rect 22558 59463 22614 59472
rect 22468 56840 22520 56846
rect 22468 56782 22520 56788
rect 22284 49768 22336 49774
rect 22284 49710 22336 49716
rect 22192 47592 22244 47598
rect 22192 47534 22244 47540
rect 22008 43444 22060 43450
rect 22008 43386 22060 43392
rect 21640 37120 21692 37126
rect 21640 37062 21692 37068
rect 21548 36032 21600 36038
rect 21548 35974 21600 35980
rect 21454 22128 21510 22137
rect 21454 22063 21510 22072
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21100 19378 21128 21286
rect 21192 19854 21220 21558
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 20942 21312 21286
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21284 20602 21312 20742
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 21100 18290 21128 18566
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21192 17338 21220 19790
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18358 21312 18566
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21468 17746 21496 19314
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 9926 21128 11086
rect 20996 9920 21048 9926
rect 20640 9846 20944 9874
rect 20996 9862 21048 9868
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 20442 9823 20498 9832
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20364 8838 20392 8978
rect 20456 8906 20484 9823
rect 20718 9752 20774 9761
rect 20718 9687 20774 9696
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20640 9489 20668 9522
rect 20626 9480 20682 9489
rect 20732 9450 20760 9687
rect 20916 9654 20944 9846
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20824 9450 20852 9590
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20626 9415 20682 9424
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20626 9208 20682 9217
rect 20682 9166 20760 9194
rect 20626 9143 20682 9152
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20640 8922 20668 8978
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20548 8894 20668 8922
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20442 8800 20498 8809
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20272 8401 20300 8434
rect 20258 8392 20314 8401
rect 20258 8327 20314 8336
rect 20258 7984 20314 7993
rect 20258 7919 20260 7928
rect 20312 7919 20314 7928
rect 20260 7890 20312 7896
rect 20272 7410 20300 7890
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20272 6905 20300 7210
rect 20258 6896 20314 6905
rect 20258 6831 20314 6840
rect 20272 6798 20300 6831
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20364 6662 20392 8774
rect 20442 8735 20498 8744
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20456 6361 20484 8735
rect 20548 8129 20576 8894
rect 20732 8378 20760 9166
rect 20916 8906 20944 9454
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8566 20852 8774
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20640 8350 20760 8378
rect 20534 8120 20590 8129
rect 20534 8055 20590 8064
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20548 6474 20576 7958
rect 20640 6798 20668 8350
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20732 7274 20760 8026
rect 20916 7954 20944 8842
rect 21008 8430 21036 9862
rect 21086 8664 21142 8673
rect 21086 8599 21142 8608
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21100 8090 21128 8599
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20812 7880 20864 7886
rect 20810 7848 20812 7857
rect 20864 7848 20866 7857
rect 20810 7783 20866 7792
rect 20824 7410 20852 7783
rect 20902 7576 20958 7585
rect 20902 7511 20904 7520
rect 20956 7511 20958 7520
rect 21088 7540 21140 7546
rect 20904 7482 20956 7488
rect 21088 7482 21140 7488
rect 20916 7410 20944 7482
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20718 6896 20774 6905
rect 20718 6831 20774 6840
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20548 6446 20668 6474
rect 20536 6384 20588 6390
rect 20442 6352 20498 6361
rect 20260 6316 20312 6322
rect 20536 6326 20588 6332
rect 20442 6287 20498 6296
rect 20260 6258 20312 6264
rect 19892 6190 19944 6196
rect 19904 5778 19932 6190
rect 20088 6174 20208 6202
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19352 5302 19380 5714
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19996 5234 20024 5578
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19260 5098 19288 5170
rect 19338 5128 19394 5137
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 19248 5092 19300 5098
rect 19338 5063 19394 5072
rect 19248 5034 19300 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 4690 19104 4966
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18984 2774 19012 3402
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18892 2746 19012 2774
rect 6184 750 6236 756
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 18892 542 18920 2746
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18984 610 19012 2586
rect 19076 800 19104 3334
rect 19168 2514 19196 5034
rect 19352 4604 19380 5063
rect 19444 4826 19472 5170
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19260 4576 19380 4604
rect 19616 4616 19668 4622
rect 19260 4214 19288 4576
rect 19616 4558 19668 4564
rect 19628 4468 19656 4558
rect 19628 4457 20024 4468
rect 19628 4448 20038 4457
rect 19628 4440 19982 4448
rect 19574 4380 19882 4389
rect 19982 4383 20038 4392
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19708 4276 19760 4282
rect 20088 4264 20116 6174
rect 20272 5914 20300 6258
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20272 5710 20300 5850
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20260 5568 20312 5574
rect 20166 5536 20222 5545
rect 20260 5510 20312 5516
rect 20166 5471 20222 5480
rect 19708 4218 19760 4224
rect 19812 4236 20116 4264
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 19352 3738 19380 4218
rect 19720 4162 19748 4218
rect 19812 4162 19840 4236
rect 19616 4140 19668 4146
rect 19720 4134 19840 4162
rect 19616 4082 19668 4088
rect 19432 4072 19484 4078
rect 19430 4040 19432 4049
rect 19484 4040 19486 4049
rect 19430 3975 19486 3984
rect 19628 3992 19656 4082
rect 19628 3964 19758 3992
rect 19614 3768 19670 3777
rect 19340 3732 19392 3738
rect 19730 3754 19758 3964
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19614 3703 19670 3712
rect 19720 3726 19758 3754
rect 19340 3674 19392 3680
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3194 19288 3538
rect 19628 3534 19656 3703
rect 19720 3670 19748 3726
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19996 3602 20024 3878
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19352 3346 19380 3470
rect 20180 3448 20208 5471
rect 20272 5409 20300 5510
rect 20258 5400 20314 5409
rect 20258 5335 20314 5344
rect 20350 5128 20406 5137
rect 20260 5092 20312 5098
rect 20350 5063 20406 5072
rect 20260 5034 20312 5040
rect 20272 3720 20300 5034
rect 20364 4282 20392 5063
rect 20442 4312 20498 4321
rect 20352 4276 20404 4282
rect 20442 4247 20498 4256
rect 20352 4218 20404 4224
rect 20456 4214 20484 4247
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20272 3692 20484 3720
rect 19830 3420 20208 3448
rect 19708 3392 19760 3398
rect 19352 3318 19472 3346
rect 19830 3380 19858 3420
rect 19760 3352 19858 3380
rect 19708 3334 19760 3340
rect 19444 3233 19472 3318
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19430 3224 19486 3233
rect 19574 3227 19882 3236
rect 19248 3188 19300 3194
rect 19430 3159 19486 3168
rect 20074 3224 20130 3233
rect 20456 3210 20484 3692
rect 20074 3159 20130 3168
rect 20180 3182 20484 3210
rect 19248 3130 19300 3136
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 1630 19288 2246
rect 19248 1624 19300 1630
rect 19248 1566 19300 1572
rect 19444 1442 19472 2790
rect 19536 2378 19564 2994
rect 19720 2650 19748 2994
rect 19812 2961 19840 2994
rect 19984 2984 20036 2990
rect 19798 2952 19854 2961
rect 19798 2887 19854 2896
rect 19982 2952 19984 2961
rect 20036 2952 20038 2961
rect 19982 2887 20038 2896
rect 20088 2825 20116 3159
rect 20074 2816 20130 2825
rect 20074 2751 20130 2760
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19982 2544 20038 2553
rect 19982 2479 20038 2488
rect 19996 2446 20024 2479
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19524 2372 19576 2378
rect 19524 2314 19576 2320
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 19248 1420 19300 1426
rect 19444 1414 19656 1442
rect 19248 1362 19300 1368
rect 19260 1306 19288 1362
rect 19260 1278 19380 1306
rect 19352 800 19380 1278
rect 19628 800 19656 1414
rect 19904 800 19932 1838
rect 20088 1426 20116 2314
rect 20076 1420 20128 1426
rect 20076 1362 20128 1368
rect 20180 800 20208 3182
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20272 1902 20300 2314
rect 20260 1896 20312 1902
rect 20260 1838 20312 1844
rect 20364 1494 20392 2858
rect 20456 1873 20484 3062
rect 20548 3058 20576 6326
rect 20640 5234 20668 6446
rect 20732 6322 20760 6831
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20916 5574 20944 7346
rect 21100 6798 21128 7482
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21100 6458 21128 6734
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 21008 5166 21036 5850
rect 21100 5778 21128 6394
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20824 4622 20852 5102
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20640 4146 20668 4490
rect 20732 4321 20760 4558
rect 20718 4312 20774 4321
rect 20718 4247 20774 4256
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20626 3768 20682 3777
rect 20626 3703 20682 3712
rect 20640 3534 20668 3703
rect 20824 3534 20852 4082
rect 20916 3534 20944 4218
rect 21008 4146 21036 4694
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20732 2990 20760 3402
rect 20824 3058 20852 3470
rect 20904 3392 20956 3398
rect 20902 3360 20904 3369
rect 20956 3360 20958 3369
rect 20902 3295 20958 3304
rect 21008 3194 21036 3946
rect 21100 3466 21128 4626
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20812 2916 20864 2922
rect 20812 2858 20864 2864
rect 20718 2816 20774 2825
rect 20824 2802 20852 2858
rect 20902 2816 20958 2825
rect 20824 2774 20902 2802
rect 20718 2751 20774 2760
rect 20902 2751 20958 2760
rect 20626 2680 20682 2689
rect 20626 2615 20682 2624
rect 20442 1864 20498 1873
rect 20442 1799 20498 1808
rect 20640 1766 20668 2615
rect 20444 1760 20496 1766
rect 20444 1702 20496 1708
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 20352 1488 20404 1494
rect 20352 1430 20404 1436
rect 20456 800 20484 1702
rect 20732 800 20760 2751
rect 20902 2680 20958 2689
rect 20902 2615 20958 2624
rect 20916 2446 20944 2615
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 21192 2310 21220 15982
rect 21376 15502 21404 17070
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 11830 21312 12378
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21270 11112 21326 11121
rect 21270 11047 21326 11056
rect 21284 10742 21312 11047
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21284 9926 21312 9998
rect 21376 9926 21404 11698
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21284 7818 21312 9862
rect 21376 9586 21404 9862
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 7868 21404 9318
rect 21468 8634 21496 13126
rect 21560 13025 21588 35974
rect 21652 32978 21680 37062
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 21836 35290 21864 35430
rect 21824 35284 21876 35290
rect 21824 35226 21876 35232
rect 22020 33522 22048 43386
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 22112 38593 22140 39374
rect 22098 38584 22154 38593
rect 22098 38519 22154 38528
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 22112 35086 22140 37402
rect 22204 35698 22232 47534
rect 22296 36106 22324 49710
rect 22376 40996 22428 41002
rect 22376 40938 22428 40944
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22098 34640 22154 34649
rect 22098 34575 22100 34584
rect 22152 34575 22154 34584
rect 22100 34546 22152 34552
rect 22204 34513 22232 35634
rect 22388 34746 22416 40938
rect 22756 38350 22784 59978
rect 23584 59770 23612 59978
rect 23572 59764 23624 59770
rect 23572 59706 23624 59712
rect 23572 55752 23624 55758
rect 23572 55694 23624 55700
rect 23584 54738 23612 55694
rect 23572 54732 23624 54738
rect 23572 54674 23624 54680
rect 22836 54596 22888 54602
rect 22836 54538 22888 54544
rect 22848 44878 22876 54538
rect 23572 52896 23624 52902
rect 23572 52838 23624 52844
rect 22836 44872 22888 44878
rect 22836 44814 22888 44820
rect 23480 42356 23532 42362
rect 23480 42298 23532 42304
rect 23202 38584 23258 38593
rect 23202 38519 23258 38528
rect 23216 38350 23244 38519
rect 23492 38418 23520 42298
rect 23480 38412 23532 38418
rect 23480 38354 23532 38360
rect 22744 38344 22796 38350
rect 22744 38286 22796 38292
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 22940 38010 22968 38286
rect 23020 38276 23072 38282
rect 23020 38218 23072 38224
rect 22928 38004 22980 38010
rect 22928 37946 22980 37952
rect 22560 37732 22612 37738
rect 22560 37674 22612 37680
rect 22468 36304 22520 36310
rect 22468 36246 22520 36252
rect 22480 36174 22508 36246
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22190 34504 22246 34513
rect 22190 34439 22246 34448
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 22112 33522 22140 34342
rect 22296 33862 22324 34546
rect 22480 33998 22508 34886
rect 22572 34610 22600 37674
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22848 36174 22876 36654
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22652 36100 22704 36106
rect 22652 36042 22704 36048
rect 22664 36009 22692 36042
rect 22650 36000 22706 36009
rect 22650 35935 22706 35944
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22560 34060 22612 34066
rect 22560 34002 22612 34008
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21836 25838 21864 31962
rect 22572 28529 22600 34002
rect 22664 31346 22692 35022
rect 22756 34678 22784 35430
rect 23032 35057 23060 38218
rect 23296 36304 23348 36310
rect 23296 36246 23348 36252
rect 23018 35048 23074 35057
rect 23018 34983 23074 34992
rect 22744 34672 22796 34678
rect 22744 34614 22796 34620
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22744 34536 22796 34542
rect 22744 34478 22796 34484
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22664 31142 22692 31282
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22558 28520 22614 28529
rect 22558 28455 22614 28464
rect 21824 25832 21876 25838
rect 21824 25774 21876 25780
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21638 19544 21694 19553
rect 21638 19479 21694 19488
rect 21652 19378 21680 19479
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21744 18766 21772 22102
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21730 17640 21786 17649
rect 21730 17575 21786 17584
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21546 13016 21602 13025
rect 21546 12951 21602 12960
rect 21652 12889 21680 13262
rect 21638 12880 21694 12889
rect 21638 12815 21694 12824
rect 21744 12434 21772 17575
rect 21836 13802 21864 25774
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22020 20516 22048 21082
rect 22112 20942 22140 22374
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22100 20528 22152 20534
rect 22020 20488 22100 20516
rect 22100 20470 22152 20476
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21928 17134 21956 20402
rect 22112 19825 22140 20470
rect 22098 19816 22154 19825
rect 22098 19751 22154 19760
rect 22006 19348 22062 19357
rect 22006 19283 22062 19292
rect 22020 18970 22048 19283
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22112 18034 22140 19751
rect 22190 19544 22246 19553
rect 22190 19479 22246 19488
rect 22204 18154 22232 19479
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22112 18006 22232 18034
rect 22204 17202 22232 18006
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 22296 16182 22324 23258
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 22480 22098 22508 22986
rect 22468 22092 22520 22098
rect 22664 22094 22692 29786
rect 22756 22681 22784 34478
rect 22848 30394 22876 34546
rect 23204 34468 23256 34474
rect 23204 34410 23256 34416
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22940 30734 22968 31690
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 22836 30388 22888 30394
rect 22836 30330 22888 30336
rect 22742 22672 22798 22681
rect 22742 22607 22798 22616
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22468 22034 22520 22040
rect 22572 22066 22692 22094
rect 22480 21486 22508 22034
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 22388 19242 22416 20266
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 19145 22416 19178
rect 22374 19136 22430 19145
rect 22374 19071 22430 19080
rect 22480 18970 22508 19722
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22006 15464 22062 15473
rect 22006 15399 22062 15408
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21928 13326 21956 13466
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 22020 12866 22048 15399
rect 22112 15026 22140 16118
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22098 14920 22154 14929
rect 22098 14855 22154 14864
rect 22112 14550 22140 14855
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22020 12838 22140 12866
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21652 12406 21772 12434
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21560 10985 21588 11086
rect 21546 10976 21602 10985
rect 21546 10911 21602 10920
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21560 9178 21588 10066
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21456 7880 21508 7886
rect 21376 7840 21456 7868
rect 21456 7822 21508 7828
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 7324 21312 7754
rect 21468 7585 21496 7822
rect 21454 7576 21510 7585
rect 21560 7546 21588 9114
rect 21454 7511 21510 7520
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21364 7336 21416 7342
rect 21284 7296 21364 7324
rect 21284 6730 21312 7296
rect 21364 7278 21416 7284
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21272 6724 21324 6730
rect 21272 6666 21324 6672
rect 21284 6322 21312 6666
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5642 21312 6258
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21284 4690 21312 5578
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21270 3632 21326 3641
rect 21270 3567 21326 3576
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 20996 1420 21048 1426
rect 20996 1362 21048 1368
rect 21008 800 21036 1362
rect 21284 800 21312 3567
rect 21376 3126 21404 4966
rect 21468 4690 21496 7210
rect 21560 7177 21588 7278
rect 21546 7168 21602 7177
rect 21546 7103 21602 7112
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21546 4312 21602 4321
rect 21546 4247 21602 4256
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21376 2310 21404 2926
rect 21468 2650 21496 3062
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21560 800 21588 4247
rect 21652 4010 21680 12406
rect 22020 12170 22048 12718
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21732 11280 21784 11286
rect 21732 11222 21784 11228
rect 21744 7954 21772 11222
rect 21836 8498 21864 11766
rect 22020 11762 22048 12106
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 21916 11688 21968 11694
rect 22112 11642 22140 12838
rect 22204 11744 22232 13806
rect 22296 12918 22324 14758
rect 22480 13870 22508 15030
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22388 12434 22416 13738
rect 22480 13326 22508 13806
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22388 12406 22508 12434
rect 22284 11756 22336 11762
rect 22204 11716 22284 11744
rect 22284 11698 22336 11704
rect 21916 11630 21968 11636
rect 21928 11529 21956 11630
rect 22020 11614 22140 11642
rect 21914 11520 21970 11529
rect 21914 11455 21970 11464
rect 21914 11112 21970 11121
rect 21914 11047 21916 11056
rect 21968 11047 21970 11056
rect 21916 11018 21968 11024
rect 21914 10704 21970 10713
rect 21914 10639 21970 10648
rect 21928 10130 21956 10639
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21928 9042 21956 9522
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21744 6390 21772 7686
rect 21732 6384 21784 6390
rect 21732 6326 21784 6332
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21744 4214 21772 6190
rect 21836 5710 21864 8026
rect 21928 7993 21956 8978
rect 21914 7984 21970 7993
rect 21914 7919 21970 7928
rect 22020 7698 22048 11614
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22112 10062 22140 11154
rect 22192 11144 22244 11150
rect 22190 11112 22192 11121
rect 22244 11112 22246 11121
rect 22190 11047 22246 11056
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22388 10713 22416 10746
rect 22190 10704 22246 10713
rect 22190 10639 22192 10648
rect 22244 10639 22246 10648
rect 22374 10704 22430 10713
rect 22374 10639 22430 10648
rect 22192 10610 22244 10616
rect 22284 10600 22336 10606
rect 22204 10548 22284 10554
rect 22204 10542 22336 10548
rect 22204 10526 22324 10542
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22112 9738 22140 9998
rect 22204 9926 22232 10526
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 9994 22324 10406
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22112 9710 22324 9738
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22112 8974 22140 9454
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 22100 8832 22152 8838
rect 22098 8800 22100 8809
rect 22152 8800 22154 8809
rect 22098 8735 22154 8744
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 21928 7670 22048 7698
rect 21928 6254 21956 7670
rect 22006 7576 22062 7585
rect 22006 7511 22062 7520
rect 22020 7410 22048 7511
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22112 6934 22140 7890
rect 22204 7206 22232 9522
rect 22296 8838 22324 9710
rect 22480 9602 22508 12406
rect 22572 10606 22600 22066
rect 22848 21690 22876 22578
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22664 19417 22692 21490
rect 22940 20890 22968 30670
rect 23032 23254 23060 31962
rect 23216 29578 23244 34410
rect 23204 29572 23256 29578
rect 23204 29514 23256 29520
rect 23020 23248 23072 23254
rect 23020 23190 23072 23196
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 23032 21554 23060 21898
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 22940 20862 23060 20890
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22742 19544 22798 19553
rect 22742 19479 22798 19488
rect 22756 19446 22784 19479
rect 22744 19440 22796 19446
rect 22650 19408 22706 19417
rect 22744 19382 22796 19388
rect 22940 19378 22968 20742
rect 22650 19343 22706 19352
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22742 18048 22798 18057
rect 22742 17983 22798 17992
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22664 13734 22692 14418
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22572 9722 22600 10542
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22480 9574 22600 9602
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22374 8800 22430 8809
rect 22296 7818 22324 8774
rect 22374 8735 22430 8744
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22296 7721 22324 7754
rect 22282 7712 22338 7721
rect 22282 7647 22338 7656
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22100 6928 22152 6934
rect 22296 6882 22324 7482
rect 22100 6870 22152 6876
rect 22204 6854 22324 6882
rect 22204 6798 22232 6854
rect 22192 6792 22244 6798
rect 22098 6760 22154 6769
rect 22304 6792 22356 6798
rect 22192 6734 22244 6740
rect 22296 6740 22304 6746
rect 22296 6734 22356 6740
rect 22098 6695 22154 6704
rect 22296 6718 22344 6734
rect 22112 6390 22140 6695
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21916 6112 21968 6118
rect 21914 6080 21916 6089
rect 21968 6080 21970 6089
rect 21914 6015 21970 6024
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21640 4004 21692 4010
rect 21640 3946 21692 3952
rect 21836 3942 21864 5170
rect 22020 4758 22048 6258
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22098 6080 22154 6089
rect 22098 6015 22154 6024
rect 22112 5574 22140 6015
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22204 4622 22232 6122
rect 22296 6118 22324 6718
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22112 4282 22140 4558
rect 22204 4282 22232 4558
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21914 3904 21970 3913
rect 21836 3777 21864 3878
rect 21970 3862 22048 3890
rect 21914 3839 21970 3848
rect 21822 3768 21878 3777
rect 21822 3703 21878 3712
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 18972 604 19024 610
rect 18972 546 19024 552
rect 18880 536 18932 542
rect 18880 478 18932 484
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21546 0 21602 800
rect 21652 678 21680 3402
rect 22020 2774 22048 3862
rect 22296 3534 22324 6054
rect 22388 4146 22416 8735
rect 22480 8090 22508 8910
rect 22572 8401 22600 9574
rect 22558 8392 22614 8401
rect 22558 8327 22614 8336
rect 22558 8120 22614 8129
rect 22468 8084 22520 8090
rect 22558 8055 22614 8064
rect 22468 8026 22520 8032
rect 22572 7954 22600 8055
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22466 6896 22522 6905
rect 22466 6831 22522 6840
rect 22480 6798 22508 6831
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22466 6488 22522 6497
rect 22466 6423 22522 6432
rect 22480 6322 22508 6423
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22468 5228 22520 5234
rect 22572 5216 22600 7890
rect 22664 6458 22692 10610
rect 22756 9518 22784 17983
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 16182 22968 16390
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22848 14414 22876 14758
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22834 13288 22890 13297
rect 22834 13223 22890 13232
rect 22848 10810 22876 13223
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22926 9344 22982 9353
rect 22926 9279 22982 9288
rect 22940 8974 22968 9279
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22836 8424 22888 8430
rect 23032 8412 23060 20862
rect 23124 20262 23152 21422
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23124 18630 23152 18906
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 23124 16590 23152 17002
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 14414 23152 16390
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23124 12102 23152 13670
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23124 11694 23152 11834
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 22888 8384 23060 8412
rect 22836 8366 22888 8372
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22756 6304 22784 7482
rect 22848 6866 22876 8366
rect 23124 7857 23152 9998
rect 23110 7848 23166 7857
rect 23110 7783 23166 7792
rect 23124 7546 23152 7783
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22520 5188 22600 5216
rect 22664 6276 22784 6304
rect 22468 5170 22520 5176
rect 22480 4457 22508 5170
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22466 4448 22522 4457
rect 22466 4383 22522 4392
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22284 3528 22336 3534
rect 22190 3496 22246 3505
rect 22284 3470 22336 3476
rect 22190 3431 22192 3440
rect 22244 3431 22246 3440
rect 22192 3402 22244 3408
rect 22480 3398 22508 4150
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22572 3126 22600 4626
rect 22664 4570 22692 6276
rect 22848 5953 22876 6394
rect 22834 5944 22890 5953
rect 22834 5879 22890 5888
rect 22848 5778 22876 5879
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22834 5264 22890 5273
rect 22834 5199 22836 5208
rect 22888 5199 22890 5208
rect 22836 5170 22888 5176
rect 22664 4542 22876 4570
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22560 3120 22612 3126
rect 22098 3088 22154 3097
rect 22560 3062 22612 3068
rect 22098 3023 22154 3032
rect 21836 2746 22048 2774
rect 21836 800 21864 2746
rect 22006 2680 22062 2689
rect 22006 2615 22062 2624
rect 22020 2582 22048 2615
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22112 800 22140 3023
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22296 1426 22324 2382
rect 22284 1420 22336 1426
rect 22284 1362 22336 1368
rect 22388 800 22416 2790
rect 22480 2514 22508 2858
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22664 800 22692 4422
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22756 4049 22784 4082
rect 22742 4040 22798 4049
rect 22742 3975 22798 3984
rect 22848 3942 22876 4542
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22940 3738 22968 6938
rect 23112 6792 23164 6798
rect 23018 6760 23074 6769
rect 23112 6734 23164 6740
rect 23018 6695 23074 6704
rect 23032 6662 23060 6695
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23124 6474 23152 6734
rect 23032 6446 23152 6474
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23032 3602 23060 6446
rect 23216 6322 23244 29514
rect 23308 26926 23336 36246
rect 23480 36100 23532 36106
rect 23480 36042 23532 36048
rect 23492 35834 23520 36042
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23478 35048 23534 35057
rect 23478 34983 23534 34992
rect 23492 34610 23520 34983
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 23492 29850 23520 34546
rect 23480 29844 23532 29850
rect 23480 29786 23532 29792
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23492 29306 23520 29582
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23584 29170 23612 52838
rect 23768 41750 23796 60998
rect 24596 60790 24624 63294
rect 25134 63200 25190 64000
rect 25870 63200 25926 64000
rect 26606 63200 26662 64000
rect 27342 63322 27398 64000
rect 27342 63294 27568 63322
rect 27342 63200 27398 63294
rect 24952 61668 25004 61674
rect 24952 61610 25004 61616
rect 24584 60784 24636 60790
rect 24584 60726 24636 60732
rect 24676 60716 24728 60722
rect 24676 60658 24728 60664
rect 24492 60580 24544 60586
rect 24492 60522 24544 60528
rect 24400 60512 24452 60518
rect 24400 60454 24452 60460
rect 23848 60104 23900 60110
rect 23848 60046 23900 60052
rect 23940 60104 23992 60110
rect 23940 60046 23992 60052
rect 23860 59945 23888 60046
rect 23846 59936 23902 59945
rect 23846 59871 23902 59880
rect 23860 53106 23888 59871
rect 23952 55706 23980 60046
rect 23952 55678 24072 55706
rect 23940 54664 23992 54670
rect 23940 54606 23992 54612
rect 23952 53242 23980 54606
rect 23940 53236 23992 53242
rect 23940 53178 23992 53184
rect 23848 53100 23900 53106
rect 23848 53042 23900 53048
rect 23756 41744 23808 41750
rect 23756 41686 23808 41692
rect 24044 41614 24072 55678
rect 24308 53100 24360 53106
rect 24308 53042 24360 53048
rect 24216 50380 24268 50386
rect 24216 50322 24268 50328
rect 24228 45554 24256 50322
rect 24136 45526 24256 45554
rect 24136 45490 24164 45526
rect 24124 45484 24176 45490
rect 24124 45426 24176 45432
rect 24124 41676 24176 41682
rect 24124 41618 24176 41624
rect 24032 41608 24084 41614
rect 24032 41550 24084 41556
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23676 36174 23704 38150
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35630 23704 35974
rect 23768 35766 23796 36722
rect 23848 36576 23900 36582
rect 23848 36518 23900 36524
rect 23756 35760 23808 35766
rect 23756 35702 23808 35708
rect 23664 35624 23716 35630
rect 23664 35566 23716 35572
rect 23860 35494 23888 36518
rect 24032 36100 24084 36106
rect 24032 36042 24084 36048
rect 23848 35488 23900 35494
rect 23848 35430 23900 35436
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23664 35216 23716 35222
rect 23664 35158 23716 35164
rect 23676 33522 23704 35158
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 23860 34649 23888 34682
rect 23846 34640 23902 34649
rect 23846 34575 23902 34584
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23676 30190 23704 32846
rect 23952 31754 23980 35430
rect 24044 32434 24072 36042
rect 24136 35698 24164 41618
rect 24228 41414 24256 45526
rect 24320 42770 24348 53042
rect 24308 42764 24360 42770
rect 24308 42706 24360 42712
rect 24228 41386 24348 41414
rect 24320 37874 24348 41386
rect 24308 37868 24360 37874
rect 24308 37810 24360 37816
rect 24320 36786 24348 37810
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24124 35692 24176 35698
rect 24124 35634 24176 35640
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 23860 31726 23980 31754
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 23308 22574 23336 23190
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23308 10062 23336 22510
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23400 19446 23428 20946
rect 23584 20466 23612 22170
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23400 18834 23428 19382
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23400 16658 23428 18770
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23492 15638 23520 20334
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23570 14920 23626 14929
rect 23570 14855 23626 14864
rect 23584 14822 23612 14855
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23400 12646 23428 14758
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23492 12306 23520 12650
rect 23570 12472 23626 12481
rect 23570 12407 23626 12416
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23400 9908 23428 10066
rect 23308 9880 23428 9908
rect 23308 8809 23336 9880
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23294 8800 23350 8809
rect 23294 8735 23350 8744
rect 23294 8392 23350 8401
rect 23294 8327 23350 8336
rect 23308 6458 23336 8327
rect 23400 6730 23428 9454
rect 23492 6905 23520 10474
rect 23478 6896 23534 6905
rect 23478 6831 23534 6840
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23294 6352 23350 6361
rect 23204 6316 23256 6322
rect 23294 6287 23296 6296
rect 23204 6258 23256 6264
rect 23348 6287 23350 6296
rect 23296 6258 23348 6264
rect 23216 5846 23244 6258
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 23110 4312 23166 4321
rect 23110 4247 23166 4256
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 23124 3505 23152 4247
rect 23308 4146 23336 6258
rect 23400 6089 23428 6666
rect 23386 6080 23442 6089
rect 23386 6015 23442 6024
rect 23492 5642 23520 6831
rect 23584 5914 23612 12407
rect 23676 10985 23704 30126
rect 23860 29646 23888 31726
rect 23940 30320 23992 30326
rect 23940 30262 23992 30268
rect 24032 30320 24084 30326
rect 24032 30262 24084 30268
rect 23952 30161 23980 30262
rect 23938 30152 23994 30161
rect 23938 30087 23994 30096
rect 24044 29866 24072 30262
rect 23952 29838 24072 29866
rect 23952 29782 23980 29838
rect 23940 29776 23992 29782
rect 23940 29718 23992 29724
rect 24032 29776 24084 29782
rect 24032 29718 24084 29724
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23860 23497 23888 29582
rect 24044 29102 24072 29718
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 24136 27334 24164 35634
rect 24216 30388 24268 30394
rect 24216 30330 24268 30336
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 23846 23488 23902 23497
rect 23846 23423 23902 23432
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23940 21956 23992 21962
rect 23940 21898 23992 21904
rect 23768 21350 23796 21898
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23768 19281 23796 19450
rect 23754 19272 23810 19281
rect 23754 19207 23810 19216
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23768 17542 23796 18022
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23768 13569 23796 17002
rect 23754 13560 23810 13569
rect 23754 13495 23810 13504
rect 23846 11248 23902 11257
rect 23846 11183 23902 11192
rect 23662 10976 23718 10985
rect 23662 10911 23718 10920
rect 23664 10056 23716 10062
rect 23662 10024 23664 10033
rect 23716 10024 23718 10033
rect 23662 9959 23718 9968
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23676 9353 23704 9386
rect 23662 9344 23718 9353
rect 23662 9279 23718 9288
rect 23768 8673 23796 9930
rect 23754 8664 23810 8673
rect 23754 8599 23810 8608
rect 23754 8528 23810 8537
rect 23754 8463 23756 8472
rect 23808 8463 23810 8472
rect 23756 8434 23808 8440
rect 23768 8022 23796 8434
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23756 6928 23808 6934
rect 23756 6870 23808 6876
rect 23768 6798 23796 6870
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23756 6656 23808 6662
rect 23676 6616 23756 6644
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23676 5545 23704 6616
rect 23756 6598 23808 6604
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23662 5536 23718 5545
rect 23662 5471 23718 5480
rect 23768 5370 23796 6054
rect 23860 5846 23888 11183
rect 23952 9178 23980 21898
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24136 20534 24164 21490
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24044 18154 24072 18294
rect 24032 18148 24084 18154
rect 24032 18090 24084 18096
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 24044 16590 24072 17546
rect 24136 17338 24164 19994
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24228 17218 24256 30330
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24320 29238 24348 29990
rect 24412 29578 24440 60454
rect 24504 34542 24532 60522
rect 24688 60466 24716 60658
rect 24596 60438 24716 60466
rect 24596 59702 24624 60438
rect 24768 60104 24820 60110
rect 24768 60046 24820 60052
rect 24674 59936 24730 59945
rect 24674 59871 24730 59880
rect 24584 59696 24636 59702
rect 24584 59638 24636 59644
rect 24688 59616 24716 59871
rect 24780 59786 24808 60046
rect 24964 60042 24992 61610
rect 25148 61198 25176 63200
rect 25884 61198 25912 63200
rect 26620 61198 26648 63200
rect 25136 61192 25188 61198
rect 25136 61134 25188 61140
rect 25872 61192 25924 61198
rect 25872 61134 25924 61140
rect 26608 61192 26660 61198
rect 26608 61134 26660 61140
rect 26884 61124 26936 61130
rect 26884 61066 26936 61072
rect 25228 60580 25280 60586
rect 25228 60522 25280 60528
rect 25240 60110 25268 60522
rect 25964 60308 26016 60314
rect 25964 60250 26016 60256
rect 26792 60308 26844 60314
rect 26792 60250 26844 60256
rect 25872 60240 25924 60246
rect 25872 60182 25924 60188
rect 25136 60104 25188 60110
rect 25136 60046 25188 60052
rect 25228 60104 25280 60110
rect 25228 60046 25280 60052
rect 25504 60104 25556 60110
rect 25504 60046 25556 60052
rect 24952 60036 25004 60042
rect 24952 59978 25004 59984
rect 24780 59758 24900 59786
rect 24768 59628 24820 59634
rect 24688 59588 24768 59616
rect 24768 59570 24820 59576
rect 24872 59378 24900 59758
rect 25148 59498 25176 60046
rect 25516 59770 25544 60046
rect 25884 59974 25912 60182
rect 25976 60110 26004 60250
rect 26056 60240 26108 60246
rect 26056 60182 26108 60188
rect 25964 60104 26016 60110
rect 25964 60046 26016 60052
rect 25872 59968 25924 59974
rect 25872 59910 25924 59916
rect 25870 59800 25926 59809
rect 25504 59764 25556 59770
rect 25870 59735 25926 59744
rect 25504 59706 25556 59712
rect 25884 59702 25912 59735
rect 25872 59696 25924 59702
rect 25872 59638 25924 59644
rect 25780 59628 25832 59634
rect 25700 59588 25780 59616
rect 25136 59492 25188 59498
rect 25136 59434 25188 59440
rect 25596 59492 25648 59498
rect 25700 59480 25728 59588
rect 25780 59570 25832 59576
rect 25648 59452 25728 59480
rect 25778 59528 25834 59537
rect 25778 59463 25780 59472
rect 25596 59434 25648 59440
rect 24780 59350 24900 59378
rect 24780 48278 24808 59350
rect 25700 56778 25728 59452
rect 25832 59463 25834 59472
rect 25780 59434 25832 59440
rect 25964 59424 26016 59430
rect 25964 59366 26016 59372
rect 25688 56772 25740 56778
rect 25688 56714 25740 56720
rect 25700 51074 25728 56714
rect 25516 51046 25728 51074
rect 24768 48272 24820 48278
rect 24768 48214 24820 48220
rect 25412 48272 25464 48278
rect 25412 48214 25464 48220
rect 24860 46980 24912 46986
rect 24860 46922 24912 46928
rect 24582 41576 24638 41585
rect 24582 41511 24584 41520
rect 24636 41511 24638 41520
rect 24584 41482 24636 41488
rect 24768 35216 24820 35222
rect 24768 35158 24820 35164
rect 24780 35086 24808 35158
rect 24768 35080 24820 35086
rect 24768 35022 24820 35028
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24676 34536 24728 34542
rect 24676 34478 24728 34484
rect 24688 30326 24716 34478
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24504 29782 24532 30194
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24400 29572 24452 29578
rect 24400 29514 24452 29520
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 24400 23248 24452 23254
rect 24400 23190 24452 23196
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24320 18970 24348 19178
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24412 18426 24440 23190
rect 24504 18442 24532 28902
rect 24596 28422 24624 29582
rect 24688 29578 24716 30262
rect 24780 30054 24808 33458
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24872 29646 24900 46922
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 31822 25360 32166
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25134 30288 25190 30297
rect 25134 30223 25136 30232
rect 25188 30223 25190 30232
rect 25136 30194 25188 30200
rect 25136 30048 25188 30054
rect 25136 29990 25188 29996
rect 25148 29714 25176 29990
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 25240 29458 25268 31282
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 25332 30326 25360 30874
rect 25320 30320 25372 30326
rect 25320 30262 25372 30268
rect 25332 29578 25360 30262
rect 25320 29572 25372 29578
rect 25320 29514 25372 29520
rect 25148 29238 25176 29446
rect 25240 29430 25360 29458
rect 25136 29232 25188 29238
rect 25136 29174 25188 29180
rect 25332 29102 25360 29430
rect 25424 29102 25452 48214
rect 25516 31958 25544 51046
rect 25594 37904 25650 37913
rect 25594 37839 25650 37848
rect 25504 31952 25556 31958
rect 25504 31894 25556 31900
rect 25608 31414 25636 37839
rect 25976 34610 26004 59366
rect 26068 54738 26096 60182
rect 26424 60104 26476 60110
rect 26424 60046 26476 60052
rect 26436 59974 26464 60046
rect 26240 59968 26292 59974
rect 26240 59910 26292 59916
rect 26424 59968 26476 59974
rect 26424 59910 26476 59916
rect 26252 59634 26280 59910
rect 26240 59628 26292 59634
rect 26240 59570 26292 59576
rect 26148 59560 26200 59566
rect 26148 59502 26200 59508
rect 26056 54732 26108 54738
rect 26056 54674 26108 54680
rect 26160 51074 26188 59502
rect 26332 51808 26384 51814
rect 26332 51750 26384 51756
rect 26068 51046 26188 51074
rect 26068 41414 26096 51046
rect 26068 41386 26188 41414
rect 26056 38888 26108 38894
rect 26056 38830 26108 38836
rect 26068 37913 26096 38830
rect 26054 37904 26110 37913
rect 26054 37839 26110 37848
rect 26160 35834 26188 41386
rect 26148 35828 26200 35834
rect 26148 35770 26200 35776
rect 26160 35018 26188 35770
rect 26148 35012 26200 35018
rect 26148 34954 26200 34960
rect 26344 34678 26372 51750
rect 26436 47705 26464 59910
rect 26804 59770 26832 60250
rect 26896 60110 26924 61066
rect 27344 61056 27396 61062
rect 27344 60998 27396 61004
rect 27160 60852 27212 60858
rect 27160 60794 27212 60800
rect 26976 60172 27028 60178
rect 26976 60114 27028 60120
rect 26884 60104 26936 60110
rect 26884 60046 26936 60052
rect 26792 59764 26844 59770
rect 26792 59706 26844 59712
rect 26988 59702 27016 60114
rect 27172 60110 27200 60794
rect 27356 60734 27384 60998
rect 27540 60790 27568 63294
rect 28078 63200 28134 64000
rect 28814 63322 28870 64000
rect 29550 63322 29606 64000
rect 28814 63294 28948 63322
rect 28814 63200 28870 63294
rect 28092 61198 28120 63200
rect 28356 61600 28408 61606
rect 28356 61542 28408 61548
rect 28264 61260 28316 61266
rect 28264 61202 28316 61208
rect 28080 61192 28132 61198
rect 28080 61134 28132 61140
rect 27528 60784 27580 60790
rect 27356 60706 27476 60734
rect 27528 60726 27580 60732
rect 27160 60104 27212 60110
rect 27160 60046 27212 60052
rect 27252 60104 27304 60110
rect 27252 60046 27304 60052
rect 27264 59945 27292 60046
rect 27250 59936 27306 59945
rect 27250 59871 27306 59880
rect 26976 59696 27028 59702
rect 26976 59638 27028 59644
rect 26884 59084 26936 59090
rect 26884 59026 26936 59032
rect 26896 58857 26924 59026
rect 26882 58848 26938 58857
rect 26882 58783 26938 58792
rect 26976 57044 27028 57050
rect 26976 56986 27028 56992
rect 26608 55684 26660 55690
rect 26608 55626 26660 55632
rect 26422 47696 26478 47705
rect 26422 47631 26478 47640
rect 26620 40118 26648 55626
rect 26608 40112 26660 40118
rect 26608 40054 26660 40060
rect 26332 34672 26384 34678
rect 26332 34614 26384 34620
rect 26884 34672 26936 34678
rect 26884 34614 26936 34620
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 26148 34604 26200 34610
rect 26148 34546 26200 34552
rect 26056 34468 26108 34474
rect 26056 34410 26108 34416
rect 26068 32026 26096 34410
rect 26160 32434 26188 34546
rect 26608 34400 26660 34406
rect 26608 34342 26660 34348
rect 26620 33046 26648 34342
rect 26608 33040 26660 33046
rect 26608 32982 26660 32988
rect 26700 32904 26752 32910
rect 26700 32846 26752 32852
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 25964 31952 26016 31958
rect 25964 31894 26016 31900
rect 25780 31748 25832 31754
rect 25780 31690 25832 31696
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25608 30938 25636 31350
rect 25792 31346 25820 31690
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25596 30932 25648 30938
rect 25596 30874 25648 30880
rect 25686 30288 25742 30297
rect 25686 30223 25742 30232
rect 25700 30190 25728 30223
rect 25688 30184 25740 30190
rect 25688 30126 25740 30132
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 29850 25912 29990
rect 25976 29850 26004 31894
rect 26068 31822 26096 31962
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26712 31482 26740 32846
rect 26700 31476 26752 31482
rect 26700 31418 26752 31424
rect 26330 30152 26386 30161
rect 26330 30087 26332 30096
rect 26384 30087 26386 30096
rect 26332 30058 26384 30064
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 25964 29844 26016 29850
rect 25964 29786 26016 29792
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 25596 29504 25648 29510
rect 25596 29446 25648 29452
rect 25608 29170 25636 29446
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25320 29096 25372 29102
rect 25320 29038 25372 29044
rect 25412 29096 25464 29102
rect 25412 29038 25464 29044
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22030 24624 22918
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24688 21010 24716 23054
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24596 20262 24624 20402
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24596 20058 24624 20198
rect 24780 20074 24808 20198
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24688 20046 24808 20074
rect 24688 19854 24716 20046
rect 24766 19952 24822 19961
rect 24766 19887 24822 19896
rect 24860 19916 24912 19922
rect 24780 19854 24808 19887
rect 24860 19858 24912 19864
rect 24676 19848 24728 19854
rect 24582 19816 24638 19825
rect 24676 19790 24728 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24582 19751 24584 19760
rect 24636 19751 24638 19760
rect 24584 19722 24636 19728
rect 24596 18630 24624 19722
rect 24780 19417 24808 19790
rect 24766 19408 24822 19417
rect 24766 19343 24822 19352
rect 24872 18766 24900 19858
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24504 18414 24808 18442
rect 24320 18329 24348 18362
rect 24306 18320 24362 18329
rect 24306 18255 24362 18264
rect 24504 18034 24532 18414
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24412 18006 24532 18034
rect 24412 17814 24440 18006
rect 24400 17808 24452 17814
rect 24584 17808 24636 17814
rect 24400 17750 24452 17756
rect 24582 17776 24584 17785
rect 24636 17776 24638 17785
rect 24492 17740 24544 17746
rect 24582 17711 24638 17720
rect 24492 17682 24544 17688
rect 24504 17270 24532 17682
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24492 17264 24544 17270
rect 24228 17190 24440 17218
rect 24492 17206 24544 17212
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 14385 24072 15846
rect 24030 14376 24086 14385
rect 24030 14311 24086 14320
rect 24044 12889 24072 14311
rect 24136 14113 24164 16934
rect 24216 15972 24268 15978
rect 24216 15914 24268 15920
rect 24122 14104 24178 14113
rect 24122 14039 24178 14048
rect 24030 12880 24086 12889
rect 24030 12815 24032 12824
rect 24084 12815 24086 12824
rect 24032 12786 24084 12792
rect 24044 11898 24072 12786
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24032 10736 24084 10742
rect 24030 10704 24032 10713
rect 24084 10704 24086 10713
rect 24030 10639 24086 10648
rect 24136 10305 24164 14039
rect 24228 13002 24256 15914
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24320 13938 24348 14486
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24320 13190 24348 13874
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24228 12974 24348 13002
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24228 11898 24256 12718
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24320 11762 24348 12974
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24320 11626 24348 11698
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 24122 10296 24178 10305
rect 24032 10260 24084 10266
rect 24412 10266 24440 17190
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24504 15910 24532 16186
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24596 14618 24624 17614
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24596 12238 24624 12378
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 12073 24624 12174
rect 24582 12064 24638 12073
rect 24582 11999 24638 12008
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24504 11286 24532 11698
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24492 11144 24544 11150
rect 24544 11092 24624 11098
rect 24492 11086 24624 11092
rect 24504 11070 24624 11086
rect 24122 10231 24178 10240
rect 24400 10260 24452 10266
rect 24032 10202 24084 10208
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23952 6798 23980 8910
rect 24044 8430 24072 10202
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24136 6798 24164 10231
rect 24400 10202 24452 10208
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24228 8809 24256 9522
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24214 8800 24270 8809
rect 24214 8735 24270 8744
rect 24398 8528 24454 8537
rect 24398 8463 24454 8472
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7206 24256 7686
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24216 6996 24268 7002
rect 24216 6938 24268 6944
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 23952 6644 23980 6734
rect 23952 6616 24164 6644
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 23492 4758 23520 5063
rect 23480 4752 23532 4758
rect 23480 4694 23532 4700
rect 23768 4690 23796 5306
rect 24032 5296 24084 5302
rect 24032 5238 24084 5244
rect 24044 5030 24072 5238
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23216 3534 23244 3878
rect 23400 3670 23428 4082
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23204 3528 23256 3534
rect 23110 3496 23166 3505
rect 23204 3470 23256 3476
rect 23110 3431 23166 3440
rect 23124 3398 23152 3431
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23112 3188 23164 3194
rect 23216 3176 23244 3334
rect 23164 3148 23244 3176
rect 23112 3130 23164 3136
rect 22926 3088 22982 3097
rect 22926 3023 22928 3032
rect 22980 3023 22982 3032
rect 22928 2994 22980 3000
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22756 882 22784 2858
rect 23124 2825 23152 3130
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23110 2816 23166 2825
rect 23110 2751 23166 2760
rect 23018 2680 23074 2689
rect 23018 2615 23074 2624
rect 23032 2582 23060 2615
rect 23124 2582 23152 2751
rect 23308 2650 23336 2994
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23020 2576 23072 2582
rect 23020 2518 23072 2524
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 23204 2440 23256 2446
rect 23400 2428 23428 3606
rect 23584 3194 23612 4422
rect 23952 3398 23980 4626
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23938 3224 23994 3233
rect 23572 3188 23624 3194
rect 23938 3159 23994 3168
rect 23572 3130 23624 3136
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23256 2400 23428 2428
rect 23204 2382 23256 2388
rect 23572 2372 23624 2378
rect 23572 2314 23624 2320
rect 23480 2304 23532 2310
rect 23400 2264 23480 2292
rect 22928 1964 22980 1970
rect 22928 1906 22980 1912
rect 22744 876 22796 882
rect 22744 818 22796 824
rect 22940 800 22968 1906
rect 23204 1488 23256 1494
rect 23204 1430 23256 1436
rect 23216 800 23244 1430
rect 23400 950 23428 2264
rect 23480 2246 23532 2252
rect 23480 1760 23532 1766
rect 23480 1702 23532 1708
rect 23388 944 23440 950
rect 23388 886 23440 892
rect 23492 800 23520 1702
rect 23584 1290 23612 2314
rect 23572 1284 23624 1290
rect 23572 1226 23624 1232
rect 23768 800 23796 2926
rect 23952 1578 23980 3159
rect 24044 3058 24072 4966
rect 24136 3233 24164 6616
rect 24228 6254 24256 6938
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24412 5710 24440 8463
rect 24504 5953 24532 9318
rect 24596 8974 24624 11070
rect 24688 10266 24716 18090
rect 24780 17678 24808 18414
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24872 17490 24900 17614
rect 24780 17462 24900 17490
rect 24780 16998 24808 17462
rect 24964 17218 24992 24210
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19922 25176 20334
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25240 19961 25268 19994
rect 25226 19952 25282 19961
rect 25136 19916 25188 19922
rect 25226 19887 25282 19896
rect 25136 19858 25188 19864
rect 24872 17190 24992 17218
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24780 14414 24808 15574
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24780 10470 24808 11494
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24688 10033 24716 10066
rect 24674 10024 24730 10033
rect 24674 9959 24730 9968
rect 24674 9888 24730 9897
rect 24674 9823 24730 9832
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24688 7886 24716 9823
rect 24780 8974 24808 10406
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24584 7812 24636 7818
rect 24584 7754 24636 7760
rect 24596 7342 24624 7754
rect 24780 7426 24808 8910
rect 24688 7398 24808 7426
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24688 6746 24716 7398
rect 24872 6798 24900 17190
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 25056 16250 25084 16458
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25056 15366 25084 15438
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25148 15162 25176 15506
rect 25240 15366 25268 15574
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 13734 25268 13874
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24964 10606 24992 11018
rect 25056 10674 25084 12854
rect 25148 12238 25176 13262
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 24964 9926 24992 10202
rect 25148 10130 25176 12174
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25240 10044 25268 11086
rect 25332 10266 25360 29038
rect 25412 27328 25464 27334
rect 25412 27270 25464 27276
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25320 10056 25372 10062
rect 25240 10016 25320 10044
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 9738 25084 9862
rect 24964 9722 25084 9738
rect 24952 9716 25084 9722
rect 25004 9710 25084 9716
rect 24952 9658 25004 9664
rect 25044 9648 25096 9654
rect 25096 9608 25176 9636
rect 25044 9590 25096 9596
rect 25148 9518 25176 9608
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24964 8634 24992 9114
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25056 8430 25084 9454
rect 25148 9382 25176 9454
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25240 9042 25268 10016
rect 25320 9998 25372 10004
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24964 7342 24992 8366
rect 25056 7834 25084 8366
rect 25134 7984 25190 7993
rect 25240 7954 25268 8978
rect 25424 8634 25452 27270
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25516 19514 25544 22986
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25516 14890 25544 15302
rect 25608 14958 25636 21490
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25700 19825 25728 19858
rect 25686 19816 25742 19825
rect 25686 19751 25742 19760
rect 25792 17338 25820 22578
rect 25872 22500 25924 22506
rect 25872 22442 25924 22448
rect 25884 21690 25912 22442
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25700 16998 25728 17206
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25884 15366 25912 18294
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25504 14884 25556 14890
rect 25504 14826 25556 14832
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25504 14408 25556 14414
rect 25502 14376 25504 14385
rect 25556 14376 25558 14385
rect 25608 14346 25636 14554
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25502 14311 25558 14320
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 25516 13530 25544 13670
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25792 12434 25820 14447
rect 25700 12406 25820 12434
rect 25594 11520 25650 11529
rect 25594 11455 25650 11464
rect 25608 11218 25636 11455
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25134 7919 25136 7928
rect 25188 7919 25190 7928
rect 25228 7948 25280 7954
rect 25136 7890 25188 7896
rect 25228 7890 25280 7896
rect 25056 7806 25176 7834
rect 25148 7750 25176 7806
rect 25516 7750 25544 10202
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25608 8090 25636 9522
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 24964 6934 24992 7278
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24596 6718 24716 6746
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24490 5944 24546 5953
rect 24490 5879 24546 5888
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24320 5545 24348 5646
rect 24306 5536 24362 5545
rect 24306 5471 24362 5480
rect 24504 5234 24532 5879
rect 24596 5692 24624 6718
rect 24950 6624 25006 6633
rect 24950 6559 25006 6568
rect 24964 6322 24992 6559
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 25056 6186 25084 7142
rect 25148 6882 25176 7686
rect 25228 7268 25280 7274
rect 25228 7210 25280 7216
rect 25240 7002 25268 7210
rect 25228 6996 25280 7002
rect 25228 6938 25280 6944
rect 25148 6854 25268 6882
rect 25044 6180 25096 6186
rect 25044 6122 25096 6128
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 24676 5704 24728 5710
rect 24596 5664 24676 5692
rect 24676 5646 24728 5652
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24872 5370 24900 5578
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24412 4282 24440 5102
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 24584 4548 24636 4554
rect 24584 4490 24636 4496
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24122 3224 24178 3233
rect 24122 3159 24178 3168
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24228 1766 24256 4014
rect 24216 1760 24268 1766
rect 24216 1702 24268 1708
rect 24320 1680 24348 4150
rect 24398 3904 24454 3913
rect 24398 3839 24454 3848
rect 24412 3738 24440 3839
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24398 3632 24454 3641
rect 24398 3567 24454 3576
rect 24412 2922 24440 3567
rect 24400 2916 24452 2922
rect 24400 2858 24452 2864
rect 24320 1652 24440 1680
rect 23952 1550 24072 1578
rect 24044 800 24072 1550
rect 24412 1018 24440 1652
rect 24400 1012 24452 1018
rect 24400 954 24452 960
rect 24228 836 24348 864
rect 21640 672 21692 678
rect 21640 614 21692 620
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24228 542 24256 836
rect 24320 800 24348 836
rect 24504 814 24532 4490
rect 24596 3738 24624 4490
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24688 3602 24716 5102
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24780 3074 24808 4558
rect 24872 4214 24900 4626
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24872 4078 24900 4150
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24872 3534 24900 3674
rect 24964 3641 24992 5238
rect 25148 5234 25176 5714
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25148 4690 25176 5170
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 4146 25176 4626
rect 25136 4140 25188 4146
rect 25136 4082 25188 4088
rect 25044 4004 25096 4010
rect 25044 3946 25096 3952
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24780 3046 24992 3074
rect 24964 2774 24992 3046
rect 25056 2836 25084 3946
rect 25148 3641 25176 4082
rect 25134 3632 25190 3641
rect 25134 3567 25190 3576
rect 25240 3398 25268 6854
rect 25516 6186 25544 7686
rect 25608 6866 25636 7890
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 25608 5914 25636 6802
rect 25700 6730 25728 12406
rect 25778 12064 25834 12073
rect 25778 11999 25834 12008
rect 25792 9489 25820 11999
rect 25976 10985 26004 29582
rect 26160 25702 26188 29582
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 26056 22432 26108 22438
rect 26056 22374 26108 22380
rect 26068 20942 26096 22374
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26252 20330 26280 21422
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26068 18970 26096 19790
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 26068 18630 26096 18770
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26056 18216 26108 18222
rect 26054 18184 26056 18193
rect 26108 18184 26110 18193
rect 26160 18154 26188 19314
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26054 18119 26110 18128
rect 26148 18148 26200 18154
rect 26148 18090 26200 18096
rect 26252 17678 26280 18566
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26344 17202 26372 26250
rect 26896 24857 26924 34614
rect 26988 32910 27016 56986
rect 27344 56296 27396 56302
rect 27344 56238 27396 56244
rect 27356 55758 27384 56238
rect 27344 55752 27396 55758
rect 27344 55694 27396 55700
rect 27448 53106 27476 60706
rect 28080 60512 28132 60518
rect 28080 60454 28132 60460
rect 28172 60512 28224 60518
rect 28172 60454 28224 60460
rect 28092 60110 28120 60454
rect 28184 60178 28212 60454
rect 28172 60172 28224 60178
rect 28172 60114 28224 60120
rect 27988 60104 28040 60110
rect 27988 60046 28040 60052
rect 28080 60104 28132 60110
rect 28080 60046 28132 60052
rect 27528 59968 27580 59974
rect 27528 59910 27580 59916
rect 27540 55826 27568 59910
rect 28000 59430 28028 60046
rect 27988 59424 28040 59430
rect 27988 59366 28040 59372
rect 27620 56704 27672 56710
rect 27620 56646 27672 56652
rect 27632 56438 27660 56646
rect 27620 56432 27672 56438
rect 27620 56374 27672 56380
rect 27528 55820 27580 55826
rect 27528 55762 27580 55768
rect 27528 54528 27580 54534
rect 27528 54470 27580 54476
rect 27540 53174 27568 54470
rect 27528 53168 27580 53174
rect 27528 53110 27580 53116
rect 27436 53100 27488 53106
rect 27436 53042 27488 53048
rect 27436 33448 27488 33454
rect 27436 33390 27488 33396
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 26976 29096 27028 29102
rect 26976 29038 27028 29044
rect 26882 24848 26938 24857
rect 26882 24783 26938 24792
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 26516 22228 26568 22234
rect 26516 22170 26568 22176
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26436 20602 26464 22034
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26436 18358 26464 18838
rect 26424 18352 26476 18358
rect 26424 18294 26476 18300
rect 26422 17776 26478 17785
rect 26422 17711 26478 17720
rect 26436 17678 26464 17711
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26056 16720 26108 16726
rect 26056 16662 26108 16668
rect 26068 15570 26096 16662
rect 26528 15638 26556 22170
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 26620 14550 26648 23054
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26712 20466 26740 21286
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 17882 26832 19654
rect 26896 18766 26924 20198
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26896 17882 26924 18022
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26712 16726 26740 17070
rect 26700 16720 26752 16726
rect 26700 16662 26752 16668
rect 26896 16590 26924 17478
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 26608 14544 26660 14550
rect 26608 14486 26660 14492
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26068 12918 26096 13330
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26148 13184 26200 13190
rect 26528 13161 26556 13262
rect 26148 13126 26200 13132
rect 26514 13152 26570 13161
rect 26056 12912 26108 12918
rect 26056 12854 26108 12860
rect 26160 11830 26188 13126
rect 26514 13087 26570 13096
rect 26528 12918 26556 13087
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26148 11824 26200 11830
rect 26148 11766 26200 11772
rect 25962 10976 26018 10985
rect 25962 10911 26018 10920
rect 25872 9648 25924 9654
rect 25976 9636 26004 10911
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 25924 9608 26004 9636
rect 25872 9590 25924 9596
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 25872 9512 25924 9518
rect 25778 9480 25834 9489
rect 25872 9454 25924 9460
rect 25778 9415 25834 9424
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25792 8498 25820 9318
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25884 8430 25912 9454
rect 26068 9217 26096 9522
rect 26148 9444 26200 9450
rect 26148 9386 26200 9392
rect 26054 9208 26110 9217
rect 26054 9143 26110 9152
rect 26160 8498 26188 9386
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 26344 8362 26372 10542
rect 26436 9761 26464 12786
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26422 9752 26478 9761
rect 26422 9687 26478 9696
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26436 9042 26464 9454
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 25792 7426 25820 8026
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 25884 7546 25912 7754
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25792 7398 25912 7426
rect 25780 7336 25832 7342
rect 25778 7304 25780 7313
rect 25832 7304 25834 7313
rect 25778 7239 25834 7248
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25608 5545 25636 5578
rect 25594 5536 25650 5545
rect 25594 5471 25650 5480
rect 25792 4146 25820 7239
rect 25884 5030 25912 7398
rect 26068 6730 26096 8026
rect 26528 7546 26556 11834
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26620 9722 26648 10950
rect 26712 10849 26740 13262
rect 26698 10840 26754 10849
rect 26698 10775 26754 10784
rect 26698 10024 26754 10033
rect 26698 9959 26754 9968
rect 26712 9722 26740 9959
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26620 9178 26648 9658
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 7546 26740 8774
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 26804 6458 26832 13942
rect 26792 6452 26844 6458
rect 26792 6394 26844 6400
rect 26608 6180 26660 6186
rect 26608 6122 26660 6128
rect 26620 5846 26648 6122
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25780 4140 25832 4146
rect 26160 4128 26188 5510
rect 26422 4176 26478 4185
rect 26160 4100 26280 4128
rect 26422 4111 26478 4120
rect 25780 4082 25832 4088
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25424 3194 25452 4082
rect 25502 3768 25558 3777
rect 25502 3703 25558 3712
rect 25516 3194 25544 3703
rect 25778 3632 25834 3641
rect 25778 3567 25780 3576
rect 25832 3567 25834 3576
rect 25780 3538 25832 3544
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 25700 2990 25728 3470
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25688 2984 25740 2990
rect 25688 2926 25740 2932
rect 25136 2848 25188 2854
rect 25056 2808 25136 2836
rect 25136 2790 25188 2796
rect 24964 2746 25084 2774
rect 25056 2650 25084 2746
rect 25608 2666 25636 2926
rect 25516 2650 25636 2666
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 25504 2644 25636 2650
rect 25556 2638 25636 2644
rect 25504 2586 25556 2592
rect 24584 1828 24636 1834
rect 24584 1770 24636 1776
rect 24492 808 24544 814
rect 24216 536 24268 542
rect 24216 478 24268 484
rect 24306 0 24362 800
rect 24596 800 24624 1770
rect 24780 1086 24808 2586
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 25608 2310 25636 2518
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 25134 1864 25190 1873
rect 25134 1799 25190 1808
rect 24768 1080 24820 1086
rect 24768 1022 24820 1028
rect 24780 836 24900 864
rect 24492 750 24544 756
rect 24582 0 24638 800
rect 24674 776 24730 785
rect 24780 762 24808 836
rect 24872 800 24900 836
rect 25148 800 25176 1799
rect 25410 1592 25466 1601
rect 25410 1527 25466 1536
rect 25424 800 25452 1527
rect 25686 1456 25742 1465
rect 25686 1391 25742 1400
rect 25700 800 25728 1391
rect 25884 836 26004 864
rect 24730 734 24808 762
rect 24674 711 24730 720
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25884 762 25912 836
rect 25976 800 26004 836
rect 26252 800 26280 4100
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26344 3126 26372 3334
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 26344 2378 26372 2450
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 26436 1714 26464 4111
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26528 1834 26556 2246
rect 26516 1828 26568 1834
rect 26516 1770 26568 1776
rect 26436 1686 26556 1714
rect 26528 800 26556 1686
rect 26804 800 26832 2790
rect 26896 2514 26924 16186
rect 26988 12986 27016 29038
rect 27172 27033 27200 32710
rect 27158 27024 27214 27033
rect 27158 26959 27214 26968
rect 27448 22166 27476 33390
rect 27712 31204 27764 31210
rect 27712 31146 27764 31152
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27632 22574 27660 23122
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27436 22160 27488 22166
rect 27436 22102 27488 22108
rect 27448 22001 27476 22102
rect 27434 21992 27490 22001
rect 27434 21927 27490 21936
rect 27540 21622 27568 22374
rect 27724 22094 27752 31146
rect 28276 31142 28304 61202
rect 28368 60518 28396 61542
rect 28448 61124 28500 61130
rect 28448 61066 28500 61072
rect 28356 60512 28408 60518
rect 28356 60454 28408 60460
rect 28356 56976 28408 56982
rect 28356 56918 28408 56924
rect 28368 33114 28396 56918
rect 28356 33108 28408 33114
rect 28356 33050 28408 33056
rect 28264 31136 28316 31142
rect 28264 31078 28316 31084
rect 28460 22817 28488 61066
rect 28920 61044 28948 63294
rect 29550 63294 29868 63322
rect 29550 63200 29606 63294
rect 29840 61198 29868 63294
rect 30286 63200 30342 64000
rect 31022 63322 31078 64000
rect 31022 63294 31248 63322
rect 31022 63200 31078 63294
rect 29828 61192 29880 61198
rect 29828 61134 29880 61140
rect 29920 61056 29972 61062
rect 28920 61016 29040 61044
rect 29012 60790 29040 61016
rect 29920 60998 29972 61004
rect 29000 60784 29052 60790
rect 29000 60726 29052 60732
rect 29092 60512 29144 60518
rect 29092 60454 29144 60460
rect 28724 60240 28776 60246
rect 28724 60182 28776 60188
rect 28816 60240 28868 60246
rect 28816 60182 28868 60188
rect 28540 60172 28592 60178
rect 28540 60114 28592 60120
rect 28552 60081 28580 60114
rect 28736 60110 28764 60182
rect 28724 60104 28776 60110
rect 28538 60072 28594 60081
rect 28724 60046 28776 60052
rect 28828 60042 28856 60182
rect 29000 60104 29052 60110
rect 28998 60072 29000 60081
rect 29052 60072 29054 60081
rect 28538 60007 28594 60016
rect 28816 60036 28868 60042
rect 29104 60042 29132 60454
rect 29734 60344 29790 60353
rect 29734 60279 29736 60288
rect 29788 60279 29790 60288
rect 29736 60250 29788 60256
rect 29642 60208 29698 60217
rect 29642 60143 29644 60152
rect 29696 60143 29698 60152
rect 29644 60114 29696 60120
rect 29184 60104 29236 60110
rect 29184 60046 29236 60052
rect 28998 60007 29054 60016
rect 29092 60036 29144 60042
rect 28816 59978 28868 59984
rect 29092 59978 29144 59984
rect 29196 59770 29224 60046
rect 29276 59968 29328 59974
rect 29276 59910 29328 59916
rect 29184 59764 29236 59770
rect 29184 59706 29236 59712
rect 29288 56370 29316 59910
rect 29828 59424 29880 59430
rect 29828 59366 29880 59372
rect 29644 57248 29696 57254
rect 29644 57190 29696 57196
rect 29656 56370 29684 57190
rect 29276 56364 29328 56370
rect 29276 56306 29328 56312
rect 29644 56364 29696 56370
rect 29644 56306 29696 56312
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 28446 22808 28502 22817
rect 28446 22743 28502 22752
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27632 22066 27752 22094
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27160 21072 27212 21078
rect 27160 21014 27212 21020
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 27080 17954 27108 18362
rect 27172 18290 27200 21014
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27080 17926 27200 17954
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 26988 12617 27016 12922
rect 26974 12608 27030 12617
rect 26974 12543 27030 12552
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26988 9110 27016 9454
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 26974 8664 27030 8673
rect 27080 8634 27108 17138
rect 27172 16114 27200 17926
rect 27264 16574 27292 20742
rect 27356 17202 27384 21082
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27448 19378 27476 20402
rect 27632 19718 27660 22066
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27724 21690 27752 21830
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27816 20262 27844 22646
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28460 22030 28488 22510
rect 27896 22024 27948 22030
rect 27896 21966 27948 21972
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 27908 20806 27936 21966
rect 28172 21684 28224 21690
rect 28172 21626 28224 21632
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27896 20324 27948 20330
rect 27896 20266 27948 20272
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27632 19446 27660 19654
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27620 19440 27672 19446
rect 27620 19382 27672 19388
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 27632 18970 27660 19178
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27528 18352 27580 18358
rect 27526 18320 27528 18329
rect 27580 18320 27582 18329
rect 27632 18290 27660 18634
rect 27526 18255 27582 18264
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27436 18216 27488 18222
rect 27434 18184 27436 18193
rect 27488 18184 27490 18193
rect 27434 18119 27490 18128
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 17354 27660 17478
rect 27448 17338 27660 17354
rect 27436 17332 27660 17338
rect 27488 17326 27660 17332
rect 27436 17274 27488 17280
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27632 16658 27660 17070
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27264 16546 27384 16574
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27160 15700 27212 15706
rect 27160 15642 27212 15648
rect 27172 15434 27200 15642
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27264 13841 27292 14962
rect 27356 14822 27384 16546
rect 27618 16416 27674 16425
rect 27618 16351 27674 16360
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27540 15366 27568 16118
rect 27632 15978 27660 16351
rect 27724 16182 27752 19450
rect 27816 18086 27844 20198
rect 27908 18426 27936 20266
rect 27988 19236 28040 19242
rect 27988 19178 28040 19184
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27908 18086 27936 18226
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27908 17882 27936 18022
rect 27896 17876 27948 17882
rect 27896 17818 27948 17824
rect 27894 17776 27950 17785
rect 27894 17711 27896 17720
rect 27948 17711 27950 17720
rect 27896 17682 27948 17688
rect 28000 16250 28028 19178
rect 28080 19168 28132 19174
rect 28080 19110 28132 19116
rect 27988 16244 28040 16250
rect 27988 16186 28040 16192
rect 27712 16176 27764 16182
rect 27712 16118 27764 16124
rect 27620 15972 27672 15978
rect 27620 15914 27672 15920
rect 28092 15570 28120 19110
rect 28184 17542 28212 21626
rect 28460 21486 28488 21966
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28736 21554 28764 21830
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 28448 21480 28500 21486
rect 28816 21480 28868 21486
rect 28448 21422 28500 21428
rect 28736 21428 28816 21434
rect 28736 21422 28868 21428
rect 28540 21412 28592 21418
rect 28540 21354 28592 21360
rect 28736 21406 28856 21422
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28264 20800 28316 20806
rect 28264 20742 28316 20748
rect 28276 18290 28304 20742
rect 28460 20466 28488 21286
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28356 19236 28408 19242
rect 28356 19178 28408 19184
rect 28368 18902 28396 19178
rect 28356 18896 28408 18902
rect 28356 18838 28408 18844
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 28276 16454 28304 18226
rect 28356 18080 28408 18086
rect 28356 18022 28408 18028
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28080 15564 28132 15570
rect 28080 15506 28132 15512
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 28368 15162 28396 18022
rect 28460 17678 28488 18702
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 27250 13832 27306 13841
rect 27250 13767 27306 13776
rect 27528 13184 27580 13190
rect 27526 13152 27528 13161
rect 27580 13152 27582 13161
rect 27526 13087 27582 13096
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27620 12980 27672 12986
rect 27672 12940 27752 12968
rect 27620 12922 27672 12928
rect 27356 12850 27384 12922
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 27158 12608 27214 12617
rect 27158 12543 27214 12552
rect 27172 10470 27200 12543
rect 27356 12170 27384 12650
rect 27574 12640 27626 12646
rect 27448 12588 27574 12594
rect 27448 12582 27626 12588
rect 27448 12566 27614 12582
rect 27344 12164 27396 12170
rect 27344 12106 27396 12112
rect 27448 11898 27476 12566
rect 27724 12102 27752 12940
rect 27816 12918 27844 14758
rect 27988 13388 28040 13394
rect 27988 13330 28040 13336
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27816 12617 27844 12854
rect 27802 12608 27858 12617
rect 27802 12543 27858 12552
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27724 11898 27752 12038
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27344 11824 27396 11830
rect 27344 11766 27396 11772
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 26974 8599 26976 8608
rect 27028 8599 27030 8608
rect 27068 8628 27120 8634
rect 26976 8570 27028 8576
rect 27068 8570 27120 8576
rect 27172 8566 27200 8910
rect 27264 8566 27292 11290
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 27252 8560 27304 8566
rect 27252 8502 27304 8508
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 26988 6662 27016 7822
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27264 7478 27292 7686
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 27080 5914 27108 6734
rect 27356 6662 27384 11766
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27448 11354 27476 11494
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27632 11286 27660 11630
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27448 9450 27476 9522
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27448 9081 27476 9114
rect 27434 9072 27490 9081
rect 27434 9007 27490 9016
rect 27448 8498 27476 9007
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27540 8378 27568 11154
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27632 10305 27660 10610
rect 27618 10296 27674 10305
rect 27618 10231 27674 10240
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27632 9654 27660 9862
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 27448 8350 27568 8378
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27160 6248 27212 6254
rect 27448 6236 27476 8350
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27540 7342 27568 8230
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27540 7177 27568 7278
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 27526 7168 27582 7177
rect 27526 7103 27582 7112
rect 27526 6896 27582 6905
rect 27526 6831 27582 6840
rect 27540 6798 27568 6831
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27540 6322 27568 6598
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27212 6208 27476 6236
rect 27160 6190 27212 6196
rect 27342 5944 27398 5953
rect 27068 5908 27120 5914
rect 27342 5879 27344 5888
rect 27068 5850 27120 5856
rect 27396 5879 27398 5888
rect 27344 5850 27396 5856
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27540 4690 27568 4966
rect 27528 4684 27580 4690
rect 27448 4644 27528 4672
rect 26976 4480 27028 4486
rect 26976 4422 27028 4428
rect 26988 3466 27016 4422
rect 27448 4214 27476 4644
rect 27528 4626 27580 4632
rect 27632 4214 27660 7210
rect 27816 5642 27844 11630
rect 27894 9752 27950 9761
rect 27894 9687 27950 9696
rect 27908 6662 27936 9687
rect 28000 8430 28028 13330
rect 28092 11694 28120 14758
rect 28356 14476 28408 14482
rect 28356 14418 28408 14424
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28184 13530 28212 13738
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28184 12850 28212 13466
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28276 12850 28304 13126
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28368 12434 28396 14418
rect 28184 12406 28396 12434
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28184 10674 28212 12406
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28184 9110 28212 10610
rect 28276 9518 28304 11154
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28356 8900 28408 8906
rect 28356 8842 28408 8848
rect 28368 8634 28396 8842
rect 28460 8634 28488 15370
rect 28552 14498 28580 21354
rect 28736 20262 28764 21406
rect 29000 21344 29052 21350
rect 29000 21286 29052 21292
rect 28908 21004 28960 21010
rect 28908 20946 28960 20952
rect 28724 20256 28776 20262
rect 28724 20198 28776 20204
rect 28736 16658 28764 20198
rect 28816 19712 28868 19718
rect 28816 19654 28868 19660
rect 28828 17542 28856 19654
rect 28920 17678 28948 20946
rect 29012 20466 29040 21286
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17785 29040 18022
rect 29196 17882 29224 21490
rect 29274 19136 29330 19145
rect 29274 19071 29330 19080
rect 29184 17876 29236 17882
rect 29184 17818 29236 17824
rect 28998 17776 29054 17785
rect 28998 17711 29054 17720
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28552 14482 28672 14498
rect 28540 14476 28672 14482
rect 28592 14470 28672 14476
rect 28540 14418 28592 14424
rect 28538 14376 28594 14385
rect 28538 14311 28594 14320
rect 28552 11626 28580 14311
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28644 10130 28672 14470
rect 28736 12374 28764 16594
rect 28920 14822 28948 17614
rect 29000 17604 29052 17610
rect 29000 17546 29052 17552
rect 29012 15609 29040 17546
rect 29288 16250 29316 19071
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 16726 29408 17478
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29276 16244 29328 16250
rect 29276 16186 29328 16192
rect 28998 15600 29054 15609
rect 28998 15535 29054 15544
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 29012 15094 29040 15438
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 29380 14482 29408 16662
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29472 15366 29500 16050
rect 29460 15360 29512 15366
rect 29460 15302 29512 15308
rect 29368 14476 29420 14482
rect 29368 14418 29420 14424
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 28736 11218 28764 12310
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 29196 11898 29224 12038
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28724 10464 28776 10470
rect 28724 10406 28776 10412
rect 28814 10432 28870 10441
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 28632 9716 28684 9722
rect 28632 9658 28684 9664
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 27988 7744 28040 7750
rect 27986 7712 27988 7721
rect 28040 7712 28042 7721
rect 27986 7647 28042 7656
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 27988 6724 28040 6730
rect 27988 6666 28040 6672
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 28000 6458 28028 6666
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 27712 5636 27764 5642
rect 27712 5578 27764 5584
rect 27804 5636 27856 5642
rect 27804 5578 27856 5584
rect 28080 5636 28132 5642
rect 28080 5578 28132 5584
rect 27724 5370 27752 5578
rect 27802 5536 27858 5545
rect 27802 5471 27858 5480
rect 27712 5364 27764 5370
rect 27712 5306 27764 5312
rect 27816 4554 27844 5471
rect 28092 5370 28120 5578
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28080 5364 28132 5370
rect 28080 5306 28132 5312
rect 28184 5166 28212 5510
rect 28276 5234 28304 7142
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 28172 5160 28224 5166
rect 28172 5102 28224 5108
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27804 4548 27856 4554
rect 27804 4490 27856 4496
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27172 3534 27200 3878
rect 27264 3534 27292 4082
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27066 1728 27122 1737
rect 27066 1663 27122 1672
rect 27080 800 27108 1663
rect 27356 800 27384 3878
rect 27448 3194 27476 4150
rect 27908 4078 27936 5034
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 28000 4321 28028 4558
rect 27986 4312 28042 4321
rect 27986 4247 28042 4256
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27540 3074 27568 3402
rect 27632 3398 27660 4014
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 27448 3058 27568 3074
rect 27620 3120 27672 3126
rect 28092 3108 28120 4762
rect 28184 4593 28212 5102
rect 28170 4584 28226 4593
rect 28170 4519 28226 4528
rect 28276 3466 28304 5170
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 28368 4622 28396 4655
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 28368 3670 28396 4014
rect 28460 3942 28488 5714
rect 28552 3942 28580 9454
rect 28644 8294 28672 9658
rect 28736 8974 28764 10406
rect 28814 10367 28870 10376
rect 28828 9568 28856 10367
rect 28920 10146 28948 11086
rect 29092 11076 29144 11082
rect 29092 11018 29144 11024
rect 29104 10810 29132 11018
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 28920 10118 29132 10146
rect 29104 10062 29132 10118
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 29012 9722 29040 9998
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 29000 9580 29052 9586
rect 28828 9540 29000 9568
rect 29000 9522 29052 9528
rect 28906 9480 28962 9489
rect 29196 9466 29224 11630
rect 28906 9415 28962 9424
rect 29012 9438 29224 9466
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28920 8906 28948 9415
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 28724 8424 28776 8430
rect 28920 8401 28948 8842
rect 28724 8366 28776 8372
rect 28906 8392 28962 8401
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28632 7948 28684 7954
rect 28736 7936 28764 8366
rect 28906 8327 28962 8336
rect 28684 7908 28764 7936
rect 28816 7948 28868 7954
rect 28632 7890 28684 7896
rect 29012 7936 29040 9438
rect 29288 9330 29316 13806
rect 29380 12306 29408 14418
rect 29368 12300 29420 12306
rect 29368 12242 29420 12248
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 29380 10810 29408 10950
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29196 9302 29316 9330
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29104 8634 29132 8910
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29104 7954 29132 8230
rect 28816 7890 28868 7896
rect 28920 7908 29040 7936
rect 29092 7948 29144 7954
rect 28644 7342 28672 7890
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28644 6254 28672 7278
rect 28828 7206 28856 7890
rect 28920 7750 28948 7908
rect 29092 7890 29144 7896
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 28816 7200 28868 7206
rect 28816 7142 28868 7148
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 28632 6248 28684 6254
rect 28632 6190 28684 6196
rect 28644 5166 28672 6190
rect 28736 5574 28764 6666
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28828 6390 28856 6598
rect 28816 6384 28868 6390
rect 28816 6326 28868 6332
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 29012 5710 29040 6054
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28906 5400 28962 5409
rect 28906 5335 28962 5344
rect 28724 5296 28776 5302
rect 28724 5238 28776 5244
rect 28632 5160 28684 5166
rect 28632 5102 28684 5108
rect 28632 4752 28684 4758
rect 28630 4720 28632 4729
rect 28684 4720 28686 4729
rect 28630 4655 28686 4664
rect 28736 4214 28764 5238
rect 28920 5234 28948 5335
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 28814 4856 28870 4865
rect 28814 4791 28870 4800
rect 28828 4672 28856 4791
rect 28954 4684 29006 4690
rect 28828 4644 28954 4672
rect 28954 4626 29006 4632
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29012 4214 29040 4422
rect 28724 4208 28776 4214
rect 28724 4150 28776 4156
rect 28908 4208 28960 4214
rect 28908 4150 28960 4156
rect 29000 4208 29052 4214
rect 29000 4150 29052 4156
rect 28632 4072 28684 4078
rect 28632 4014 28684 4020
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28540 3936 28592 3942
rect 28644 3913 28672 4014
rect 28540 3878 28592 3884
rect 28630 3904 28686 3913
rect 28630 3839 28686 3848
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 28264 3460 28316 3466
rect 28264 3402 28316 3408
rect 28264 3120 28316 3126
rect 28092 3080 28264 3108
rect 27620 3062 27672 3068
rect 28264 3062 28316 3068
rect 27436 3052 27568 3058
rect 27488 3046 27568 3052
rect 27436 2994 27488 3000
rect 27632 800 27660 3062
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 27816 1057 27844 2382
rect 28172 1692 28224 1698
rect 28172 1634 28224 1640
rect 27896 1624 27948 1630
rect 27896 1566 27948 1572
rect 27802 1048 27858 1057
rect 27802 983 27858 992
rect 27908 800 27936 1566
rect 28184 800 28212 1634
rect 28276 1562 28304 3062
rect 28368 3058 28396 3606
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 28552 3097 28580 3402
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28538 3088 28594 3097
rect 28356 3052 28408 3058
rect 28538 3023 28594 3032
rect 28356 2994 28408 3000
rect 28644 2922 28672 3334
rect 28356 2916 28408 2922
rect 28356 2858 28408 2864
rect 28632 2916 28684 2922
rect 28632 2858 28684 2864
rect 28368 2446 28396 2858
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28448 2032 28500 2038
rect 28448 1974 28500 1980
rect 28264 1556 28316 1562
rect 28264 1498 28316 1504
rect 28460 800 28488 1974
rect 25792 734 25912 762
rect 25792 610 25820 734
rect 25780 604 25832 610
rect 25780 546 25832 552
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28644 746 28672 2858
rect 28920 2774 28948 4150
rect 28998 3632 29054 3641
rect 28998 3567 29054 3576
rect 29012 3398 29040 3567
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 28736 2746 28948 2774
rect 28736 800 28764 2746
rect 29000 2100 29052 2106
rect 29000 2042 29052 2048
rect 29012 800 29040 2042
rect 29104 1329 29132 7686
rect 29196 6390 29224 9302
rect 29472 9217 29500 9590
rect 29458 9208 29514 9217
rect 29288 9166 29458 9194
rect 29288 7274 29316 9166
rect 29458 9143 29514 9152
rect 29458 9072 29514 9081
rect 29458 9007 29514 9016
rect 29368 8900 29420 8906
rect 29368 8842 29420 8848
rect 29276 7268 29328 7274
rect 29276 7210 29328 7216
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29184 6384 29236 6390
rect 29182 6352 29184 6361
rect 29236 6352 29238 6361
rect 29182 6287 29238 6296
rect 29184 6112 29236 6118
rect 29288 6100 29316 6734
rect 29380 6322 29408 8842
rect 29472 8362 29500 9007
rect 29564 8906 29592 26930
rect 29840 25770 29868 59366
rect 29932 32570 29960 60998
rect 30300 60874 30328 63200
rect 31220 61198 31248 63294
rect 31758 63200 31814 64000
rect 32494 63200 32550 64000
rect 33230 63322 33286 64000
rect 33966 63322 34022 64000
rect 33230 63294 33548 63322
rect 33230 63200 33286 63294
rect 31772 61198 31800 63200
rect 32508 61198 32536 63200
rect 33520 61198 33548 63294
rect 33966 63294 34284 63322
rect 33966 63200 34022 63294
rect 34256 61198 34284 63294
rect 34702 63200 34758 64000
rect 35438 63322 35494 64000
rect 36174 63322 36230 64000
rect 35438 63294 35848 63322
rect 35438 63200 35494 63294
rect 31208 61192 31260 61198
rect 31760 61192 31812 61198
rect 31208 61134 31260 61140
rect 31574 61160 31630 61169
rect 31760 61134 31812 61140
rect 32496 61192 32548 61198
rect 32496 61134 32548 61140
rect 33508 61192 33560 61198
rect 33508 61134 33560 61140
rect 34244 61192 34296 61198
rect 34244 61134 34296 61140
rect 34716 61130 34744 63200
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 35072 61192 35124 61198
rect 35820 61180 35848 63294
rect 36174 63294 36400 63322
rect 36174 63200 36230 63294
rect 35900 61192 35952 61198
rect 35820 61152 35900 61180
rect 35072 61134 35124 61140
rect 35900 61134 35952 61140
rect 31574 61095 31576 61104
rect 31628 61095 31630 61104
rect 34704 61124 34756 61130
rect 31576 61066 31628 61072
rect 34704 61066 34756 61072
rect 33508 61056 33560 61062
rect 33508 60998 33560 61004
rect 34244 61056 34296 61062
rect 34244 60998 34296 61004
rect 30300 60846 30420 60874
rect 30392 60790 30420 60846
rect 30380 60784 30432 60790
rect 30380 60726 30432 60732
rect 30010 60344 30066 60353
rect 30010 60279 30012 60288
rect 30064 60279 30066 60288
rect 30012 60250 30064 60256
rect 30010 60208 30066 60217
rect 30010 60143 30066 60152
rect 30104 60172 30156 60178
rect 30024 60042 30052 60143
rect 30104 60114 30156 60120
rect 30012 60036 30064 60042
rect 30012 59978 30064 59984
rect 30116 59702 30144 60114
rect 30196 60104 30248 60110
rect 30194 60072 30196 60081
rect 30248 60072 30250 60081
rect 30194 60007 30250 60016
rect 30656 59968 30708 59974
rect 30656 59910 30708 59916
rect 33232 59968 33284 59974
rect 33232 59910 33284 59916
rect 30668 59770 30696 59910
rect 30656 59764 30708 59770
rect 30656 59706 30708 59712
rect 30104 59696 30156 59702
rect 30104 59638 30156 59644
rect 30012 59628 30064 59634
rect 30012 59570 30064 59576
rect 30024 59430 30052 59570
rect 30012 59424 30064 59430
rect 30012 59366 30064 59372
rect 30012 56364 30064 56370
rect 30012 56306 30064 56312
rect 30024 55758 30052 56306
rect 30012 55752 30064 55758
rect 30012 55694 30064 55700
rect 30024 54670 30052 55694
rect 30012 54664 30064 54670
rect 30012 54606 30064 54612
rect 30024 53582 30052 54606
rect 30012 53576 30064 53582
rect 30012 53518 30064 53524
rect 30564 45348 30616 45354
rect 30564 45290 30616 45296
rect 30576 45082 30604 45290
rect 30564 45076 30616 45082
rect 30564 45018 30616 45024
rect 30288 40112 30340 40118
rect 30288 40054 30340 40060
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 29828 25764 29880 25770
rect 29828 25706 29880 25712
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 29736 20528 29788 20534
rect 29736 20470 29788 20476
rect 29748 16658 29776 20470
rect 30116 20262 30144 20742
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29840 18766 29868 20198
rect 30116 19854 30144 20198
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 30300 19718 30328 40054
rect 30668 22778 30696 59706
rect 32404 56160 32456 56166
rect 32404 56102 32456 56108
rect 30748 44872 30800 44878
rect 30748 44814 30800 44820
rect 30656 22772 30708 22778
rect 30656 22714 30708 22720
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30392 19938 30420 19994
rect 30392 19922 30604 19938
rect 30392 19916 30616 19922
rect 30392 19910 30564 19916
rect 30564 19858 30616 19864
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30208 18970 30236 19314
rect 30012 18964 30064 18970
rect 30012 18906 30064 18912
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 30024 18698 30052 18906
rect 30300 18737 30328 19654
rect 30286 18728 30342 18737
rect 30012 18692 30064 18698
rect 30286 18663 30342 18672
rect 30012 18634 30064 18640
rect 30668 18290 30696 20402
rect 30760 18630 30788 44814
rect 31024 44804 31076 44810
rect 31024 44746 31076 44752
rect 30932 29504 30984 29510
rect 30932 29446 30984 29452
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30852 18698 30880 19654
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30748 18624 30800 18630
rect 30748 18566 30800 18572
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 29840 17338 29868 18226
rect 30472 18216 30524 18222
rect 30472 18158 30524 18164
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30300 17338 30328 17614
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 29644 16448 29696 16454
rect 29644 16390 29696 16396
rect 29656 16114 29684 16390
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29748 16028 29776 16594
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29840 16182 29868 16526
rect 29828 16176 29880 16182
rect 29828 16118 29880 16124
rect 29828 16040 29880 16046
rect 29748 16000 29828 16028
rect 29828 15982 29880 15988
rect 30010 16008 30066 16017
rect 29840 14414 29868 15982
rect 30010 15943 30066 15952
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29840 13938 29868 14350
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29734 13152 29790 13161
rect 29734 13087 29790 13096
rect 29748 12714 29776 13087
rect 29736 12708 29788 12714
rect 29736 12650 29788 12656
rect 29840 12238 29868 13874
rect 29932 13394 29960 15506
rect 30024 14346 30052 15943
rect 30104 15904 30156 15910
rect 30104 15846 30156 15852
rect 30012 14340 30064 14346
rect 30012 14282 30064 14288
rect 30012 14000 30064 14006
rect 30012 13942 30064 13948
rect 29920 13388 29972 13394
rect 29920 13330 29972 13336
rect 30024 13161 30052 13942
rect 30116 13569 30144 15846
rect 30194 15056 30250 15065
rect 30194 14991 30250 15000
rect 30208 14006 30236 14991
rect 30196 14000 30248 14006
rect 30196 13942 30248 13948
rect 30102 13560 30158 13569
rect 30102 13495 30158 13504
rect 30104 13184 30156 13190
rect 30010 13152 30066 13161
rect 30104 13126 30156 13132
rect 30010 13087 30066 13096
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 29840 11626 29868 12174
rect 30024 12170 30052 13087
rect 30116 12209 30144 13126
rect 30300 12434 30328 16934
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30392 15745 30420 16730
rect 30378 15736 30434 15745
rect 30378 15671 30434 15680
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30208 12406 30328 12434
rect 30102 12200 30158 12209
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 30012 12164 30064 12170
rect 30102 12135 30158 12144
rect 30012 12106 30064 12112
rect 29828 11620 29880 11626
rect 29828 11562 29880 11568
rect 29932 11529 29960 12106
rect 30208 12102 30236 12406
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 29918 11520 29974 11529
rect 29918 11455 29974 11464
rect 30024 11286 30052 11834
rect 30104 11620 30156 11626
rect 30104 11562 30156 11568
rect 30012 11280 30064 11286
rect 30012 11222 30064 11228
rect 30116 11150 30144 11562
rect 30104 11144 30156 11150
rect 29918 11112 29974 11121
rect 30104 11086 30156 11092
rect 29918 11047 29974 11056
rect 29736 9716 29788 9722
rect 29736 9658 29788 9664
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29656 9081 29684 9590
rect 29642 9072 29698 9081
rect 29642 9007 29698 9016
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29552 8900 29604 8906
rect 29552 8842 29604 8848
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29564 7002 29592 7142
rect 29552 6996 29604 7002
rect 29552 6938 29604 6944
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29472 6458 29500 6802
rect 29460 6452 29512 6458
rect 29460 6394 29512 6400
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29236 6072 29316 6100
rect 29184 6054 29236 6060
rect 29196 5710 29224 6054
rect 29368 5840 29420 5846
rect 29368 5782 29420 5788
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29196 5234 29224 5646
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29196 4622 29224 5170
rect 29184 4616 29236 4622
rect 29380 4593 29408 5782
rect 29564 5234 29592 6938
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29184 4558 29236 4564
rect 29366 4584 29422 4593
rect 29366 4519 29422 4528
rect 29184 4480 29236 4486
rect 29380 4434 29408 4519
rect 29184 4422 29236 4428
rect 29196 4282 29224 4422
rect 29288 4406 29408 4434
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 29184 3936 29236 3942
rect 29184 3878 29236 3884
rect 29196 3738 29224 3878
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29090 1320 29146 1329
rect 29090 1255 29146 1264
rect 29196 1154 29224 3130
rect 29288 2446 29316 4406
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29380 2650 29408 4218
rect 29472 4185 29500 5102
rect 29458 4176 29514 4185
rect 29458 4111 29514 4120
rect 29460 4072 29512 4078
rect 29458 4040 29460 4049
rect 29512 4040 29514 4049
rect 29458 3975 29514 3984
rect 29564 3602 29592 5170
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29276 2440 29328 2446
rect 29276 2382 29328 2388
rect 29380 2106 29408 2586
rect 29368 2100 29420 2106
rect 29368 2042 29420 2048
rect 29276 1896 29328 1902
rect 29276 1838 29328 1844
rect 29184 1148 29236 1154
rect 29184 1090 29236 1096
rect 29288 800 29316 1838
rect 29472 1714 29500 3538
rect 29552 3460 29604 3466
rect 29552 3402 29604 3408
rect 29564 3194 29592 3402
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29656 1902 29684 8910
rect 29748 8498 29776 9658
rect 29828 9444 29880 9450
rect 29828 9386 29880 9392
rect 29840 8974 29868 9386
rect 29932 9353 29960 11047
rect 30010 10840 30066 10849
rect 30010 10775 30066 10784
rect 29918 9344 29974 9353
rect 29918 9279 29974 9288
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29734 6896 29790 6905
rect 29734 6831 29790 6840
rect 29748 6322 29776 6831
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29932 6254 29960 9279
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 30024 6202 30052 10775
rect 30104 10532 30156 10538
rect 30104 10474 30156 10480
rect 30116 9761 30144 10474
rect 30102 9752 30158 9761
rect 30102 9687 30158 9696
rect 30102 9344 30158 9353
rect 30102 9279 30158 9288
rect 30116 8498 30144 9279
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30102 8256 30158 8265
rect 30102 8191 30158 8200
rect 30116 7886 30144 8191
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7478 30144 7686
rect 30104 7472 30156 7478
rect 30104 7414 30156 7420
rect 30208 6866 30236 12038
rect 30392 11830 30420 13194
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30300 9722 30328 10066
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30300 8022 30328 9522
rect 30288 8016 30340 8022
rect 30288 7958 30340 7964
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30300 7721 30328 7822
rect 30392 7750 30420 11766
rect 30484 9722 30512 18158
rect 30852 18086 30880 18634
rect 30840 18080 30892 18086
rect 30840 18022 30892 18028
rect 30748 16992 30800 16998
rect 30748 16934 30800 16940
rect 30760 16658 30788 16934
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 30748 16652 30800 16658
rect 30748 16594 30800 16600
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30576 14958 30604 15302
rect 30668 15026 30696 15846
rect 30748 15360 30800 15366
rect 30748 15302 30800 15308
rect 30656 15020 30708 15026
rect 30656 14962 30708 14968
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30760 14793 30788 15302
rect 30852 15162 30880 16730
rect 30944 15502 30972 29446
rect 31036 26353 31064 44746
rect 32128 36372 32180 36378
rect 32128 36314 32180 36320
rect 31760 34196 31812 34202
rect 31760 34138 31812 34144
rect 31772 32502 31800 34138
rect 31760 32496 31812 32502
rect 31760 32438 31812 32444
rect 31022 26344 31078 26353
rect 31022 26279 31078 26288
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31404 18426 31432 20742
rect 31852 20256 31904 20262
rect 31852 20198 31904 20204
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31392 18420 31444 18426
rect 31392 18362 31444 18368
rect 31588 18222 31616 19246
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 31036 16590 31064 18022
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 31128 16454 31156 18158
rect 31392 18080 31444 18086
rect 31392 18022 31444 18028
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31312 17202 31340 17614
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31208 17128 31260 17134
rect 31206 17096 31208 17105
rect 31260 17096 31262 17105
rect 31206 17031 31262 17040
rect 31116 16448 31168 16454
rect 31114 16416 31116 16425
rect 31168 16416 31170 16425
rect 31114 16351 31170 16360
rect 31300 15632 31352 15638
rect 31300 15574 31352 15580
rect 30932 15496 30984 15502
rect 30932 15438 30984 15444
rect 30944 15162 30972 15438
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 30746 14784 30802 14793
rect 30746 14719 30802 14728
rect 30760 14618 30788 14719
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30932 14544 30984 14550
rect 30932 14486 30984 14492
rect 30944 13870 30972 14486
rect 31036 14006 31064 15030
rect 31116 14952 31168 14958
rect 31116 14894 31168 14900
rect 31128 14550 31156 14894
rect 31208 14884 31260 14890
rect 31208 14826 31260 14832
rect 31116 14544 31168 14550
rect 31116 14486 31168 14492
rect 31024 14000 31076 14006
rect 31024 13942 31076 13948
rect 30932 13864 30984 13870
rect 30932 13806 30984 13812
rect 31128 13734 31156 14486
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30576 10810 30604 11698
rect 30944 11558 30972 11834
rect 30656 11552 30708 11558
rect 30656 11494 30708 11500
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30932 11552 30984 11558
rect 30932 11494 30984 11500
rect 30668 11014 30696 11494
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30472 9716 30524 9722
rect 30472 9658 30524 9664
rect 30380 7744 30432 7750
rect 30286 7712 30342 7721
rect 30380 7686 30432 7692
rect 30286 7647 30342 7656
rect 30300 7002 30328 7647
rect 30288 6996 30340 7002
rect 30288 6938 30340 6944
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30102 6216 30158 6225
rect 30024 6174 30102 6202
rect 30102 6151 30158 6160
rect 30010 5944 30066 5953
rect 30010 5879 30066 5888
rect 29736 5772 29788 5778
rect 29736 5714 29788 5720
rect 29748 4078 29776 5714
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29840 4826 29868 5170
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29736 4072 29788 4078
rect 29920 4072 29972 4078
rect 29736 4014 29788 4020
rect 29840 4032 29920 4060
rect 29736 3596 29788 3602
rect 29840 3584 29868 4032
rect 30024 4049 30052 5879
rect 30116 4622 30144 6151
rect 30300 5817 30328 6258
rect 30286 5808 30342 5817
rect 30286 5743 30342 5752
rect 30196 5296 30248 5302
rect 30196 5238 30248 5244
rect 30208 5030 30236 5238
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30300 4690 30328 4966
rect 30288 4684 30340 4690
rect 30288 4626 30340 4632
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 29920 4014 29972 4020
rect 30010 4040 30066 4049
rect 30010 3975 30066 3984
rect 29920 3936 29972 3942
rect 29920 3878 29972 3884
rect 29788 3556 29868 3584
rect 29736 3538 29788 3544
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29840 3194 29868 3402
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 29932 3058 29960 3878
rect 30024 3194 30052 3975
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 30208 2990 30236 3334
rect 30392 3074 30420 6598
rect 30484 5778 30512 6802
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 30576 5658 30604 10610
rect 30656 10532 30708 10538
rect 30656 10474 30708 10480
rect 30668 5953 30696 10474
rect 30746 9208 30802 9217
rect 30746 9143 30802 9152
rect 30760 9110 30788 9143
rect 30748 9104 30800 9110
rect 30748 9046 30800 9052
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30760 7206 30788 8910
rect 30852 8838 30880 11494
rect 31036 11150 31064 12174
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31128 10810 31156 10950
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31220 10130 31248 14826
rect 31312 14346 31340 15574
rect 31300 14340 31352 14346
rect 31300 14282 31352 14288
rect 31404 12782 31432 18022
rect 31588 17134 31616 18158
rect 31760 18148 31812 18154
rect 31760 18090 31812 18096
rect 31772 17746 31800 18090
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31576 17128 31628 17134
rect 31496 17088 31576 17116
rect 31496 15638 31524 17088
rect 31576 17070 31628 17076
rect 31484 15632 31536 15638
rect 31484 15574 31536 15580
rect 31496 15366 31524 15574
rect 31864 15434 31892 20198
rect 32140 16289 32168 36314
rect 32416 20874 32444 56102
rect 32956 42560 33008 42566
rect 32956 42502 33008 42508
rect 32772 27872 32824 27878
rect 32772 27814 32824 27820
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32404 20868 32456 20874
rect 32404 20810 32456 20816
rect 32508 20618 32536 25842
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32600 22094 32628 22918
rect 32600 22066 32720 22094
rect 32508 20590 32628 20618
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32508 17882 32536 20402
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32404 16992 32456 16998
rect 32404 16934 32456 16940
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32126 16280 32182 16289
rect 32126 16215 32182 16224
rect 32232 16182 32260 16458
rect 32220 16176 32272 16182
rect 32220 16118 32272 16124
rect 32416 16114 32444 16934
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32324 15502 32352 16050
rect 32600 15994 32628 20590
rect 32692 17202 32720 22066
rect 32680 17196 32732 17202
rect 32680 17138 32732 17144
rect 32692 16726 32720 17138
rect 32680 16720 32732 16726
rect 32680 16662 32732 16668
rect 32508 15966 32628 15994
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31852 15428 31904 15434
rect 31852 15370 31904 15376
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31484 14884 31536 14890
rect 31484 14826 31536 14832
rect 31496 12782 31524 14826
rect 31588 14822 31616 15370
rect 32218 15192 32274 15201
rect 32218 15127 32274 15136
rect 32036 15020 32088 15026
rect 32036 14962 32088 14968
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 31392 12776 31444 12782
rect 31392 12718 31444 12724
rect 31484 12776 31536 12782
rect 31536 12736 31708 12764
rect 31484 12718 31536 12724
rect 31680 12306 31708 12736
rect 31576 12300 31628 12306
rect 31576 12242 31628 12248
rect 31668 12300 31720 12306
rect 31668 12242 31720 12248
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31312 11694 31340 11834
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31298 10840 31354 10849
rect 31298 10775 31300 10784
rect 31352 10775 31354 10784
rect 31300 10746 31352 10752
rect 31404 10690 31432 11630
rect 31312 10662 31432 10690
rect 31208 10124 31260 10130
rect 31208 10066 31260 10072
rect 30932 9716 30984 9722
rect 30932 9658 30984 9664
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 30748 7200 30800 7206
rect 30748 7142 30800 7148
rect 30654 5944 30710 5953
rect 30654 5879 30710 5888
rect 30576 5630 30788 5658
rect 30656 5568 30708 5574
rect 30654 5536 30656 5545
rect 30708 5536 30710 5545
rect 30654 5471 30710 5480
rect 30564 5092 30616 5098
rect 30564 5034 30616 5040
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 30484 4185 30512 4626
rect 30470 4176 30526 4185
rect 30470 4111 30526 4120
rect 30484 3126 30512 4111
rect 30300 3058 30420 3074
rect 30472 3120 30524 3126
rect 30472 3062 30524 3068
rect 30288 3052 30420 3058
rect 30340 3046 30420 3052
rect 30288 2994 30340 3000
rect 30196 2984 30248 2990
rect 30102 2952 30158 2961
rect 30196 2926 30248 2932
rect 30102 2887 30158 2896
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 29644 1896 29696 1902
rect 29644 1838 29696 1844
rect 29472 1686 29592 1714
rect 29564 800 29592 1686
rect 29840 800 29868 2314
rect 30116 800 30144 2887
rect 30208 2774 30236 2926
rect 30208 2746 30328 2774
rect 30300 2009 30328 2746
rect 30576 2553 30604 5034
rect 30668 4826 30696 5471
rect 30656 4820 30708 4826
rect 30656 4762 30708 4768
rect 30760 3126 30788 5630
rect 30852 4554 30880 7686
rect 30840 4548 30892 4554
rect 30840 4490 30892 4496
rect 30944 3534 30972 9658
rect 31116 9648 31168 9654
rect 31116 9590 31168 9596
rect 31206 9616 31262 9625
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 31036 8430 31064 9522
rect 31128 9330 31156 9590
rect 31206 9551 31208 9560
rect 31260 9551 31262 9560
rect 31208 9522 31260 9528
rect 31312 9450 31340 10662
rect 31300 9444 31352 9450
rect 31300 9386 31352 9392
rect 31128 9302 31340 9330
rect 31312 8634 31340 9302
rect 31392 8968 31444 8974
rect 31392 8910 31444 8916
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31036 7274 31064 7822
rect 31114 7712 31170 7721
rect 31114 7647 31170 7656
rect 31128 7546 31156 7647
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31024 7268 31076 7274
rect 31024 7210 31076 7216
rect 31220 7206 31248 8230
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31114 6896 31170 6905
rect 31114 6831 31170 6840
rect 31128 6798 31156 6831
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 31036 6089 31064 6666
rect 31220 6633 31248 6734
rect 31206 6624 31262 6633
rect 31206 6559 31262 6568
rect 31116 6112 31168 6118
rect 31022 6080 31078 6089
rect 31116 6054 31168 6060
rect 31022 6015 31078 6024
rect 31036 5817 31064 6015
rect 31022 5808 31078 5817
rect 31022 5743 31078 5752
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 31036 5302 31064 5646
rect 31024 5296 31076 5302
rect 31024 5238 31076 5244
rect 31128 5098 31156 6054
rect 31116 5092 31168 5098
rect 31116 5034 31168 5040
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 31312 3058 31340 8570
rect 31404 5250 31432 8910
rect 31496 8498 31524 12038
rect 31588 11694 31616 12242
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31576 10600 31628 10606
rect 31680 10554 31708 12242
rect 31956 12102 31984 13466
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31628 10548 31800 10554
rect 31576 10542 31800 10548
rect 31588 10538 31800 10542
rect 31588 10532 31812 10538
rect 31588 10526 31760 10532
rect 31760 10474 31812 10480
rect 31850 10160 31906 10169
rect 31850 10095 31852 10104
rect 31904 10095 31906 10104
rect 31852 10066 31904 10072
rect 31574 9616 31630 9625
rect 31760 9580 31812 9586
rect 31574 9551 31576 9560
rect 31628 9551 31630 9560
rect 31576 9522 31628 9528
rect 31680 9540 31760 9568
rect 31576 9444 31628 9450
rect 31576 9386 31628 9392
rect 31588 8809 31616 9386
rect 31574 8800 31630 8809
rect 31574 8735 31630 8744
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 31680 8129 31708 9540
rect 31760 9522 31812 9528
rect 31944 9376 31996 9382
rect 31944 9318 31996 9324
rect 31758 9208 31814 9217
rect 31758 9143 31814 9152
rect 31772 9110 31800 9143
rect 31760 9104 31812 9110
rect 31760 9046 31812 9052
rect 31760 8832 31812 8838
rect 31760 8774 31812 8780
rect 31666 8120 31722 8129
rect 31666 8055 31722 8064
rect 31772 7290 31800 8774
rect 31956 8401 31984 9318
rect 31942 8392 31998 8401
rect 31942 8327 31998 8336
rect 31772 7262 31892 7290
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31760 7200 31812 7206
rect 31760 7142 31812 7148
rect 31496 6662 31524 7142
rect 31576 6724 31628 6730
rect 31576 6666 31628 6672
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 31484 6112 31536 6118
rect 31484 6054 31536 6060
rect 31496 5846 31524 6054
rect 31484 5840 31536 5846
rect 31484 5782 31536 5788
rect 31484 5568 31536 5574
rect 31484 5510 31536 5516
rect 31496 5370 31524 5510
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 31404 5222 31524 5250
rect 31392 5160 31444 5166
rect 31390 5128 31392 5137
rect 31444 5128 31446 5137
rect 31496 5098 31524 5222
rect 31390 5063 31446 5072
rect 31484 5092 31536 5098
rect 31404 3738 31432 5063
rect 31484 5034 31536 5040
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 30562 2544 30618 2553
rect 30380 2508 30432 2514
rect 30562 2479 30618 2488
rect 30380 2450 30432 2456
rect 30286 2000 30342 2009
rect 30286 1935 30342 1944
rect 30392 800 30420 2450
rect 30656 2372 30708 2378
rect 30656 2314 30708 2320
rect 30932 2372 30984 2378
rect 30932 2314 30984 2320
rect 30668 800 30696 2314
rect 30944 800 30972 2314
rect 31220 800 31248 2926
rect 31484 2372 31536 2378
rect 31484 2314 31536 2320
rect 31496 800 31524 2314
rect 31588 1970 31616 6666
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 31680 6390 31708 6598
rect 31668 6384 31720 6390
rect 31668 6326 31720 6332
rect 31668 5636 31720 5642
rect 31668 5578 31720 5584
rect 31680 5545 31708 5578
rect 31666 5536 31722 5545
rect 31666 5471 31722 5480
rect 31772 5234 31800 7142
rect 31864 6118 31892 7262
rect 31852 6112 31904 6118
rect 31852 6054 31904 6060
rect 31852 5636 31904 5642
rect 31852 5578 31904 5584
rect 31864 5545 31892 5578
rect 31850 5536 31906 5545
rect 31850 5471 31906 5480
rect 31850 5400 31906 5409
rect 31850 5335 31906 5344
rect 31864 5234 31892 5335
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 31852 5228 31904 5234
rect 31852 5170 31904 5176
rect 31956 5166 31984 8327
rect 32048 8090 32076 14962
rect 32232 12442 32260 15127
rect 32312 13456 32364 13462
rect 32312 13398 32364 13404
rect 32220 12436 32272 12442
rect 32220 12378 32272 12384
rect 32324 11150 32352 13398
rect 32402 13288 32458 13297
rect 32402 13223 32458 13232
rect 32416 11830 32444 13223
rect 32508 12918 32536 15966
rect 32784 15094 32812 27814
rect 32968 22438 32996 42502
rect 33140 36712 33192 36718
rect 33140 36654 33192 36660
rect 33152 35698 33180 36654
rect 33140 35692 33192 35698
rect 33140 35634 33192 35640
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33060 18834 33088 19790
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 33152 18086 33180 19110
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 33244 16574 33272 59910
rect 33324 56704 33376 56710
rect 33322 56672 33324 56681
rect 33376 56672 33378 56681
rect 33322 56607 33378 56616
rect 33520 42770 33548 60998
rect 34256 60734 34284 60998
rect 34164 60706 34284 60734
rect 35084 60722 35112 61134
rect 35348 61056 35400 61062
rect 35348 60998 35400 61004
rect 36084 61056 36136 61062
rect 36084 60998 36136 61004
rect 35072 60716 35124 60722
rect 34164 60110 34192 60706
rect 35072 60658 35124 60664
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 33784 60104 33836 60110
rect 33784 60046 33836 60052
rect 34152 60104 34204 60110
rect 34152 60046 34204 60052
rect 33796 59770 33824 60046
rect 33784 59764 33836 59770
rect 33784 59706 33836 59712
rect 33796 56846 33824 59706
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 34520 58948 34572 58954
rect 34520 58890 34572 58896
rect 34532 57050 34560 58890
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34520 57044 34572 57050
rect 34520 56986 34572 56992
rect 33784 56840 33836 56846
rect 33784 56782 33836 56788
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34612 52556 34664 52562
rect 34612 52498 34664 52504
rect 34244 46368 34296 46374
rect 34244 46310 34296 46316
rect 34060 43716 34112 43722
rect 34060 43658 34112 43664
rect 33968 43648 34020 43654
rect 33968 43590 34020 43596
rect 33980 43314 34008 43590
rect 34072 43314 34100 43658
rect 34256 43382 34284 46310
rect 34244 43376 34296 43382
rect 34244 43318 34296 43324
rect 33968 43308 34020 43314
rect 33968 43250 34020 43256
rect 34060 43308 34112 43314
rect 34060 43250 34112 43256
rect 34072 43194 34100 43250
rect 33980 43166 34100 43194
rect 33508 42764 33560 42770
rect 33508 42706 33560 42712
rect 33980 42702 34008 43166
rect 34520 43104 34572 43110
rect 34520 43046 34572 43052
rect 34532 42945 34560 43046
rect 34518 42936 34574 42945
rect 34518 42871 34574 42880
rect 33968 42696 34020 42702
rect 33968 42638 34020 42644
rect 33324 40112 33376 40118
rect 33324 40054 33376 40060
rect 33336 17678 33364 40054
rect 33980 36854 34008 42638
rect 34060 39092 34112 39098
rect 34060 39034 34112 39040
rect 34072 38962 34100 39034
rect 34060 38956 34112 38962
rect 34060 38898 34112 38904
rect 34428 38956 34480 38962
rect 34428 38898 34480 38904
rect 33968 36848 34020 36854
rect 33968 36790 34020 36796
rect 34440 35834 34468 38898
rect 34624 38826 34652 52498
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34796 49156 34848 49162
rect 34796 49098 34848 49104
rect 34612 38820 34664 38826
rect 34612 38762 34664 38768
rect 34428 35828 34480 35834
rect 34428 35770 34480 35776
rect 34440 34542 34468 35770
rect 33600 34536 33652 34542
rect 33600 34478 33652 34484
rect 34428 34536 34480 34542
rect 34428 34478 34480 34484
rect 33508 20596 33560 20602
rect 33508 20538 33560 20544
rect 33520 19514 33548 20538
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 33508 18080 33560 18086
rect 33508 18022 33560 18028
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 33244 16546 33364 16574
rect 33048 16448 33100 16454
rect 33048 16390 33100 16396
rect 33060 16250 33088 16390
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32772 15088 32824 15094
rect 32772 15030 32824 15036
rect 32784 13920 32812 15030
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32968 13938 32996 14894
rect 32692 13892 32812 13920
rect 32956 13932 33008 13938
rect 32692 13394 32720 13892
rect 32956 13874 33008 13880
rect 32864 13456 32916 13462
rect 32864 13398 32916 13404
rect 32680 13388 32732 13394
rect 32680 13330 32732 13336
rect 32586 13152 32642 13161
rect 32586 13087 32642 13096
rect 32600 12918 32628 13087
rect 32496 12912 32548 12918
rect 32494 12880 32496 12889
rect 32588 12912 32640 12918
rect 32548 12880 32550 12889
rect 32588 12854 32640 12860
rect 32494 12815 32550 12824
rect 32876 12714 32904 13398
rect 32968 13258 32996 13874
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 32956 13252 33008 13258
rect 32956 13194 33008 13200
rect 32968 12850 32996 13194
rect 33138 13016 33194 13025
rect 33138 12951 33194 12960
rect 33046 12880 33102 12889
rect 32956 12844 33008 12850
rect 33046 12815 33102 12824
rect 32956 12786 33008 12792
rect 32864 12708 32916 12714
rect 32864 12650 32916 12656
rect 32680 12640 32732 12646
rect 32678 12608 32680 12617
rect 32732 12608 32734 12617
rect 32678 12543 32734 12552
rect 32770 12472 32826 12481
rect 32770 12407 32826 12416
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32404 11824 32456 11830
rect 32404 11766 32456 11772
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32416 10810 32444 11562
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 32508 10674 32536 12038
rect 32680 11008 32732 11014
rect 32680 10950 32732 10956
rect 32586 10704 32642 10713
rect 32496 10668 32548 10674
rect 32586 10639 32588 10648
rect 32496 10610 32548 10616
rect 32640 10639 32642 10648
rect 32588 10610 32640 10616
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 32416 9722 32444 10066
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32128 9376 32180 9382
rect 32128 9318 32180 9324
rect 32140 8537 32168 9318
rect 32312 8560 32364 8566
rect 32126 8528 32182 8537
rect 32312 8502 32364 8508
rect 32126 8463 32182 8472
rect 32036 8084 32088 8090
rect 32036 8026 32088 8032
rect 32036 7404 32088 7410
rect 32036 7346 32088 7352
rect 31944 5160 31996 5166
rect 31944 5102 31996 5108
rect 32048 5098 32076 7346
rect 32036 5092 32088 5098
rect 32036 5034 32088 5040
rect 32140 4978 32168 8463
rect 32324 7954 32352 8502
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32312 7948 32364 7954
rect 32312 7890 32364 7896
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 32232 5574 32260 6598
rect 32324 6322 32352 7890
rect 32416 7313 32444 8366
rect 32402 7304 32458 7313
rect 32402 7239 32458 7248
rect 32508 6390 32536 10610
rect 32588 10532 32640 10538
rect 32588 10474 32640 10480
rect 32600 8566 32628 10474
rect 32692 9926 32720 10950
rect 32784 10130 32812 12407
rect 32956 12164 33008 12170
rect 32956 12106 33008 12112
rect 32862 11520 32918 11529
rect 32862 11455 32918 11464
rect 32876 10742 32904 11455
rect 32968 11014 32996 12106
rect 33060 11694 33088 12815
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 33152 10742 33180 12951
rect 33244 12442 33272 13466
rect 33232 12436 33284 12442
rect 33232 12378 33284 12384
rect 33336 12050 33364 16546
rect 33428 15910 33456 17478
rect 33520 17270 33548 18022
rect 33508 17264 33560 17270
rect 33508 17206 33560 17212
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33428 15638 33456 15846
rect 33416 15632 33468 15638
rect 33416 15574 33468 15580
rect 33612 13326 33640 34478
rect 34808 26234 34836 49098
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35164 43716 35216 43722
rect 35360 43704 35388 60998
rect 35624 60512 35676 60518
rect 35624 60454 35676 60460
rect 35716 60512 35768 60518
rect 35716 60454 35768 60460
rect 35530 60072 35586 60081
rect 35636 60042 35664 60454
rect 35530 60007 35586 60016
rect 35624 60036 35676 60042
rect 35544 59634 35572 60007
rect 35624 59978 35676 59984
rect 35532 59628 35584 59634
rect 35532 59570 35584 59576
rect 35544 56370 35572 59570
rect 35728 56930 35756 60454
rect 35728 56902 35940 56930
rect 35912 56846 35940 56902
rect 35624 56840 35676 56846
rect 35624 56782 35676 56788
rect 35900 56840 35952 56846
rect 35900 56782 35952 56788
rect 35992 56840 36044 56846
rect 35992 56782 36044 56788
rect 35636 56506 35664 56782
rect 35624 56500 35676 56506
rect 35624 56442 35676 56448
rect 35532 56364 35584 56370
rect 35532 56306 35584 56312
rect 36004 52562 36032 56782
rect 35992 52556 36044 52562
rect 35992 52498 36044 52504
rect 35440 43920 35492 43926
rect 35440 43862 35492 43868
rect 35216 43676 35388 43704
rect 35164 43658 35216 43664
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35348 33992 35400 33998
rect 35348 33934 35400 33940
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34624 26206 34836 26234
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34440 22094 34468 22374
rect 34164 22066 34468 22094
rect 33784 20868 33836 20874
rect 33784 20810 33836 20816
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33704 17270 33732 17478
rect 33692 17264 33744 17270
rect 33692 17206 33744 17212
rect 33690 17096 33746 17105
rect 33690 17031 33746 17040
rect 33704 16250 33732 17031
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33704 14958 33732 15982
rect 33692 14952 33744 14958
rect 33692 14894 33744 14900
rect 33796 14657 33824 20810
rect 33968 18692 34020 18698
rect 33968 18634 34020 18640
rect 33876 18080 33928 18086
rect 33876 18022 33928 18028
rect 33782 14648 33838 14657
rect 33782 14583 33838 14592
rect 33888 14550 33916 18022
rect 33980 17134 34008 18634
rect 33968 17128 34020 17134
rect 33968 17070 34020 17076
rect 33968 15904 34020 15910
rect 33968 15846 34020 15852
rect 33980 15094 34008 15846
rect 34058 15736 34114 15745
rect 34058 15671 34114 15680
rect 34072 15638 34100 15671
rect 34060 15632 34112 15638
rect 34060 15574 34112 15580
rect 34072 15502 34100 15574
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33968 15088 34020 15094
rect 33968 15030 34020 15036
rect 34058 14920 34114 14929
rect 34058 14855 34114 14864
rect 33966 14648 34022 14657
rect 33966 14583 34022 14592
rect 33876 14544 33928 14550
rect 33876 14486 33928 14492
rect 33876 14408 33928 14414
rect 33876 14350 33928 14356
rect 33888 14226 33916 14350
rect 33980 14346 34008 14583
rect 33968 14340 34020 14346
rect 33968 14282 34020 14288
rect 34072 14226 34100 14855
rect 33888 14198 34100 14226
rect 33876 13864 33928 13870
rect 33876 13806 33928 13812
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 33416 13252 33468 13258
rect 33416 13194 33468 13200
rect 33428 12322 33456 13194
rect 33612 12617 33640 13262
rect 33598 12608 33654 12617
rect 33598 12543 33654 12552
rect 33428 12294 33732 12322
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33506 12200 33562 12209
rect 33244 12022 33364 12050
rect 32864 10736 32916 10742
rect 32864 10678 32916 10684
rect 33140 10736 33192 10742
rect 33140 10678 33192 10684
rect 32862 10432 32918 10441
rect 32862 10367 32918 10376
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32678 9752 32734 9761
rect 32678 9687 32680 9696
rect 32732 9687 32734 9696
rect 32680 9658 32732 9664
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32784 9178 32812 9522
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 32680 9104 32732 9110
rect 32680 9046 32732 9052
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32600 7426 32628 8502
rect 32692 7546 32720 9046
rect 32772 8016 32824 8022
rect 32772 7958 32824 7964
rect 32784 7750 32812 7958
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 32600 7398 32720 7426
rect 32588 7336 32640 7342
rect 32588 7278 32640 7284
rect 32600 6497 32628 7278
rect 32692 7274 32720 7398
rect 32680 7268 32732 7274
rect 32680 7210 32732 7216
rect 32678 6896 32734 6905
rect 32876 6882 32904 10367
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 32956 9716 33008 9722
rect 32956 9658 33008 9664
rect 32968 9625 32996 9658
rect 32954 9616 33010 9625
rect 32954 9551 33010 9560
rect 32956 9444 33008 9450
rect 32956 9386 33008 9392
rect 32968 9178 32996 9386
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32968 8945 32996 8978
rect 32954 8936 33010 8945
rect 32954 8871 33010 8880
rect 32956 8560 33008 8566
rect 32956 8502 33008 8508
rect 32968 8090 32996 8502
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32784 6866 32904 6882
rect 32678 6831 32734 6840
rect 32772 6860 32904 6866
rect 32692 6798 32720 6831
rect 32824 6854 32904 6860
rect 32772 6802 32824 6808
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32586 6488 32642 6497
rect 32586 6423 32642 6432
rect 32496 6384 32548 6390
rect 32496 6326 32548 6332
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 31864 4950 32168 4978
rect 31758 4176 31814 4185
rect 31758 4111 31814 4120
rect 31772 4010 31800 4111
rect 31760 4004 31812 4010
rect 31760 3946 31812 3952
rect 31760 2984 31812 2990
rect 31760 2926 31812 2932
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 31680 2650 31708 2790
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 31576 1964 31628 1970
rect 31576 1906 31628 1912
rect 31772 800 31800 2926
rect 31864 2774 31892 4950
rect 32324 4622 32352 6258
rect 32402 5944 32458 5953
rect 32402 5879 32458 5888
rect 32416 5681 32444 5879
rect 32402 5672 32458 5681
rect 32402 5607 32458 5616
rect 32416 5574 32444 5607
rect 32600 5574 32628 6423
rect 32404 5568 32456 5574
rect 32404 5510 32456 5516
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32402 5264 32458 5273
rect 32402 5199 32458 5208
rect 32416 5030 32444 5199
rect 32404 5024 32456 5030
rect 32404 4966 32456 4972
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32324 4434 32352 4558
rect 32324 4406 32444 4434
rect 32312 4276 32364 4282
rect 32312 4218 32364 4224
rect 32324 3466 32352 4218
rect 32416 3466 32444 4406
rect 32600 4282 32628 5510
rect 32680 5024 32732 5030
rect 32784 5001 32812 6802
rect 32680 4966 32732 4972
rect 32770 4992 32826 5001
rect 32692 4729 32720 4966
rect 32770 4927 32826 4936
rect 32678 4720 32734 4729
rect 32968 4672 32996 8026
rect 33060 7818 33088 10066
rect 33048 7812 33100 7818
rect 33048 7754 33100 7760
rect 33060 6730 33088 7754
rect 33152 7478 33180 10134
rect 33244 8634 33272 12022
rect 33428 11898 33456 12174
rect 33506 12135 33562 12144
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33336 11642 33364 11834
rect 33336 11626 33456 11642
rect 33336 11620 33468 11626
rect 33336 11614 33416 11620
rect 33416 11562 33468 11568
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 33336 11286 33364 11494
rect 33520 11286 33548 12135
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33324 11280 33376 11286
rect 33324 11222 33376 11228
rect 33508 11280 33560 11286
rect 33508 11222 33560 11228
rect 33324 11144 33376 11150
rect 33322 11112 33324 11121
rect 33376 11112 33378 11121
rect 33322 11047 33378 11056
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33336 9081 33364 10950
rect 33506 9752 33562 9761
rect 33506 9687 33562 9696
rect 33416 9580 33468 9586
rect 33416 9522 33468 9528
rect 33428 9353 33456 9522
rect 33414 9344 33470 9353
rect 33414 9279 33470 9288
rect 33416 9104 33468 9110
rect 33322 9072 33378 9081
rect 33416 9046 33468 9052
rect 33520 9058 33548 9687
rect 33612 9178 33640 11494
rect 33704 10985 33732 12294
rect 33784 12300 33836 12306
rect 33784 12242 33836 12248
rect 33796 11218 33824 12242
rect 33888 12238 33916 13806
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33876 11280 33928 11286
rect 33876 11222 33928 11228
rect 33784 11212 33836 11218
rect 33784 11154 33836 11160
rect 33690 10976 33746 10985
rect 33690 10911 33746 10920
rect 33796 10792 33824 11154
rect 33704 10764 33824 10792
rect 33704 9466 33732 10764
rect 33784 10668 33836 10674
rect 33784 10610 33836 10616
rect 33796 9994 33824 10610
rect 33784 9988 33836 9994
rect 33784 9930 33836 9936
rect 33796 9654 33824 9930
rect 33784 9648 33836 9654
rect 33784 9590 33836 9596
rect 33888 9586 33916 11222
rect 33980 10810 34008 14198
rect 34060 12436 34112 12442
rect 34060 12378 34112 12384
rect 34072 12306 34100 12378
rect 34060 12300 34112 12306
rect 34060 12242 34112 12248
rect 34060 11620 34112 11626
rect 34060 11562 34112 11568
rect 34072 11393 34100 11562
rect 34058 11384 34114 11393
rect 34058 11319 34114 11328
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 33968 10668 34020 10674
rect 33968 10610 34020 10616
rect 33980 10305 34008 10610
rect 34060 10532 34112 10538
rect 34060 10474 34112 10480
rect 34072 10441 34100 10474
rect 34058 10432 34114 10441
rect 34058 10367 34114 10376
rect 33966 10296 34022 10305
rect 33966 10231 34022 10240
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33704 9438 33824 9466
rect 33692 9376 33744 9382
rect 33692 9318 33744 9324
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33322 9007 33378 9016
rect 33232 8628 33284 8634
rect 33232 8570 33284 8576
rect 33244 8294 33272 8570
rect 33428 8566 33456 9046
rect 33520 9030 33640 9058
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33416 8560 33468 8566
rect 33416 8502 33468 8508
rect 33324 8424 33376 8430
rect 33324 8366 33376 8372
rect 33232 8288 33284 8294
rect 33232 8230 33284 8236
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33140 7268 33192 7274
rect 33140 7210 33192 7216
rect 33152 6934 33180 7210
rect 33336 7002 33364 8366
rect 33324 6996 33376 7002
rect 33324 6938 33376 6944
rect 33140 6928 33192 6934
rect 33140 6870 33192 6876
rect 33230 6896 33286 6905
rect 33230 6831 33286 6840
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33048 6724 33100 6730
rect 33048 6666 33100 6672
rect 33152 5930 33180 6734
rect 33244 6662 33272 6831
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33336 6089 33364 6938
rect 33322 6080 33378 6089
rect 33322 6015 33378 6024
rect 33152 5902 33456 5930
rect 33232 5840 33284 5846
rect 33232 5782 33284 5788
rect 33324 5840 33376 5846
rect 33324 5782 33376 5788
rect 33244 5681 33272 5782
rect 33230 5672 33286 5681
rect 33230 5607 33286 5616
rect 32678 4655 32734 4664
rect 32784 4644 32996 4672
rect 32588 4276 32640 4282
rect 32588 4218 32640 4224
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32310 3224 32366 3233
rect 32036 3188 32088 3194
rect 32310 3159 32366 3168
rect 32036 3130 32088 3136
rect 32048 2854 32076 3130
rect 32324 3058 32352 3159
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32312 3052 32364 3058
rect 32312 2994 32364 3000
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 32508 2774 32536 3062
rect 31864 2746 31984 2774
rect 31956 2446 31984 2746
rect 32324 2746 32536 2774
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 32036 2304 32088 2310
rect 32036 2246 32088 2252
rect 32048 800 32076 2246
rect 32324 800 32352 2746
rect 32784 2446 32812 4644
rect 32954 4584 33010 4593
rect 32954 4519 32956 4528
rect 33008 4519 33010 4528
rect 33140 4548 33192 4554
rect 32956 4490 33008 4496
rect 33140 4490 33192 4496
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32588 1420 32640 1426
rect 32588 1362 32640 1368
rect 32600 800 32628 1362
rect 32876 800 32904 3402
rect 33152 2836 33180 4490
rect 33232 4140 33284 4146
rect 33232 4082 33284 4088
rect 33244 3670 33272 4082
rect 33232 3664 33284 3670
rect 33230 3632 33232 3641
rect 33284 3632 33286 3641
rect 33230 3567 33286 3576
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33060 2808 33180 2836
rect 33060 2582 33088 2808
rect 33244 2774 33272 3130
rect 33152 2746 33272 2774
rect 33048 2576 33100 2582
rect 33048 2518 33100 2524
rect 33152 800 33180 2746
rect 33336 921 33364 5782
rect 33428 5710 33456 5902
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 33428 2854 33456 5510
rect 33520 5098 33548 8910
rect 33612 7274 33640 9030
rect 33704 8498 33732 9318
rect 33796 8974 33824 9438
rect 33888 9178 33916 9522
rect 33980 9518 34008 9998
rect 34058 9888 34114 9897
rect 34058 9823 34114 9832
rect 34072 9625 34100 9823
rect 34058 9616 34114 9625
rect 34058 9551 34060 9560
rect 34112 9551 34114 9560
rect 34060 9522 34112 9528
rect 33968 9512 34020 9518
rect 34164 9466 34192 22066
rect 34426 19272 34482 19281
rect 34426 19207 34482 19216
rect 34440 18970 34468 19207
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34244 18216 34296 18222
rect 34244 18158 34296 18164
rect 34256 16046 34284 18158
rect 34428 17604 34480 17610
rect 34428 17546 34480 17552
rect 34440 16182 34468 17546
rect 34428 16176 34480 16182
rect 34428 16118 34480 16124
rect 34244 16040 34296 16046
rect 34244 15982 34296 15988
rect 34440 15570 34468 16118
rect 34532 16114 34560 18566
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 34428 15564 34480 15570
rect 34428 15506 34480 15512
rect 34336 15088 34388 15094
rect 34336 15030 34388 15036
rect 34244 14544 34296 14550
rect 34244 14486 34296 14492
rect 34256 14113 34284 14486
rect 34348 14482 34376 15030
rect 34336 14476 34388 14482
rect 34336 14418 34388 14424
rect 34242 14104 34298 14113
rect 34242 14039 34298 14048
rect 34518 14104 34574 14113
rect 34518 14039 34574 14048
rect 34336 14000 34388 14006
rect 34336 13942 34388 13948
rect 34348 13818 34376 13942
rect 34348 13790 34468 13818
rect 34244 13728 34296 13734
rect 34244 13670 34296 13676
rect 34336 13728 34388 13734
rect 34336 13670 34388 13676
rect 34256 13190 34284 13670
rect 34348 13462 34376 13670
rect 34336 13456 34388 13462
rect 34336 13398 34388 13404
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34256 11121 34284 12174
rect 34334 11928 34390 11937
rect 34334 11863 34390 11872
rect 34348 11762 34376 11863
rect 34336 11756 34388 11762
rect 34336 11698 34388 11704
rect 34242 11112 34298 11121
rect 34242 11047 34298 11056
rect 34348 10962 34376 11698
rect 34440 11150 34468 13790
rect 34532 12481 34560 14039
rect 34518 12472 34574 12481
rect 34518 12407 34574 12416
rect 34520 12300 34572 12306
rect 34520 12242 34572 12248
rect 34532 11898 34560 12242
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34624 11393 34652 26206
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35070 19544 35126 19553
rect 35070 19479 35072 19488
rect 35124 19479 35126 19488
rect 35072 19450 35124 19456
rect 34796 19440 34848 19446
rect 34796 19382 34848 19388
rect 34808 18766 34836 19382
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34886 18864 34942 18873
rect 34886 18799 34942 18808
rect 34900 18766 34928 18799
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34888 18760 34940 18766
rect 34888 18702 34940 18708
rect 34704 18692 34756 18698
rect 34704 18634 34756 18640
rect 34716 16454 34744 18634
rect 34808 18426 34836 18702
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34886 17776 34942 17785
rect 34886 17711 34942 17720
rect 34900 17678 34928 17711
rect 34888 17672 34940 17678
rect 34888 17614 34940 17620
rect 34796 17332 34848 17338
rect 34796 17274 34848 17280
rect 34704 16448 34756 16454
rect 34704 16390 34756 16396
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34716 14618 34744 15438
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 34716 13977 34744 14418
rect 34808 14414 34836 17274
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34980 16720 35032 16726
rect 34980 16662 35032 16668
rect 34992 16454 35020 16662
rect 35360 16590 35388 33934
rect 35452 33930 35480 43862
rect 35532 39296 35584 39302
rect 35532 39238 35584 39244
rect 35440 33924 35492 33930
rect 35440 33866 35492 33872
rect 35544 19718 35572 39238
rect 35992 35556 36044 35562
rect 35992 35498 36044 35504
rect 36004 35086 36032 35498
rect 36096 35086 36124 60998
rect 36372 60790 36400 63294
rect 36910 63200 36966 64000
rect 37646 63200 37702 64000
rect 38382 63322 38438 64000
rect 39118 63322 39174 64000
rect 39854 63322 39910 64000
rect 40590 63322 40646 64000
rect 38382 63294 38608 63322
rect 38382 63200 38438 63294
rect 36924 61198 36952 63200
rect 37660 61198 37688 63200
rect 36912 61192 36964 61198
rect 36912 61134 36964 61140
rect 37648 61192 37700 61198
rect 38580 61180 38608 63294
rect 39118 63294 39528 63322
rect 39118 63200 39174 63294
rect 39500 61198 39528 63294
rect 39854 63294 39988 63322
rect 39854 63200 39910 63294
rect 39580 61260 39632 61266
rect 39580 61202 39632 61208
rect 38660 61192 38712 61198
rect 38580 61152 38660 61180
rect 37648 61134 37700 61140
rect 38660 61134 38712 61140
rect 39488 61192 39540 61198
rect 39488 61134 39540 61140
rect 37280 61056 37332 61062
rect 37280 60998 37332 61004
rect 39120 61056 39172 61062
rect 39120 60998 39172 61004
rect 36360 60784 36412 60790
rect 36360 60726 36412 60732
rect 36636 60648 36688 60654
rect 36636 60590 36688 60596
rect 36648 60110 36676 60590
rect 37188 60172 37240 60178
rect 37188 60114 37240 60120
rect 36636 60104 36688 60110
rect 36636 60046 36688 60052
rect 37200 59022 37228 60114
rect 37292 59022 37320 60998
rect 37188 59016 37240 59022
rect 37188 58958 37240 58964
rect 37280 59016 37332 59022
rect 37280 58958 37332 58964
rect 37556 59016 37608 59022
rect 37556 58958 37608 58964
rect 37200 56506 37228 58958
rect 36452 56500 36504 56506
rect 36452 56442 36504 56448
rect 37188 56500 37240 56506
rect 37188 56442 37240 56448
rect 36464 56370 36492 56442
rect 36452 56364 36504 56370
rect 36452 56306 36504 56312
rect 36452 53576 36504 53582
rect 36452 53518 36504 53524
rect 36268 48000 36320 48006
rect 36268 47942 36320 47948
rect 36176 43716 36228 43722
rect 36176 43658 36228 43664
rect 36188 42838 36216 43658
rect 36176 42832 36228 42838
rect 36176 42774 36228 42780
rect 36188 35630 36216 42774
rect 36176 35624 36228 35630
rect 36176 35566 36228 35572
rect 35992 35080 36044 35086
rect 35992 35022 36044 35028
rect 36084 35080 36136 35086
rect 36084 35022 36136 35028
rect 35900 33924 35952 33930
rect 35900 33866 35952 33872
rect 35532 19712 35584 19718
rect 35532 19654 35584 19660
rect 35544 19310 35572 19654
rect 35806 19544 35862 19553
rect 35806 19479 35862 19488
rect 35820 19446 35848 19479
rect 35808 19440 35860 19446
rect 35808 19382 35860 19388
rect 35532 19304 35584 19310
rect 35532 19246 35584 19252
rect 35716 19304 35768 19310
rect 35716 19246 35768 19252
rect 35728 16697 35756 19246
rect 35808 18964 35860 18970
rect 35808 18906 35860 18912
rect 35820 18766 35848 18906
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 35714 16688 35770 16697
rect 35714 16623 35716 16632
rect 35768 16623 35770 16632
rect 35716 16594 35768 16600
rect 35164 16584 35216 16590
rect 35164 16526 35216 16532
rect 35348 16584 35400 16590
rect 35728 16563 35756 16594
rect 35348 16526 35400 16532
rect 34980 16448 35032 16454
rect 34980 16390 35032 16396
rect 35176 16182 35204 16526
rect 35164 16176 35216 16182
rect 35164 16118 35216 16124
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15722 35388 16526
rect 35624 16448 35676 16454
rect 35624 16390 35676 16396
rect 35636 16250 35664 16390
rect 35624 16244 35676 16250
rect 35624 16186 35676 16192
rect 35624 16040 35676 16046
rect 35624 15982 35676 15988
rect 35268 15694 35388 15722
rect 35268 15586 35296 15694
rect 34992 15558 35296 15586
rect 35440 15564 35492 15570
rect 34888 15360 34940 15366
rect 34992 15348 35020 15558
rect 35440 15506 35492 15512
rect 35072 15496 35124 15502
rect 35072 15438 35124 15444
rect 34940 15320 35020 15348
rect 34888 15302 34940 15308
rect 35084 15201 35112 15438
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35070 15192 35126 15201
rect 35070 15127 35126 15136
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34796 14408 34848 14414
rect 34796 14350 34848 14356
rect 34702 13968 34758 13977
rect 34702 13903 34758 13912
rect 34886 13968 34942 13977
rect 34886 13903 34888 13912
rect 34940 13903 34942 13912
rect 35247 13932 35299 13938
rect 34888 13874 34940 13880
rect 35360 13920 35388 15302
rect 35299 13892 35388 13920
rect 35247 13874 35299 13880
rect 34796 13864 34848 13870
rect 35452 13852 35480 15506
rect 35532 14952 35584 14958
rect 35530 14920 35532 14929
rect 35584 14920 35586 14929
rect 35636 14890 35664 15982
rect 35806 15600 35862 15609
rect 35806 15535 35862 15544
rect 35530 14855 35586 14864
rect 35624 14884 35676 14890
rect 35624 14826 35676 14832
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35624 14272 35676 14278
rect 35624 14214 35676 14220
rect 34796 13806 34848 13812
rect 35360 13824 35480 13852
rect 34808 13462 34836 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13456 34848 13462
rect 34796 13398 34848 13404
rect 34808 12850 34836 13398
rect 35164 13388 35216 13394
rect 35360 13376 35388 13824
rect 35438 13696 35494 13705
rect 35438 13631 35494 13640
rect 35452 13530 35480 13631
rect 35440 13524 35492 13530
rect 35440 13466 35492 13472
rect 35216 13348 35388 13376
rect 35164 13330 35216 13336
rect 34980 13252 35032 13258
rect 34980 13194 35032 13200
rect 34992 13161 35020 13194
rect 34978 13152 35034 13161
rect 34978 13087 35034 13096
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34702 11520 34758 11529
rect 34702 11455 34758 11464
rect 34610 11384 34666 11393
rect 34610 11319 34666 11328
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34256 10934 34376 10962
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 34256 10010 34284 10934
rect 34336 10804 34388 10810
rect 34336 10746 34388 10752
rect 34348 10452 34376 10746
rect 34532 10742 34560 10950
rect 34716 10810 34744 11455
rect 34808 11218 34836 12786
rect 35176 12782 35204 13330
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35544 12889 35572 13194
rect 35530 12880 35586 12889
rect 35530 12815 35586 12824
rect 35164 12776 35216 12782
rect 35636 12730 35664 14214
rect 35164 12718 35216 12724
rect 35360 12702 35664 12730
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35164 12368 35216 12374
rect 35164 12310 35216 12316
rect 34886 12200 34942 12209
rect 34886 12135 34942 12144
rect 34900 12102 34928 12135
rect 34888 12096 34940 12102
rect 34888 12038 34940 12044
rect 35072 12096 35124 12102
rect 35072 12038 35124 12044
rect 34900 11694 34928 12038
rect 35084 11898 35112 12038
rect 35176 11937 35204 12310
rect 35256 12096 35308 12102
rect 35360 12084 35388 12702
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35452 12374 35480 12582
rect 35440 12368 35492 12374
rect 35440 12310 35492 12316
rect 35532 12368 35584 12374
rect 35532 12310 35584 12316
rect 35622 12336 35678 12345
rect 35440 12232 35492 12238
rect 35544 12220 35572 12310
rect 35622 12271 35624 12280
rect 35676 12271 35678 12280
rect 35624 12242 35676 12248
rect 35728 12238 35756 14418
rect 35820 13530 35848 15535
rect 35912 14226 35940 33866
rect 36280 22094 36308 47942
rect 36464 45490 36492 53518
rect 36452 45484 36504 45490
rect 36452 45426 36504 45432
rect 37096 45484 37148 45490
rect 37096 45426 37148 45432
rect 36464 43654 36492 45426
rect 37108 44810 37136 45426
rect 37568 45354 37596 58958
rect 39132 46442 39160 60998
rect 39304 58472 39356 58478
rect 39304 58414 39356 58420
rect 39316 50386 39344 58414
rect 39396 55344 39448 55350
rect 39396 55286 39448 55292
rect 39304 50380 39356 50386
rect 39304 50322 39356 50328
rect 39408 47598 39436 55286
rect 39396 47592 39448 47598
rect 39396 47534 39448 47540
rect 39120 46436 39172 46442
rect 39120 46378 39172 46384
rect 37556 45348 37608 45354
rect 37556 45290 37608 45296
rect 37648 44872 37700 44878
rect 37648 44814 37700 44820
rect 37096 44804 37148 44810
rect 37096 44746 37148 44752
rect 36452 43648 36504 43654
rect 36452 43590 36504 43596
rect 36912 42696 36964 42702
rect 36910 42664 36912 42673
rect 36964 42664 36966 42673
rect 37108 42634 37136 44746
rect 37372 44736 37424 44742
rect 37372 44678 37424 44684
rect 37188 43444 37240 43450
rect 37188 43386 37240 43392
rect 37200 42702 37228 43386
rect 37384 43314 37412 44678
rect 37372 43308 37424 43314
rect 37372 43250 37424 43256
rect 37384 42702 37412 43250
rect 37188 42696 37240 42702
rect 37188 42638 37240 42644
rect 37372 42696 37424 42702
rect 37372 42638 37424 42644
rect 36910 42599 36966 42608
rect 37096 42628 37148 42634
rect 37096 42570 37148 42576
rect 37108 42362 37136 42570
rect 37096 42356 37148 42362
rect 37096 42298 37148 42304
rect 36820 40928 36872 40934
rect 36820 40870 36872 40876
rect 36832 35086 36860 40870
rect 37280 36032 37332 36038
rect 37280 35974 37332 35980
rect 37292 35766 37320 35974
rect 37280 35760 37332 35766
rect 37280 35702 37332 35708
rect 37004 35216 37056 35222
rect 37004 35158 37056 35164
rect 36820 35080 36872 35086
rect 36820 35022 36872 35028
rect 36280 22066 36768 22094
rect 36268 20324 36320 20330
rect 36268 20266 36320 20272
rect 36280 19854 36308 20266
rect 36268 19848 36320 19854
rect 36268 19790 36320 19796
rect 36280 19310 36308 19790
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36268 19304 36320 19310
rect 36268 19246 36320 19252
rect 36280 18873 36308 19246
rect 36266 18864 36322 18873
rect 36266 18799 36322 18808
rect 35992 17672 36044 17678
rect 35992 17614 36044 17620
rect 36004 16640 36032 17614
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36096 16794 36124 17138
rect 36360 17128 36412 17134
rect 36360 17070 36412 17076
rect 36084 16788 36136 16794
rect 36084 16730 36136 16736
rect 36176 16652 36228 16658
rect 36004 16612 36176 16640
rect 36176 16594 36228 16600
rect 36176 16244 36228 16250
rect 36176 16186 36228 16192
rect 36188 15978 36216 16186
rect 36176 15972 36228 15978
rect 36176 15914 36228 15920
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 36096 15094 36124 15302
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 36188 14958 36216 15098
rect 36176 14952 36228 14958
rect 36176 14894 36228 14900
rect 36176 14612 36228 14618
rect 36176 14554 36228 14560
rect 36188 14346 36216 14554
rect 36372 14414 36400 17070
rect 36464 16250 36492 19654
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36648 18358 36676 19110
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 36544 17128 36596 17134
rect 36544 17070 36596 17076
rect 36452 16244 36504 16250
rect 36452 16186 36504 16192
rect 36452 14952 36504 14958
rect 36452 14894 36504 14900
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 36176 14340 36228 14346
rect 36176 14282 36228 14288
rect 36084 14272 36136 14278
rect 35912 14198 36032 14226
rect 36084 14214 36136 14220
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 36004 13308 36032 14198
rect 36096 13870 36124 14214
rect 36280 14074 36308 14214
rect 36268 14068 36320 14074
rect 36268 14010 36320 14016
rect 36084 13864 36136 13870
rect 36084 13806 36136 13812
rect 36268 13456 36320 13462
rect 36268 13398 36320 13404
rect 35912 13280 36032 13308
rect 35808 13184 35860 13190
rect 35806 13152 35808 13161
rect 35860 13152 35862 13161
rect 35806 13087 35862 13096
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35820 12646 35848 12786
rect 35808 12640 35860 12646
rect 35808 12582 35860 12588
rect 35492 12192 35572 12220
rect 35716 12232 35768 12238
rect 35440 12174 35492 12180
rect 35716 12174 35768 12180
rect 35808 12232 35860 12238
rect 35808 12174 35860 12180
rect 35308 12056 35388 12084
rect 35256 12038 35308 12044
rect 35162 11928 35218 11937
rect 35072 11892 35124 11898
rect 35162 11863 35218 11872
rect 35072 11834 35124 11840
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34888 11688 34940 11694
rect 34888 11630 34940 11636
rect 35360 11558 35388 11698
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 35452 10962 35480 11494
rect 35530 11112 35586 11121
rect 35530 11047 35586 11056
rect 34808 10934 35480 10962
rect 34704 10804 34756 10810
rect 34704 10746 34756 10752
rect 34520 10736 34572 10742
rect 34520 10678 34572 10684
rect 34520 10600 34572 10606
rect 34808 10588 34836 10934
rect 34572 10560 34836 10588
rect 34520 10542 34572 10548
rect 34348 10424 34652 10452
rect 34334 10296 34390 10305
rect 34334 10231 34390 10240
rect 34348 10198 34376 10231
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34520 10056 34572 10062
rect 34256 9982 34468 10010
rect 34520 9998 34572 10004
rect 34244 9648 34296 9654
rect 34242 9616 34244 9625
rect 34296 9616 34298 9625
rect 34242 9551 34298 9560
rect 33968 9454 34020 9460
rect 34072 9438 34192 9466
rect 34336 9512 34388 9518
rect 34336 9454 34388 9460
rect 33966 9344 34022 9353
rect 33966 9279 34022 9288
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 33874 8256 33930 8265
rect 33874 8191 33930 8200
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33600 6928 33652 6934
rect 33600 6870 33652 6876
rect 33612 6186 33640 6870
rect 33704 6866 33732 8026
rect 33888 7886 33916 8191
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33980 7585 34008 9279
rect 34072 9092 34100 9438
rect 34072 9064 34192 9092
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 33966 7576 34022 7585
rect 33784 7540 33836 7546
rect 33966 7511 34022 7520
rect 33784 7482 33836 7488
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33796 6798 33824 7482
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 33692 6724 33744 6730
rect 33692 6666 33744 6672
rect 33600 6180 33652 6186
rect 33600 6122 33652 6128
rect 33612 5953 33640 6122
rect 33598 5944 33654 5953
rect 33598 5879 33654 5888
rect 33598 5808 33654 5817
rect 33598 5743 33654 5752
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 33612 4622 33640 5743
rect 33600 4616 33652 4622
rect 33600 4558 33652 4564
rect 33704 4468 33732 6666
rect 33980 5817 34008 6734
rect 34072 6186 34100 8774
rect 34164 7818 34192 9064
rect 34242 8664 34298 8673
rect 34242 8599 34298 8608
rect 34256 8022 34284 8599
rect 34348 8090 34376 9454
rect 34336 8084 34388 8090
rect 34336 8026 34388 8032
rect 34244 8016 34296 8022
rect 34244 7958 34296 7964
rect 34440 7954 34468 9982
rect 34532 9058 34560 9998
rect 34624 9586 34652 10424
rect 34702 10432 34758 10441
rect 34702 10367 34758 10376
rect 34612 9580 34664 9586
rect 34612 9522 34664 9528
rect 34624 9353 34652 9522
rect 34610 9344 34666 9353
rect 34610 9279 34666 9288
rect 34716 9160 34744 10367
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34794 10296 34850 10305
rect 34934 10299 35242 10308
rect 34794 10231 34850 10240
rect 34808 10130 34836 10231
rect 34796 10124 34848 10130
rect 34796 10066 34848 10072
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 35072 10056 35124 10062
rect 35072 9998 35124 10004
rect 35256 10056 35308 10062
rect 35256 9998 35308 10004
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 9722 34836 9862
rect 34900 9722 34928 9998
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 35084 9654 35112 9998
rect 35268 9897 35296 9998
rect 35254 9888 35310 9897
rect 35254 9823 35310 9832
rect 35072 9648 35124 9654
rect 34978 9616 35034 9625
rect 34888 9580 34940 9586
rect 34808 9540 34888 9568
rect 34808 9353 34836 9540
rect 35072 9590 35124 9596
rect 34978 9551 35034 9560
rect 34888 9522 34940 9528
rect 34992 9382 35020 9551
rect 34980 9376 35032 9382
rect 34794 9344 34850 9353
rect 34980 9318 35032 9324
rect 34794 9279 34850 9288
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34716 9132 35112 9160
rect 34532 9030 34928 9058
rect 34518 8664 34574 8673
rect 34518 8599 34574 8608
rect 34532 8106 34560 8599
rect 34624 8265 34652 9030
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34796 8968 34848 8974
rect 34900 8956 34928 9030
rect 34980 8968 35032 8974
rect 34900 8928 34980 8956
rect 34796 8910 34848 8916
rect 34980 8910 35032 8916
rect 34610 8256 34666 8265
rect 34610 8191 34666 8200
rect 34532 8078 34684 8106
rect 34656 8004 34684 8078
rect 34624 7976 34684 8004
rect 34428 7948 34480 7954
rect 34428 7890 34480 7896
rect 34624 7834 34652 7976
rect 34716 7886 34744 8910
rect 34808 8514 34836 8910
rect 35084 8820 35112 9132
rect 34992 8792 35112 8820
rect 35164 8832 35216 8838
rect 34886 8528 34942 8537
rect 34808 8486 34886 8514
rect 34886 8463 34942 8472
rect 34888 8424 34940 8430
rect 34888 8366 34940 8372
rect 34900 8294 34928 8366
rect 34992 8362 35020 8792
rect 35164 8774 35216 8780
rect 35072 8560 35124 8566
rect 35072 8502 35124 8508
rect 35084 8362 35112 8502
rect 35176 8498 35204 8774
rect 35254 8664 35310 8673
rect 35360 8650 35388 10934
rect 35544 10826 35572 11047
rect 35452 10798 35572 10826
rect 35452 9976 35480 10798
rect 35532 10668 35584 10674
rect 35532 10610 35584 10616
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35544 10441 35572 10610
rect 35636 10538 35664 10610
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 35530 10432 35586 10441
rect 35530 10367 35586 10376
rect 35728 10305 35756 12174
rect 35820 11218 35848 12174
rect 35808 11212 35860 11218
rect 35808 11154 35860 11160
rect 35806 11112 35862 11121
rect 35806 11047 35862 11056
rect 35820 10606 35848 11047
rect 35912 10606 35940 13280
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 36096 12442 36124 12786
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 36096 12306 36124 12378
rect 36280 12374 36308 13398
rect 36268 12368 36320 12374
rect 36268 12310 36320 12316
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 36176 11824 36228 11830
rect 36176 11766 36228 11772
rect 36266 11792 36322 11801
rect 36084 11688 36136 11694
rect 36084 11630 36136 11636
rect 36096 11529 36124 11630
rect 36082 11520 36138 11529
rect 36082 11455 36138 11464
rect 36188 11121 36216 11766
rect 36266 11727 36268 11736
rect 36320 11727 36322 11736
rect 36268 11698 36320 11704
rect 36268 11620 36320 11626
rect 36268 11562 36320 11568
rect 36280 11393 36308 11562
rect 36266 11384 36322 11393
rect 36266 11319 36322 11328
rect 36174 11112 36230 11121
rect 36174 11047 36230 11056
rect 35992 11008 36044 11014
rect 35992 10950 36044 10956
rect 36082 10976 36138 10985
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 35808 10464 35860 10470
rect 35808 10406 35860 10412
rect 35714 10296 35770 10305
rect 35820 10266 35848 10406
rect 35714 10231 35770 10240
rect 35808 10260 35860 10266
rect 35452 9948 35572 9976
rect 35438 9888 35494 9897
rect 35438 9823 35494 9832
rect 35452 9586 35480 9823
rect 35440 9580 35492 9586
rect 35440 9522 35492 9528
rect 35440 9444 35492 9450
rect 35440 9386 35492 9392
rect 35452 8974 35480 9386
rect 35544 9160 35572 9948
rect 35624 9376 35676 9382
rect 35622 9344 35624 9353
rect 35676 9344 35678 9353
rect 35622 9279 35678 9288
rect 35544 9132 35616 9160
rect 35588 9058 35616 9132
rect 35549 9030 35616 9058
rect 35549 9024 35577 9030
rect 35544 8996 35577 9024
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35440 8832 35492 8838
rect 35440 8774 35492 8780
rect 35310 8622 35388 8650
rect 35254 8599 35310 8608
rect 35346 8528 35402 8537
rect 35164 8492 35216 8498
rect 35346 8463 35402 8472
rect 35164 8434 35216 8440
rect 34980 8356 35032 8362
rect 34980 8298 35032 8304
rect 35072 8356 35124 8362
rect 35072 8298 35124 8304
rect 34808 8266 34928 8294
rect 34152 7812 34204 7818
rect 34152 7754 34204 7760
rect 34440 7806 34652 7834
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34150 7168 34206 7177
rect 34150 7103 34206 7112
rect 34164 7002 34192 7103
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34256 6866 34284 7346
rect 34440 7342 34468 7806
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 34428 7336 34480 7342
rect 34428 7278 34480 7284
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 34256 6390 34284 6802
rect 34244 6384 34296 6390
rect 34244 6326 34296 6332
rect 34152 6248 34204 6254
rect 34152 6190 34204 6196
rect 34060 6180 34112 6186
rect 34060 6122 34112 6128
rect 33966 5808 34022 5817
rect 33966 5743 34022 5752
rect 33784 5228 33836 5234
rect 34164 5216 34192 6190
rect 34244 5228 34296 5234
rect 34164 5188 34244 5216
rect 33784 5170 33836 5176
rect 34244 5170 34296 5176
rect 33796 4826 33824 5170
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 33612 4440 33732 4468
rect 33506 4176 33562 4185
rect 33506 4111 33508 4120
rect 33560 4111 33562 4120
rect 33508 4082 33560 4088
rect 33612 4026 33640 4440
rect 33692 4140 33744 4146
rect 33692 4082 33744 4088
rect 33520 3998 33640 4026
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33416 2100 33468 2106
rect 33416 2042 33468 2048
rect 33322 912 33378 921
rect 33322 847 33378 856
rect 33428 800 33456 2042
rect 33520 1222 33548 3998
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33612 2310 33640 2586
rect 33600 2304 33652 2310
rect 33600 2246 33652 2252
rect 33508 1216 33560 1222
rect 33508 1158 33560 1164
rect 33704 800 33732 4082
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 33784 2372 33836 2378
rect 33784 2314 33836 2320
rect 33796 1426 33824 2314
rect 33784 1420 33836 1426
rect 33784 1362 33836 1368
rect 33980 800 34008 3062
rect 34072 2446 34100 5102
rect 34244 4480 34296 4486
rect 34244 4422 34296 4428
rect 34256 3738 34284 4422
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34150 3224 34206 3233
rect 34150 3159 34206 3168
rect 34164 3058 34192 3159
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 34348 2650 34376 7278
rect 34440 6186 34468 7278
rect 34532 6474 34560 7686
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34610 7032 34666 7041
rect 34610 6967 34666 6976
rect 34624 6730 34652 6967
rect 34716 6905 34744 7414
rect 34702 6896 34758 6905
rect 34808 6866 34836 8266
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35072 8084 35124 8090
rect 35072 8026 35124 8032
rect 35084 7886 35112 8026
rect 35360 8022 35388 8463
rect 35256 8016 35308 8022
rect 35256 7958 35308 7964
rect 35348 8016 35400 8022
rect 35348 7958 35400 7964
rect 35072 7880 35124 7886
rect 35268 7878 35296 7958
rect 35452 7878 35480 8774
rect 35268 7850 35480 7878
rect 35072 7822 35124 7828
rect 35348 7812 35400 7818
rect 35348 7754 35400 7760
rect 35254 7440 35310 7449
rect 35254 7375 35256 7384
rect 35308 7375 35310 7384
rect 35256 7346 35308 7352
rect 35360 7177 35388 7754
rect 35440 7472 35492 7478
rect 35544 7460 35572 8996
rect 35624 8968 35676 8974
rect 35624 8910 35676 8916
rect 35636 8412 35664 8910
rect 35728 8514 35756 10231
rect 35808 10202 35860 10208
rect 35900 10192 35952 10198
rect 35900 10134 35952 10140
rect 35806 9616 35862 9625
rect 35806 9551 35808 9560
rect 35860 9551 35862 9560
rect 35808 9522 35860 9528
rect 35912 9432 35940 10134
rect 36004 9897 36032 10950
rect 36082 10911 36138 10920
rect 36096 10282 36124 10911
rect 36188 10606 36216 11047
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 36176 10600 36228 10606
rect 36176 10542 36228 10548
rect 36280 10282 36308 10610
rect 36096 10254 36308 10282
rect 36268 10192 36320 10198
rect 36268 10134 36320 10140
rect 36176 10056 36228 10062
rect 36176 9998 36228 10004
rect 36188 9897 36216 9998
rect 35990 9888 36046 9897
rect 35990 9823 36046 9832
rect 36174 9888 36230 9897
rect 36174 9823 36230 9832
rect 36084 9580 36136 9586
rect 36084 9522 36136 9528
rect 36096 9489 36124 9522
rect 36082 9480 36138 9489
rect 35992 9444 36044 9450
rect 35912 9404 35992 9432
rect 36082 9415 36138 9424
rect 35992 9386 36044 9392
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 35990 9344 36046 9353
rect 35820 9110 35848 9318
rect 35990 9279 36046 9288
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 36004 8974 36032 9279
rect 35992 8968 36044 8974
rect 35992 8910 36044 8916
rect 35728 8486 35848 8514
rect 35716 8424 35768 8430
rect 35636 8384 35716 8412
rect 35716 8366 35768 8372
rect 35492 7432 35572 7460
rect 35440 7414 35492 7420
rect 35346 7168 35402 7177
rect 34934 7100 35242 7109
rect 35346 7103 35402 7112
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35728 7002 35756 8366
rect 35820 8294 35848 8486
rect 35808 8288 35860 8294
rect 35808 8230 35860 8236
rect 35806 8120 35862 8129
rect 35806 8055 35862 8064
rect 35820 7970 35848 8055
rect 35820 7942 35940 7970
rect 35912 7546 35940 7942
rect 35900 7540 35952 7546
rect 35900 7482 35952 7488
rect 36004 7426 36032 8910
rect 36096 8566 36124 9415
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 36280 8498 36308 10134
rect 36372 9092 36400 14350
rect 36464 13025 36492 14894
rect 36450 13016 36506 13025
rect 36450 12951 36506 12960
rect 36464 12918 36492 12951
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36556 12850 36584 17070
rect 36636 15360 36688 15366
rect 36636 15302 36688 15308
rect 36648 15162 36676 15302
rect 36636 15156 36688 15162
rect 36636 15098 36688 15104
rect 36634 15056 36690 15065
rect 36634 14991 36690 15000
rect 36648 14958 36676 14991
rect 36636 14952 36688 14958
rect 36636 14894 36688 14900
rect 36634 14648 36690 14657
rect 36634 14583 36690 14592
rect 36648 14550 36676 14583
rect 36636 14544 36688 14550
rect 36636 14486 36688 14492
rect 36636 14340 36688 14346
rect 36636 14282 36688 14288
rect 36544 12844 36596 12850
rect 36544 12786 36596 12792
rect 36544 12436 36596 12442
rect 36544 12378 36596 12384
rect 36452 12232 36504 12238
rect 36452 12174 36504 12180
rect 36464 10810 36492 12174
rect 36452 10804 36504 10810
rect 36452 10746 36504 10752
rect 36452 10464 36504 10470
rect 36452 10406 36504 10412
rect 36464 9994 36492 10406
rect 36452 9988 36504 9994
rect 36452 9930 36504 9936
rect 36556 9586 36584 12378
rect 36648 11257 36676 14282
rect 36740 11286 36768 22066
rect 36820 19712 36872 19718
rect 36820 19654 36872 19660
rect 36832 17610 36860 19654
rect 36820 17604 36872 17610
rect 36820 17546 36872 17552
rect 36912 16992 36964 16998
rect 36912 16934 36964 16940
rect 36924 16017 36952 16934
rect 36910 16008 36966 16017
rect 36910 15943 36966 15952
rect 36912 15564 36964 15570
rect 36912 15506 36964 15512
rect 36820 15020 36872 15026
rect 36820 14962 36872 14968
rect 36832 13433 36860 14962
rect 36924 14113 36952 15506
rect 36910 14104 36966 14113
rect 36910 14039 36966 14048
rect 36818 13424 36874 13433
rect 36818 13359 36874 13368
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36832 11830 36860 12786
rect 36820 11824 36872 11830
rect 36820 11766 36872 11772
rect 36728 11280 36780 11286
rect 36634 11248 36690 11257
rect 36728 11222 36780 11228
rect 36634 11183 36690 11192
rect 36740 11082 36768 11222
rect 36912 11144 36964 11150
rect 36912 11086 36964 11092
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36634 10976 36690 10985
rect 36634 10911 36690 10920
rect 36648 10130 36676 10911
rect 36728 10804 36780 10810
rect 36728 10746 36780 10752
rect 36636 10124 36688 10130
rect 36636 10066 36688 10072
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36636 9580 36688 9586
rect 36636 9522 36688 9528
rect 36648 9330 36676 9522
rect 36556 9302 36676 9330
rect 36556 9217 36584 9302
rect 36542 9208 36598 9217
rect 36740 9194 36768 10746
rect 36924 10538 36952 11086
rect 36912 10532 36964 10538
rect 36912 10474 36964 10480
rect 36910 9888 36966 9897
rect 36910 9823 36966 9832
rect 36924 9586 36952 9823
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 36924 9364 36952 9522
rect 36542 9143 36598 9152
rect 36648 9166 36768 9194
rect 36832 9336 36952 9364
rect 36372 9064 36584 9092
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 36358 8256 36414 8265
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36096 7546 36124 8026
rect 36188 7886 36216 8230
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 35912 7398 36032 7426
rect 35820 7177 35848 7346
rect 35806 7168 35862 7177
rect 35806 7103 35862 7112
rect 35256 6996 35308 7002
rect 35256 6938 35308 6944
rect 35716 6996 35768 7002
rect 35716 6938 35768 6944
rect 34888 6928 34940 6934
rect 34886 6896 34888 6905
rect 34940 6896 34942 6905
rect 34702 6831 34758 6840
rect 34796 6860 34848 6866
rect 34886 6831 34942 6840
rect 34796 6802 34848 6808
rect 34612 6724 34664 6730
rect 34612 6666 34664 6672
rect 34532 6446 34744 6474
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34428 6180 34480 6186
rect 34428 6122 34480 6128
rect 34440 5030 34468 6122
rect 34532 5953 34560 6258
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34624 6089 34652 6190
rect 34716 6118 34744 6446
rect 35268 6390 35296 6938
rect 35530 6896 35586 6905
rect 35360 6854 35530 6882
rect 35360 6798 35388 6854
rect 35530 6831 35586 6840
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 34796 6384 34848 6390
rect 34796 6326 34848 6332
rect 35256 6384 35308 6390
rect 35256 6326 35308 6332
rect 34704 6112 34756 6118
rect 34610 6080 34666 6089
rect 34704 6054 34756 6060
rect 34610 6015 34666 6024
rect 34518 5944 34574 5953
rect 34518 5879 34574 5888
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34426 4720 34482 4729
rect 34426 4655 34482 4664
rect 34440 4554 34468 4655
rect 34428 4548 34480 4554
rect 34428 4490 34480 4496
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34440 3058 34468 3674
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 34336 2644 34388 2650
rect 34336 2586 34388 2592
rect 34060 2440 34112 2446
rect 34244 2440 34296 2446
rect 34060 2382 34112 2388
rect 34164 2400 34244 2428
rect 34164 2038 34192 2400
rect 34244 2382 34296 2388
rect 34152 2032 34204 2038
rect 34152 1974 34204 1980
rect 34244 2032 34296 2038
rect 34244 1974 34296 1980
rect 34256 800 34284 1974
rect 34532 800 34560 5578
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 34624 4690 34652 5510
rect 34808 5030 34836 6326
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35176 6100 35204 6258
rect 35176 6072 35296 6100
rect 35544 6089 35572 6258
rect 35636 6254 35664 6802
rect 35716 6792 35768 6798
rect 35716 6734 35768 6740
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35268 6066 35296 6072
rect 35530 6080 35586 6089
rect 35268 6038 35388 6066
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34980 5840 35032 5846
rect 34980 5782 35032 5788
rect 34992 5710 35020 5782
rect 34980 5704 35032 5710
rect 34980 5646 35032 5652
rect 35360 5370 35388 6038
rect 35530 6015 35586 6024
rect 35624 5840 35676 5846
rect 35624 5782 35676 5788
rect 35532 5772 35584 5778
rect 35532 5714 35584 5720
rect 35438 5400 35494 5409
rect 35348 5364 35400 5370
rect 35438 5335 35494 5344
rect 35348 5306 35400 5312
rect 35072 5228 35124 5234
rect 35072 5170 35124 5176
rect 35084 5098 35112 5170
rect 35348 5160 35400 5166
rect 35348 5102 35400 5108
rect 35072 5092 35124 5098
rect 35072 5034 35124 5040
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34612 4684 34664 4690
rect 34612 4626 34664 4632
rect 35360 4146 35388 5102
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 34796 4004 34848 4010
rect 34796 3946 34848 3952
rect 34808 800 34836 3946
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34888 3596 34940 3602
rect 34888 3538 34940 3544
rect 34900 3058 34928 3538
rect 35256 3392 35308 3398
rect 35256 3334 35308 3340
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 35268 2938 35296 3334
rect 35360 3126 35388 3878
rect 35452 3369 35480 5335
rect 35544 4729 35572 5714
rect 35530 4720 35586 4729
rect 35530 4655 35532 4664
rect 35584 4655 35586 4664
rect 35532 4626 35584 4632
rect 35636 4026 35664 5782
rect 35728 4214 35756 6734
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 35820 5234 35848 6258
rect 35912 5778 35940 7398
rect 35992 7336 36044 7342
rect 35992 7278 36044 7284
rect 36004 7002 36032 7278
rect 36280 7274 36308 8230
rect 36358 8191 36414 8200
rect 36372 7313 36400 8191
rect 36358 7304 36414 7313
rect 36084 7268 36136 7274
rect 36084 7210 36136 7216
rect 36268 7268 36320 7274
rect 36358 7239 36414 7248
rect 36268 7210 36320 7216
rect 36096 7002 36124 7210
rect 35992 6996 36044 7002
rect 35992 6938 36044 6944
rect 36084 6996 36136 7002
rect 36084 6938 36136 6944
rect 36084 6792 36136 6798
rect 36360 6792 36412 6798
rect 36136 6740 36216 6746
rect 36084 6734 36216 6740
rect 36360 6734 36412 6740
rect 35992 6724 36044 6730
rect 36096 6718 36216 6734
rect 35992 6666 36044 6672
rect 36004 6186 36032 6666
rect 36084 6656 36136 6662
rect 36188 6633 36216 6718
rect 36268 6656 36320 6662
rect 36084 6598 36136 6604
rect 36174 6624 36230 6633
rect 35992 6180 36044 6186
rect 35992 6122 36044 6128
rect 36096 5794 36124 6598
rect 36268 6598 36320 6604
rect 36174 6559 36230 6568
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 36188 6118 36216 6394
rect 36280 6390 36308 6598
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 36372 6322 36400 6734
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 36176 6112 36228 6118
rect 36176 6054 36228 6060
rect 35900 5772 35952 5778
rect 36096 5766 36308 5794
rect 35900 5714 35952 5720
rect 35808 5228 35860 5234
rect 35808 5170 35860 5176
rect 35820 4570 35848 5170
rect 35912 5166 35940 5714
rect 36280 5710 36308 5766
rect 36268 5704 36320 5710
rect 36174 5672 36230 5681
rect 36268 5646 36320 5652
rect 36174 5607 36230 5616
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35900 5160 35952 5166
rect 35898 5128 35900 5137
rect 35952 5128 35954 5137
rect 35898 5063 35954 5072
rect 36096 4758 36124 5306
rect 36188 5234 36216 5607
rect 36464 5370 36492 8434
rect 36556 7177 36584 9064
rect 36542 7168 36598 7177
rect 36542 7103 36598 7112
rect 36544 6656 36596 6662
rect 36544 6598 36596 6604
rect 36556 6458 36584 6598
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36648 5250 36676 9166
rect 36728 7948 36780 7954
rect 36728 7890 36780 7896
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 36372 5222 36676 5250
rect 36266 4856 36322 4865
rect 36266 4791 36322 4800
rect 36084 4752 36136 4758
rect 36084 4694 36136 4700
rect 36176 4616 36228 4622
rect 35820 4542 36032 4570
rect 36176 4558 36228 4564
rect 36004 4486 36032 4542
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 35912 4282 35940 4422
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35716 4208 35768 4214
rect 35716 4150 35768 4156
rect 35898 4176 35954 4185
rect 35898 4111 35954 4120
rect 35912 4078 35940 4111
rect 35900 4072 35952 4078
rect 35636 3998 35756 4026
rect 35900 4014 35952 4020
rect 35624 3936 35676 3942
rect 35728 3913 35756 3998
rect 35624 3878 35676 3884
rect 35714 3904 35770 3913
rect 35438 3360 35494 3369
rect 35438 3295 35494 3304
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35268 2910 35388 2938
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35256 2372 35308 2378
rect 35256 2314 35308 2320
rect 35268 2106 35296 2314
rect 35256 2100 35308 2106
rect 35256 2042 35308 2048
rect 35360 1442 35388 2910
rect 35084 1414 35388 1442
rect 35084 800 35112 1414
rect 35452 1034 35480 3062
rect 35360 1006 35480 1034
rect 35360 800 35388 1006
rect 35636 800 35664 3878
rect 35714 3839 35770 3848
rect 35898 3768 35954 3777
rect 36188 3738 36216 4558
rect 36280 4321 36308 4791
rect 36266 4312 36322 4321
rect 36266 4247 36322 4256
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 35898 3703 35900 3712
rect 35952 3703 35954 3712
rect 36176 3732 36228 3738
rect 35900 3674 35952 3680
rect 36176 3674 36228 3680
rect 36084 3664 36136 3670
rect 36084 3606 36136 3612
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 35912 800 35940 3538
rect 36096 3534 36124 3606
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 36084 3188 36136 3194
rect 36084 3130 36136 3136
rect 36096 2514 36124 3130
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 36188 1578 36216 3674
rect 36280 3194 36308 4082
rect 36372 4078 36400 5222
rect 36544 5024 36596 5030
rect 36544 4966 36596 4972
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 36556 4622 36584 4966
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 36360 4072 36412 4078
rect 36360 4014 36412 4020
rect 36464 3738 36492 4082
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36648 3466 36676 4966
rect 36740 4282 36768 7890
rect 36832 5273 36860 9336
rect 36912 8560 36964 8566
rect 36910 8528 36912 8537
rect 36964 8528 36966 8537
rect 36910 8463 36966 8472
rect 37016 8090 37044 35158
rect 37384 35018 37412 42638
rect 37372 35012 37424 35018
rect 37372 34954 37424 34960
rect 37384 34746 37412 34954
rect 37372 34740 37424 34746
rect 37372 34682 37424 34688
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37372 19780 37424 19786
rect 37372 19722 37424 19728
rect 37384 19378 37412 19722
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37096 19304 37148 19310
rect 37096 19246 37148 19252
rect 37108 14618 37136 19246
rect 37476 18426 37504 19790
rect 37188 18420 37240 18426
rect 37188 18362 37240 18368
rect 37464 18420 37516 18426
rect 37464 18362 37516 18368
rect 37200 17202 37228 18362
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 37292 17542 37320 18226
rect 37556 18148 37608 18154
rect 37556 18090 37608 18096
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37280 17536 37332 17542
rect 37280 17478 37332 17484
rect 37188 17196 37240 17202
rect 37188 17138 37240 17144
rect 37186 16688 37242 16697
rect 37186 16623 37242 16632
rect 37200 16402 37228 16623
rect 37292 16590 37320 17478
rect 37280 16584 37332 16590
rect 37280 16526 37332 16532
rect 37200 16374 37320 16402
rect 37188 15972 37240 15978
rect 37188 15914 37240 15920
rect 37200 14958 37228 15914
rect 37188 14952 37240 14958
rect 37188 14894 37240 14900
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 37108 14074 37136 14554
rect 37188 14544 37240 14550
rect 37188 14486 37240 14492
rect 37096 14068 37148 14074
rect 37096 14010 37148 14016
rect 37200 13977 37228 14486
rect 37186 13968 37242 13977
rect 37292 13938 37320 16374
rect 37384 14074 37412 17546
rect 37476 16114 37504 17614
rect 37568 16697 37596 18090
rect 37660 17542 37688 44814
rect 38568 41472 38620 41478
rect 38568 41414 38620 41420
rect 38580 40118 38608 41414
rect 38568 40112 38620 40118
rect 38568 40054 38620 40060
rect 38568 38752 38620 38758
rect 38568 38694 38620 38700
rect 38016 38004 38068 38010
rect 38016 37946 38068 37952
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 37740 19780 37792 19786
rect 37740 19722 37792 19728
rect 37648 17536 37700 17542
rect 37648 17478 37700 17484
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37554 16688 37610 16697
rect 37554 16623 37610 16632
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37476 15094 37504 16050
rect 37568 15638 37596 16050
rect 37556 15632 37608 15638
rect 37556 15574 37608 15580
rect 37464 15088 37516 15094
rect 37464 15030 37516 15036
rect 37660 15026 37688 17138
rect 37752 16017 37780 19722
rect 37936 18222 37964 24550
rect 38028 20777 38056 37946
rect 38580 36106 38608 38694
rect 38568 36100 38620 36106
rect 38568 36042 38620 36048
rect 38844 33312 38896 33318
rect 38844 33254 38896 33260
rect 38476 22432 38528 22438
rect 38476 22374 38528 22380
rect 38014 20768 38070 20777
rect 38014 20703 38070 20712
rect 38384 20392 38436 20398
rect 38384 20334 38436 20340
rect 38108 18828 38160 18834
rect 38108 18770 38160 18776
rect 37924 18216 37976 18222
rect 37924 18158 37976 18164
rect 37832 16992 37884 16998
rect 37832 16934 37884 16940
rect 37738 16008 37794 16017
rect 37738 15943 37794 15952
rect 37740 15904 37792 15910
rect 37740 15846 37792 15852
rect 37752 15502 37780 15846
rect 37740 15496 37792 15502
rect 37738 15464 37740 15473
rect 37792 15464 37794 15473
rect 37738 15399 37794 15408
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37554 14648 37610 14657
rect 37554 14583 37556 14592
rect 37608 14583 37610 14592
rect 37556 14554 37608 14560
rect 37464 14340 37516 14346
rect 37464 14282 37516 14288
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37186 13903 37242 13912
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 37476 13870 37504 14282
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 37464 13864 37516 13870
rect 37464 13806 37516 13812
rect 37094 13560 37150 13569
rect 37094 13495 37150 13504
rect 37108 13462 37136 13495
rect 37096 13456 37148 13462
rect 37096 13398 37148 13404
rect 37280 13320 37332 13326
rect 37280 13262 37332 13268
rect 37096 12912 37148 12918
rect 37096 12854 37148 12860
rect 37108 11286 37136 12854
rect 37292 12714 37320 13262
rect 37372 12776 37424 12782
rect 37372 12718 37424 12724
rect 37280 12708 37332 12714
rect 37280 12650 37332 12656
rect 37280 12368 37332 12374
rect 37280 12310 37332 12316
rect 37292 11762 37320 12310
rect 37280 11756 37332 11762
rect 37280 11698 37332 11704
rect 37384 11694 37412 12718
rect 37568 12209 37596 13874
rect 37660 13841 37688 14962
rect 37740 14408 37792 14414
rect 37740 14350 37792 14356
rect 37646 13832 37702 13841
rect 37646 13767 37702 13776
rect 37752 13705 37780 14350
rect 37738 13696 37794 13705
rect 37738 13631 37794 13640
rect 37740 13456 37792 13462
rect 37740 13398 37792 13404
rect 37752 13326 37780 13398
rect 37740 13320 37792 13326
rect 37738 13288 37740 13297
rect 37792 13288 37794 13297
rect 37738 13223 37794 13232
rect 37740 12776 37792 12782
rect 37740 12718 37792 12724
rect 37648 12368 37700 12374
rect 37648 12310 37700 12316
rect 37554 12200 37610 12209
rect 37476 12158 37554 12186
rect 37372 11688 37424 11694
rect 37372 11630 37424 11636
rect 37370 11384 37426 11393
rect 37188 11348 37240 11354
rect 37370 11319 37372 11328
rect 37188 11290 37240 11296
rect 37424 11319 37426 11328
rect 37372 11290 37424 11296
rect 37096 11280 37148 11286
rect 37096 11222 37148 11228
rect 37200 11150 37228 11290
rect 37280 11280 37332 11286
rect 37280 11222 37332 11228
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37188 11008 37240 11014
rect 37188 10950 37240 10956
rect 37096 10056 37148 10062
rect 37096 9998 37148 10004
rect 37108 9042 37136 9998
rect 37200 9353 37228 10950
rect 37186 9344 37242 9353
rect 37186 9279 37242 9288
rect 37188 9104 37240 9110
rect 37188 9046 37240 9052
rect 37096 9036 37148 9042
rect 37096 8978 37148 8984
rect 37108 8498 37136 8978
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 37004 8084 37056 8090
rect 37004 8026 37056 8032
rect 36912 8016 36964 8022
rect 36912 7958 36964 7964
rect 36924 7546 36952 7958
rect 37004 7744 37056 7750
rect 37004 7686 37056 7692
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 37016 7478 37044 7686
rect 37004 7472 37056 7478
rect 37004 7414 37056 7420
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 36912 6928 36964 6934
rect 36912 6870 36964 6876
rect 36924 6089 36952 6870
rect 37016 6798 37044 7210
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 37004 6656 37056 6662
rect 37002 6624 37004 6633
rect 37056 6624 37058 6633
rect 37002 6559 37058 6568
rect 37108 6322 37136 8434
rect 37200 8362 37228 9046
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37292 8265 37320 11222
rect 37372 11008 37424 11014
rect 37372 10950 37424 10956
rect 37384 10606 37412 10950
rect 37372 10600 37424 10606
rect 37372 10542 37424 10548
rect 37372 10464 37424 10470
rect 37372 10406 37424 10412
rect 37384 10062 37412 10406
rect 37372 10056 37424 10062
rect 37372 9998 37424 10004
rect 37476 8650 37504 12158
rect 37554 12135 37610 12144
rect 37660 10810 37688 12310
rect 37752 11354 37780 12718
rect 37740 11348 37792 11354
rect 37740 11290 37792 11296
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 37554 10160 37610 10169
rect 37554 10095 37610 10104
rect 37568 8906 37596 10095
rect 37844 9738 37872 16934
rect 37936 12238 37964 18158
rect 38120 17785 38148 18770
rect 38106 17776 38162 17785
rect 38106 17711 38162 17720
rect 38120 16250 38148 17711
rect 38292 16992 38344 16998
rect 38292 16934 38344 16940
rect 38304 16726 38332 16934
rect 38292 16720 38344 16726
rect 38292 16662 38344 16668
rect 38200 16652 38252 16658
rect 38200 16594 38252 16600
rect 38108 16244 38160 16250
rect 38108 16186 38160 16192
rect 38120 15570 38148 16186
rect 38212 16114 38240 16594
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38108 15564 38160 15570
rect 38108 15506 38160 15512
rect 38016 15088 38068 15094
rect 38016 15030 38068 15036
rect 38028 14482 38056 15030
rect 38120 14958 38148 15506
rect 38108 14952 38160 14958
rect 38108 14894 38160 14900
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 38028 13938 38056 14418
rect 38016 13932 38068 13938
rect 38016 13874 38068 13880
rect 38016 12300 38068 12306
rect 38016 12242 38068 12248
rect 37924 12232 37976 12238
rect 37924 12174 37976 12180
rect 38028 11286 38056 12242
rect 38120 12238 38148 14894
rect 38198 13832 38254 13841
rect 38198 13767 38254 13776
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38212 11880 38240 13767
rect 38396 13530 38424 20334
rect 38488 16658 38516 22374
rect 38856 22094 38884 33254
rect 39488 28484 39540 28490
rect 39488 28426 39540 28432
rect 38856 22066 38976 22094
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38764 20058 38792 20402
rect 38752 20052 38804 20058
rect 38752 19994 38804 20000
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38856 18766 38884 19654
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38568 18624 38620 18630
rect 38568 18566 38620 18572
rect 38580 17610 38608 18566
rect 38856 18426 38884 18702
rect 38844 18420 38896 18426
rect 38844 18362 38896 18368
rect 38660 18216 38712 18222
rect 38660 18158 38712 18164
rect 38672 17678 38700 18158
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 38568 17604 38620 17610
rect 38568 17546 38620 17552
rect 38672 17338 38700 17614
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 38752 16720 38804 16726
rect 38752 16662 38804 16668
rect 38476 16652 38528 16658
rect 38476 16594 38528 16600
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 38396 13326 38424 13466
rect 38384 13320 38436 13326
rect 38120 11852 38240 11880
rect 38304 13280 38384 13308
rect 38016 11280 38068 11286
rect 38016 11222 38068 11228
rect 38016 11144 38068 11150
rect 38016 11086 38068 11092
rect 37924 10600 37976 10606
rect 37924 10542 37976 10548
rect 37936 9926 37964 10542
rect 37924 9920 37976 9926
rect 37924 9862 37976 9868
rect 38028 9761 38056 11086
rect 38120 10985 38148 11852
rect 38304 11218 38332 13280
rect 38384 13262 38436 13268
rect 38292 11212 38344 11218
rect 38292 11154 38344 11160
rect 38106 10976 38162 10985
rect 38106 10911 38162 10920
rect 38106 10432 38162 10441
rect 38106 10367 38162 10376
rect 38120 10198 38148 10367
rect 38108 10192 38160 10198
rect 38108 10134 38160 10140
rect 37752 9710 37872 9738
rect 38014 9752 38070 9761
rect 37556 8900 37608 8906
rect 37556 8842 37608 8848
rect 37384 8622 37504 8650
rect 37278 8256 37334 8265
rect 37278 8191 37334 8200
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37292 7818 37320 8026
rect 37384 8022 37412 8622
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 37384 7818 37412 7958
rect 37280 7812 37332 7818
rect 37280 7754 37332 7760
rect 37372 7812 37424 7818
rect 37372 7754 37424 7760
rect 37292 7698 37320 7754
rect 37292 7670 37412 7698
rect 37280 7404 37332 7410
rect 37280 7346 37332 7352
rect 37188 7336 37240 7342
rect 37188 7278 37240 7284
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 36910 6080 36966 6089
rect 36910 6015 36966 6024
rect 36818 5264 36874 5273
rect 36818 5199 36874 5208
rect 36924 4434 36952 6015
rect 37016 4554 37044 6258
rect 37200 6254 37228 7278
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 37096 5772 37148 5778
rect 37096 5714 37148 5720
rect 37108 4826 37136 5714
rect 37188 5568 37240 5574
rect 37188 5510 37240 5516
rect 37096 4820 37148 4826
rect 37096 4762 37148 4768
rect 37004 4548 37056 4554
rect 37004 4490 37056 4496
rect 36924 4406 37136 4434
rect 36728 4276 36780 4282
rect 36728 4218 36780 4224
rect 37004 4140 37056 4146
rect 37004 4082 37056 4088
rect 36726 4040 36782 4049
rect 36726 3975 36782 3984
rect 36740 3534 36768 3975
rect 36910 3632 36966 3641
rect 37016 3602 37044 4082
rect 36910 3567 36966 3576
rect 37004 3596 37056 3602
rect 36924 3534 36952 3567
rect 37004 3538 37056 3544
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 36912 3528 36964 3534
rect 36912 3470 36964 3476
rect 36636 3460 36688 3466
rect 36636 3402 36688 3408
rect 37004 3460 37056 3466
rect 37108 3448 37136 4406
rect 37200 3670 37228 5510
rect 37292 3670 37320 7346
rect 37384 6338 37412 7670
rect 37476 7410 37504 8502
rect 37568 8090 37596 8842
rect 37648 8832 37700 8838
rect 37648 8774 37700 8780
rect 37660 8634 37688 8774
rect 37648 8628 37700 8634
rect 37648 8570 37700 8576
rect 37556 8084 37608 8090
rect 37556 8026 37608 8032
rect 37648 8016 37700 8022
rect 37648 7958 37700 7964
rect 37556 7744 37608 7750
rect 37556 7686 37608 7692
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 37568 6905 37596 7686
rect 37660 7041 37688 7958
rect 37752 7886 37780 9710
rect 38014 9687 38070 9696
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 37844 9178 37872 9522
rect 37832 9172 37884 9178
rect 37832 9114 37884 9120
rect 37844 9042 37872 9114
rect 37832 9036 37884 9042
rect 37832 8978 37884 8984
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 37924 8900 37976 8906
rect 37924 8842 37976 8848
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 37740 7404 37792 7410
rect 37740 7346 37792 7352
rect 37646 7032 37702 7041
rect 37646 6967 37702 6976
rect 37554 6896 37610 6905
rect 37554 6831 37610 6840
rect 37648 6860 37700 6866
rect 37648 6802 37700 6808
rect 37384 6310 37596 6338
rect 37370 6216 37426 6225
rect 37370 6151 37426 6160
rect 37384 5778 37412 6151
rect 37372 5772 37424 5778
rect 37372 5714 37424 5720
rect 37372 5160 37424 5166
rect 37372 5102 37424 5108
rect 37188 3664 37240 3670
rect 37188 3606 37240 3612
rect 37280 3664 37332 3670
rect 37280 3606 37332 3612
rect 37056 3420 37136 3448
rect 37004 3402 37056 3408
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 36452 3188 36504 3194
rect 36452 3130 36504 3136
rect 36096 1550 36216 1578
rect 36096 1193 36124 1550
rect 36464 1442 36492 3130
rect 36544 2916 36596 2922
rect 36544 2858 36596 2864
rect 36188 1414 36492 1442
rect 36082 1184 36138 1193
rect 36082 1119 36138 1128
rect 36188 800 36216 1414
rect 36556 1306 36584 2858
rect 37004 2848 37056 2854
rect 37004 2790 37056 2796
rect 36728 2100 36780 2106
rect 36728 2042 36780 2048
rect 36464 1278 36584 1306
rect 36464 800 36492 1278
rect 36740 800 36768 2042
rect 37016 800 37044 2790
rect 37384 2774 37412 5102
rect 37568 4622 37596 6310
rect 37660 5914 37688 6802
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37752 5556 37780 7346
rect 37844 7342 37872 8230
rect 37832 7336 37884 7342
rect 37832 7278 37884 7284
rect 37832 6928 37884 6934
rect 37936 6916 37964 8842
rect 38028 8090 38056 8910
rect 38016 8084 38068 8090
rect 38016 8026 38068 8032
rect 37884 6888 37964 6916
rect 38120 6882 38148 8910
rect 38198 8256 38254 8265
rect 38198 8191 38254 8200
rect 38212 7410 38240 8191
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38304 7342 38332 11154
rect 38488 10810 38516 16594
rect 38660 16040 38712 16046
rect 38660 15982 38712 15988
rect 38672 14278 38700 15982
rect 38764 15366 38792 16662
rect 38842 15464 38898 15473
rect 38842 15399 38844 15408
rect 38896 15399 38898 15408
rect 38844 15370 38896 15376
rect 38752 15360 38804 15366
rect 38752 15302 38804 15308
rect 38842 15192 38898 15201
rect 38842 15127 38844 15136
rect 38896 15127 38898 15136
rect 38844 15098 38896 15104
rect 38750 15056 38806 15065
rect 38750 14991 38806 15000
rect 38764 14890 38792 14991
rect 38752 14884 38804 14890
rect 38752 14826 38804 14832
rect 38844 14816 38896 14822
rect 38844 14758 38896 14764
rect 38856 14414 38884 14758
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 38752 14340 38804 14346
rect 38752 14282 38804 14288
rect 38660 14272 38712 14278
rect 38660 14214 38712 14220
rect 38672 14074 38700 14214
rect 38764 14113 38792 14282
rect 38750 14104 38806 14113
rect 38660 14068 38712 14074
rect 38750 14039 38806 14048
rect 38660 14010 38712 14016
rect 38672 13258 38700 14010
rect 38660 13252 38712 13258
rect 38660 13194 38712 13200
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38566 12880 38622 12889
rect 38566 12815 38622 12824
rect 38580 11762 38608 12815
rect 38856 12238 38884 13194
rect 38948 12782 38976 22066
rect 39212 20392 39264 20398
rect 39212 20334 39264 20340
rect 39120 20324 39172 20330
rect 39120 20266 39172 20272
rect 39028 20256 39080 20262
rect 39028 20198 39080 20204
rect 39040 18290 39068 20198
rect 39028 18284 39080 18290
rect 39028 18226 39080 18232
rect 39028 17536 39080 17542
rect 39028 17478 39080 17484
rect 38936 12776 38988 12782
rect 38936 12718 38988 12724
rect 38844 12232 38896 12238
rect 38844 12174 38896 12180
rect 38568 11756 38620 11762
rect 38568 11698 38620 11704
rect 38568 11620 38620 11626
rect 38568 11562 38620 11568
rect 38580 11529 38608 11562
rect 38752 11552 38804 11558
rect 38566 11520 38622 11529
rect 38752 11494 38804 11500
rect 38844 11552 38896 11558
rect 38844 11494 38896 11500
rect 38566 11455 38622 11464
rect 38764 11150 38792 11494
rect 38856 11286 38884 11494
rect 38844 11280 38896 11286
rect 38844 11222 38896 11228
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38936 11076 38988 11082
rect 38936 11018 38988 11024
rect 38658 10976 38714 10985
rect 38658 10911 38714 10920
rect 38476 10804 38528 10810
rect 38476 10746 38528 10752
rect 38672 10674 38700 10911
rect 38660 10668 38712 10674
rect 38660 10610 38712 10616
rect 38752 10668 38804 10674
rect 38752 10610 38804 10616
rect 38672 10062 38700 10610
rect 38764 10305 38792 10610
rect 38948 10538 38976 11018
rect 38936 10532 38988 10538
rect 38936 10474 38988 10480
rect 38750 10296 38806 10305
rect 38750 10231 38806 10240
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38660 9920 38712 9926
rect 38660 9862 38712 9868
rect 38382 9616 38438 9625
rect 38672 9586 38700 9862
rect 38382 9551 38438 9560
rect 38660 9580 38712 9586
rect 38396 8974 38424 9551
rect 38660 9522 38712 9528
rect 38672 9489 38700 9522
rect 38658 9480 38714 9489
rect 38658 9415 38714 9424
rect 38660 9376 38712 9382
rect 38660 9318 38712 9324
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 38476 8968 38528 8974
rect 38476 8910 38528 8916
rect 38488 8566 38516 8910
rect 38476 8560 38528 8566
rect 38476 8502 38528 8508
rect 38488 7993 38516 8502
rect 38566 8256 38622 8265
rect 38566 8191 38622 8200
rect 38474 7984 38530 7993
rect 38474 7919 38530 7928
rect 38384 7880 38436 7886
rect 38384 7822 38436 7828
rect 38476 7880 38528 7886
rect 38476 7822 38528 7828
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 37832 6870 37884 6876
rect 38028 6854 38148 6882
rect 38304 6866 38332 7278
rect 38396 7274 38424 7822
rect 38384 7268 38436 7274
rect 38488 7256 38516 7822
rect 38580 7392 38608 8191
rect 38672 7392 38700 9318
rect 38764 9160 38792 10231
rect 38934 9752 38990 9761
rect 38934 9687 38990 9696
rect 38948 9586 38976 9687
rect 38936 9580 38988 9586
rect 38936 9522 38988 9528
rect 38764 9132 38976 9160
rect 38948 8974 38976 9132
rect 38936 8968 38988 8974
rect 38936 8910 38988 8916
rect 38844 8832 38896 8838
rect 38844 8774 38896 8780
rect 38750 7984 38806 7993
rect 38750 7919 38806 7928
rect 38764 7886 38792 7919
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 38580 7364 38700 7392
rect 38488 7228 38608 7256
rect 38384 7210 38436 7216
rect 38474 7168 38530 7177
rect 38474 7103 38530 7112
rect 38384 6996 38436 7002
rect 38384 6938 38436 6944
rect 38292 6860 38344 6866
rect 37832 6724 37884 6730
rect 37832 6666 37884 6672
rect 37844 5914 37872 6666
rect 37924 6656 37976 6662
rect 37924 6598 37976 6604
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37832 5568 37884 5574
rect 37752 5528 37832 5556
rect 37832 5510 37884 5516
rect 37844 4865 37872 5510
rect 37830 4856 37886 4865
rect 37936 4826 37964 6598
rect 37830 4791 37886 4800
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 37464 4208 37516 4214
rect 37464 4150 37516 4156
rect 37476 3233 37504 4150
rect 37936 4010 37964 4490
rect 37924 4004 37976 4010
rect 37924 3946 37976 3952
rect 37648 3936 37700 3942
rect 37648 3878 37700 3884
rect 37740 3936 37792 3942
rect 38028 3913 38056 6854
rect 38292 6802 38344 6808
rect 38200 6724 38252 6730
rect 38200 6666 38252 6672
rect 38212 6633 38240 6666
rect 38198 6624 38254 6633
rect 38198 6559 38254 6568
rect 38200 6452 38252 6458
rect 38200 6394 38252 6400
rect 38212 5658 38240 6394
rect 38292 6384 38344 6390
rect 38396 6372 38424 6938
rect 38488 6798 38516 7103
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38344 6344 38424 6372
rect 38292 6326 38344 6332
rect 38476 6112 38528 6118
rect 38476 6054 38528 6060
rect 38384 5772 38436 5778
rect 38384 5714 38436 5720
rect 38120 5630 38240 5658
rect 37740 3878 37792 3884
rect 38014 3904 38070 3913
rect 37556 3664 37608 3670
rect 37556 3606 37608 3612
rect 37462 3224 37518 3233
rect 37462 3159 37518 3168
rect 37292 2746 37412 2774
rect 37292 2582 37320 2746
rect 37280 2576 37332 2582
rect 37280 2518 37332 2524
rect 37280 1420 37332 1426
rect 37280 1362 37332 1368
rect 37292 800 37320 1362
rect 37568 800 37596 3606
rect 37660 2650 37688 3878
rect 37752 3534 37780 3878
rect 38014 3839 38070 3848
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 37832 2916 37884 2922
rect 37832 2858 37884 2864
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37844 800 37872 2858
rect 38120 800 38148 5630
rect 38200 5568 38252 5574
rect 38200 5510 38252 5516
rect 38212 3058 38240 5510
rect 38292 5228 38344 5234
rect 38292 5170 38344 5176
rect 38304 4690 38332 5170
rect 38396 4729 38424 5714
rect 38488 5642 38516 6054
rect 38476 5636 38528 5642
rect 38476 5578 38528 5584
rect 38580 5370 38608 7228
rect 38764 5914 38792 7822
rect 38856 7313 38884 8774
rect 38934 8664 38990 8673
rect 38934 8599 38990 8608
rect 38842 7304 38898 7313
rect 38842 7239 38898 7248
rect 38752 5908 38804 5914
rect 38752 5850 38804 5856
rect 38948 5642 38976 8599
rect 39040 6458 39068 17478
rect 39132 16658 39160 20266
rect 39224 19854 39252 20334
rect 39212 19848 39264 19854
rect 39212 19790 39264 19796
rect 39224 18766 39252 19790
rect 39396 18896 39448 18902
rect 39396 18838 39448 18844
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39212 18624 39264 18630
rect 39212 18566 39264 18572
rect 39224 17649 39252 18566
rect 39210 17640 39266 17649
rect 39210 17575 39266 17584
rect 39224 17542 39252 17575
rect 39212 17536 39264 17542
rect 39212 17478 39264 17484
rect 39120 16652 39172 16658
rect 39120 16594 39172 16600
rect 39132 16046 39160 16594
rect 39120 16040 39172 16046
rect 39120 15982 39172 15988
rect 39212 15972 39264 15978
rect 39212 15914 39264 15920
rect 39224 15502 39252 15914
rect 39212 15496 39264 15502
rect 39212 15438 39264 15444
rect 39120 15156 39172 15162
rect 39172 15116 39252 15144
rect 39120 15098 39172 15104
rect 39120 15020 39172 15026
rect 39120 14962 39172 14968
rect 39132 14929 39160 14962
rect 39118 14920 39174 14929
rect 39118 14855 39174 14864
rect 39224 14822 39252 15116
rect 39408 15094 39436 18838
rect 39396 15088 39448 15094
rect 39396 15030 39448 15036
rect 39304 14952 39356 14958
rect 39356 14912 39436 14940
rect 39304 14894 39356 14900
rect 39212 14816 39264 14822
rect 39212 14758 39264 14764
rect 39212 14476 39264 14482
rect 39212 14418 39264 14424
rect 39120 12708 39172 12714
rect 39120 12650 39172 12656
rect 39132 12442 39160 12650
rect 39120 12436 39172 12442
rect 39120 12378 39172 12384
rect 39224 10198 39252 14418
rect 39408 14278 39436 14912
rect 39396 14272 39448 14278
rect 39394 14240 39396 14249
rect 39448 14240 39450 14249
rect 39394 14175 39450 14184
rect 39396 11348 39448 11354
rect 39396 11290 39448 11296
rect 39212 10192 39264 10198
rect 39212 10134 39264 10140
rect 39120 9988 39172 9994
rect 39120 9930 39172 9936
rect 39212 9988 39264 9994
rect 39212 9930 39264 9936
rect 39132 9178 39160 9930
rect 39120 9172 39172 9178
rect 39120 9114 39172 9120
rect 39120 8900 39172 8906
rect 39120 8842 39172 8848
rect 39132 8294 39160 8842
rect 39120 8288 39172 8294
rect 39120 8230 39172 8236
rect 39120 7880 39172 7886
rect 39118 7848 39120 7857
rect 39172 7848 39174 7857
rect 39118 7783 39174 7792
rect 39120 7472 39172 7478
rect 39224 7449 39252 9930
rect 39304 9648 39356 9654
rect 39304 9590 39356 9596
rect 39120 7414 39172 7420
rect 39210 7440 39266 7449
rect 39132 7313 39160 7414
rect 39210 7375 39266 7384
rect 39118 7304 39174 7313
rect 39118 7239 39174 7248
rect 39212 7200 39264 7206
rect 39212 7142 39264 7148
rect 39028 6452 39080 6458
rect 39028 6394 39080 6400
rect 39120 5908 39172 5914
rect 39120 5850 39172 5856
rect 38936 5636 38988 5642
rect 38856 5596 38936 5624
rect 38476 5364 38528 5370
rect 38476 5306 38528 5312
rect 38568 5364 38620 5370
rect 38568 5306 38620 5312
rect 38488 5216 38516 5306
rect 38660 5296 38712 5302
rect 38660 5238 38712 5244
rect 38568 5228 38620 5234
rect 38488 5188 38568 5216
rect 38568 5170 38620 5176
rect 38476 5024 38528 5030
rect 38476 4966 38528 4972
rect 38382 4720 38438 4729
rect 38292 4684 38344 4690
rect 38382 4655 38438 4664
rect 38292 4626 38344 4632
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38292 3392 38344 3398
rect 38292 3334 38344 3340
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 38304 2990 38332 3334
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 38396 800 38424 3402
rect 38488 2582 38516 4966
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 38580 3466 38608 4558
rect 38672 4214 38700 5238
rect 38752 5092 38804 5098
rect 38752 5034 38804 5040
rect 38660 4208 38712 4214
rect 38660 4150 38712 4156
rect 38672 3602 38700 4150
rect 38764 4078 38792 5034
rect 38752 4072 38804 4078
rect 38752 4014 38804 4020
rect 38856 3942 38884 5596
rect 38936 5578 38988 5584
rect 38936 4548 38988 4554
rect 38936 4490 38988 4496
rect 38948 4146 38976 4490
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 39026 4040 39082 4049
rect 39132 4010 39160 5850
rect 39224 5030 39252 7142
rect 39212 5024 39264 5030
rect 39212 4966 39264 4972
rect 39316 4758 39344 9590
rect 39408 8634 39436 11290
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 39408 7886 39436 8570
rect 39396 7880 39448 7886
rect 39396 7822 39448 7828
rect 39396 5092 39448 5098
rect 39396 5034 39448 5040
rect 39304 4752 39356 4758
rect 39304 4694 39356 4700
rect 39408 4282 39436 5034
rect 39396 4276 39448 4282
rect 39396 4218 39448 4224
rect 39304 4140 39356 4146
rect 39304 4082 39356 4088
rect 39026 3975 39082 3984
rect 39120 4004 39172 4010
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 38844 3936 38896 3942
rect 38844 3878 38896 3884
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38672 3466 38700 3538
rect 38568 3460 38620 3466
rect 38568 3402 38620 3408
rect 38660 3460 38712 3466
rect 38660 3402 38712 3408
rect 38476 2576 38528 2582
rect 38476 2518 38528 2524
rect 38568 2576 38620 2582
rect 38568 2518 38620 2524
rect 38580 1426 38608 2518
rect 38764 2514 38792 3878
rect 38856 3058 38884 3878
rect 39040 3738 39068 3975
rect 39120 3946 39172 3952
rect 39028 3732 39080 3738
rect 39028 3674 39080 3680
rect 39316 3505 39344 4082
rect 39302 3496 39358 3505
rect 38936 3460 38988 3466
rect 39302 3431 39358 3440
rect 38936 3402 38988 3408
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38948 2938 38976 3402
rect 39500 3194 39528 28426
rect 39592 15094 39620 61202
rect 39960 61180 39988 63294
rect 40590 63294 41000 63322
rect 40590 63200 40646 63294
rect 40316 61668 40368 61674
rect 40316 61610 40368 61616
rect 40408 61668 40460 61674
rect 40408 61610 40460 61616
rect 40328 61334 40356 61610
rect 40420 61402 40448 61610
rect 40684 61600 40736 61606
rect 40684 61542 40736 61548
rect 40696 61402 40724 61542
rect 40408 61396 40460 61402
rect 40408 61338 40460 61344
rect 40684 61396 40736 61402
rect 40684 61338 40736 61344
rect 40316 61328 40368 61334
rect 40316 61270 40368 61276
rect 40972 61198 41000 63294
rect 41326 63200 41382 64000
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63200 43590 64000
rect 44270 63322 44326 64000
rect 45006 63322 45062 64000
rect 45742 63322 45798 64000
rect 46478 63322 46534 64000
rect 44270 63294 44588 63322
rect 44270 63200 44326 63294
rect 41236 61736 41288 61742
rect 41236 61678 41288 61684
rect 41144 61260 41196 61266
rect 41144 61202 41196 61208
rect 40132 61192 40184 61198
rect 39960 61152 40132 61180
rect 40132 61134 40184 61140
rect 40960 61192 41012 61198
rect 40960 61134 41012 61140
rect 39764 61124 39816 61130
rect 39764 61066 39816 61072
rect 39776 59673 39804 61066
rect 40316 61056 40368 61062
rect 40316 60998 40368 61004
rect 39762 59664 39818 59673
rect 39762 59599 39818 59608
rect 39948 56296 40000 56302
rect 39948 56238 40000 56244
rect 39960 55350 39988 56238
rect 39948 55344 40000 55350
rect 39948 55286 40000 55292
rect 40040 55208 40092 55214
rect 40040 55150 40092 55156
rect 39672 53100 39724 53106
rect 39672 53042 39724 53048
rect 39684 15450 39712 53042
rect 39856 45552 39908 45558
rect 39856 45494 39908 45500
rect 39764 20324 39816 20330
rect 39764 20266 39816 20272
rect 39776 19922 39804 20266
rect 39764 19916 39816 19922
rect 39764 19858 39816 19864
rect 39868 19009 39896 45494
rect 39948 25288 40000 25294
rect 39948 25230 40000 25236
rect 39854 19000 39910 19009
rect 39854 18935 39910 18944
rect 39960 18850 39988 25230
rect 40052 21418 40080 55150
rect 40328 35086 40356 60998
rect 41052 59968 41104 59974
rect 41052 59910 41104 59916
rect 40776 59016 40828 59022
rect 40776 58958 40828 58964
rect 40788 58546 40816 58958
rect 40868 58880 40920 58886
rect 40868 58822 40920 58828
rect 40776 58540 40828 58546
rect 40776 58482 40828 58488
rect 40408 58336 40460 58342
rect 40408 58278 40460 58284
rect 40420 58041 40448 58278
rect 40406 58032 40462 58041
rect 40406 57967 40462 57976
rect 40880 53718 40908 58822
rect 40868 53712 40920 53718
rect 40868 53654 40920 53660
rect 40408 53440 40460 53446
rect 40408 53382 40460 53388
rect 40316 35080 40368 35086
rect 40316 35022 40368 35028
rect 40224 35012 40276 35018
rect 40224 34954 40276 34960
rect 40236 34678 40264 34954
rect 40224 34672 40276 34678
rect 40224 34614 40276 34620
rect 40420 22094 40448 53382
rect 41064 40730 41092 59910
rect 41156 58546 41184 61202
rect 41248 60738 41276 61678
rect 41340 60874 41368 63200
rect 42076 61198 42104 63200
rect 42708 61668 42760 61674
rect 42708 61610 42760 61616
rect 42064 61192 42116 61198
rect 42064 61134 42116 61140
rect 41696 61056 41748 61062
rect 41696 60998 41748 61004
rect 41340 60846 41460 60874
rect 41432 60790 41460 60846
rect 41420 60784 41472 60790
rect 41248 60706 41368 60738
rect 41420 60726 41472 60732
rect 41604 60716 41656 60722
rect 41248 59022 41276 60706
rect 41604 60658 41656 60664
rect 41616 60110 41644 60658
rect 41604 60104 41656 60110
rect 41604 60046 41656 60052
rect 41236 59016 41288 59022
rect 41236 58958 41288 58964
rect 41420 59016 41472 59022
rect 41420 58958 41472 58964
rect 41432 58546 41460 58958
rect 41144 58540 41196 58546
rect 41144 58482 41196 58488
rect 41420 58540 41472 58546
rect 41420 58482 41472 58488
rect 41432 56506 41460 58482
rect 41420 56500 41472 56506
rect 41420 56442 41472 56448
rect 41432 56302 41460 56442
rect 41420 56296 41472 56302
rect 41420 56238 41472 56244
rect 41432 55350 41460 56238
rect 41420 55344 41472 55350
rect 41420 55286 41472 55292
rect 41432 53582 41460 55286
rect 41420 53576 41472 53582
rect 41420 53518 41472 53524
rect 41052 40724 41104 40730
rect 41052 40666 41104 40672
rect 40776 36236 40828 36242
rect 40776 36178 40828 36184
rect 40684 36168 40736 36174
rect 40684 36110 40736 36116
rect 40696 35630 40724 36110
rect 40684 35624 40736 35630
rect 40684 35566 40736 35572
rect 40696 35086 40724 35566
rect 40684 35080 40736 35086
rect 40684 35022 40736 35028
rect 40788 24342 40816 36178
rect 41708 36106 41736 60998
rect 41972 60512 42024 60518
rect 41972 60454 42024 60460
rect 41880 60172 41932 60178
rect 41880 60114 41932 60120
rect 41788 60104 41840 60110
rect 41788 60046 41840 60052
rect 41800 49162 41828 60046
rect 41892 59022 41920 60114
rect 41984 60110 42012 60454
rect 41972 60104 42024 60110
rect 41972 60046 42024 60052
rect 42616 60036 42668 60042
rect 42616 59978 42668 59984
rect 42628 59401 42656 59978
rect 42720 59650 42748 61610
rect 42812 61198 42840 63200
rect 42800 61192 42852 61198
rect 43548 61180 43576 63200
rect 44560 61198 44588 63294
rect 45006 63294 45508 63322
rect 45006 63200 45062 63294
rect 45480 61282 45508 63294
rect 45742 63294 46152 63322
rect 45742 63200 45798 63294
rect 45480 61254 45600 61282
rect 45572 61198 45600 61254
rect 46124 61198 46152 63294
rect 46478 63294 46704 63322
rect 46478 63200 46534 63294
rect 43628 61192 43680 61198
rect 43548 61152 43628 61180
rect 42800 61134 42852 61140
rect 43628 61134 43680 61140
rect 44548 61192 44600 61198
rect 44548 61134 44600 61140
rect 45560 61192 45612 61198
rect 45560 61134 45612 61140
rect 46112 61192 46164 61198
rect 46112 61134 46164 61140
rect 42892 61124 42944 61130
rect 42892 61066 42944 61072
rect 42720 59622 42840 59650
rect 42812 59566 42840 59622
rect 42708 59560 42760 59566
rect 42708 59502 42760 59508
rect 42800 59560 42852 59566
rect 42800 59502 42852 59508
rect 42614 59392 42670 59401
rect 42614 59327 42670 59336
rect 41880 59016 41932 59022
rect 41880 58958 41932 58964
rect 42720 57361 42748 59502
rect 42706 57352 42762 57361
rect 42706 57287 42762 57296
rect 42248 56160 42300 56166
rect 42248 56102 42300 56108
rect 41880 53712 41932 53718
rect 41880 53654 41932 53660
rect 41788 49156 41840 49162
rect 41788 49098 41840 49104
rect 41696 36100 41748 36106
rect 41696 36042 41748 36048
rect 41892 35894 41920 53654
rect 41892 35866 42012 35894
rect 41604 32564 41656 32570
rect 41604 32506 41656 32512
rect 40960 31136 41012 31142
rect 40960 31078 41012 31084
rect 40776 24336 40828 24342
rect 40776 24278 40828 24284
rect 40420 22066 40540 22094
rect 40040 21412 40092 21418
rect 40040 21354 40092 21360
rect 40224 20052 40276 20058
rect 40224 19994 40276 20000
rect 40132 19168 40184 19174
rect 40132 19110 40184 19116
rect 40144 18902 40172 19110
rect 39868 18822 39988 18850
rect 40132 18896 40184 18902
rect 40132 18838 40184 18844
rect 39868 17338 39896 18822
rect 40144 18222 40172 18838
rect 40132 18216 40184 18222
rect 40132 18158 40184 18164
rect 39856 17332 39908 17338
rect 39856 17274 39908 17280
rect 39764 16516 39816 16522
rect 39764 16458 39816 16464
rect 39776 16114 39804 16458
rect 39764 16108 39816 16114
rect 39764 16050 39816 16056
rect 39868 15502 39896 17274
rect 40236 17202 40264 19994
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 40328 18290 40356 19790
rect 40316 18284 40368 18290
rect 40316 18226 40368 18232
rect 40224 17196 40276 17202
rect 40224 17138 40276 17144
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 39960 15638 39988 17070
rect 40236 16726 40264 17138
rect 40328 17082 40356 18226
rect 40328 17054 40448 17082
rect 40420 16998 40448 17054
rect 40316 16992 40368 16998
rect 40316 16934 40368 16940
rect 40408 16992 40460 16998
rect 40408 16934 40460 16940
rect 40328 16726 40356 16934
rect 40224 16720 40276 16726
rect 40224 16662 40276 16668
rect 40316 16720 40368 16726
rect 40316 16662 40368 16668
rect 40408 16584 40460 16590
rect 40408 16526 40460 16532
rect 40132 16448 40184 16454
rect 40132 16390 40184 16396
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40052 15978 40080 16186
rect 40040 15972 40092 15978
rect 40040 15914 40092 15920
rect 39948 15632 40000 15638
rect 39948 15574 40000 15580
rect 39856 15496 39908 15502
rect 39684 15422 39804 15450
rect 39856 15438 39908 15444
rect 40144 15434 40172 16390
rect 40316 16244 40368 16250
rect 40316 16186 40368 16192
rect 40224 16108 40276 16114
rect 40328 16096 40356 16186
rect 40420 16114 40448 16526
rect 40276 16068 40356 16096
rect 40224 16050 40276 16056
rect 39580 15088 39632 15094
rect 39580 15030 39632 15036
rect 39672 14272 39724 14278
rect 39672 14214 39724 14220
rect 39684 14006 39712 14214
rect 39672 14000 39724 14006
rect 39672 13942 39724 13948
rect 39776 13258 39804 15422
rect 40132 15428 40184 15434
rect 40132 15370 40184 15376
rect 40328 15366 40356 16068
rect 40408 16108 40460 16114
rect 40408 16050 40460 16056
rect 40316 15360 40368 15366
rect 40316 15302 40368 15308
rect 40328 15201 40356 15302
rect 40314 15192 40370 15201
rect 40314 15127 40370 15136
rect 39856 15088 39908 15094
rect 39856 15030 39908 15036
rect 39764 13252 39816 13258
rect 39764 13194 39816 13200
rect 39672 12844 39724 12850
rect 39672 12786 39724 12792
rect 39580 12708 39632 12714
rect 39580 12650 39632 12656
rect 39592 12102 39620 12650
rect 39580 12096 39632 12102
rect 39580 12038 39632 12044
rect 39592 11762 39620 12038
rect 39684 11898 39712 12786
rect 39764 12776 39816 12782
rect 39764 12718 39816 12724
rect 39776 12238 39804 12718
rect 39764 12232 39816 12238
rect 39764 12174 39816 12180
rect 39672 11892 39724 11898
rect 39672 11834 39724 11840
rect 39580 11756 39632 11762
rect 39580 11698 39632 11704
rect 39592 10674 39620 11698
rect 39580 10668 39632 10674
rect 39580 10610 39632 10616
rect 39592 9761 39620 10610
rect 39578 9752 39634 9761
rect 39578 9687 39634 9696
rect 39592 9217 39620 9687
rect 39868 9654 39896 15030
rect 40316 14816 40368 14822
rect 40316 14758 40368 14764
rect 40130 14648 40186 14657
rect 40328 14634 40356 14758
rect 40130 14583 40186 14592
rect 40236 14606 40356 14634
rect 40144 13394 40172 14583
rect 40236 14414 40264 14606
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 40408 14068 40460 14074
rect 40408 14010 40460 14016
rect 40420 13870 40448 14010
rect 40408 13864 40460 13870
rect 40408 13806 40460 13812
rect 40408 13728 40460 13734
rect 40314 13696 40370 13705
rect 40408 13670 40460 13676
rect 40314 13631 40370 13640
rect 40328 13462 40356 13631
rect 40420 13462 40448 13670
rect 40316 13456 40368 13462
rect 40316 13398 40368 13404
rect 40408 13456 40460 13462
rect 40408 13398 40460 13404
rect 40132 13388 40184 13394
rect 40132 13330 40184 13336
rect 40040 13320 40092 13326
rect 40512 13308 40540 22066
rect 40868 19848 40920 19854
rect 40868 19790 40920 19796
rect 40776 19712 40828 19718
rect 40776 19654 40828 19660
rect 40684 19304 40736 19310
rect 40682 19272 40684 19281
rect 40736 19272 40738 19281
rect 40592 19236 40644 19242
rect 40682 19207 40738 19216
rect 40592 19178 40644 19184
rect 40604 19145 40632 19178
rect 40590 19136 40646 19145
rect 40590 19071 40646 19080
rect 40788 18766 40816 19654
rect 40880 19514 40908 19790
rect 40868 19508 40920 19514
rect 40868 19450 40920 19456
rect 40592 18760 40644 18766
rect 40592 18702 40644 18708
rect 40776 18760 40828 18766
rect 40776 18702 40828 18708
rect 40604 17678 40632 18702
rect 40684 18692 40736 18698
rect 40684 18634 40736 18640
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40592 17536 40644 17542
rect 40592 17478 40644 17484
rect 40604 17338 40632 17478
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 40604 16454 40632 17274
rect 40592 16448 40644 16454
rect 40592 16390 40644 16396
rect 40604 16182 40632 16390
rect 40592 16176 40644 16182
rect 40592 16118 40644 16124
rect 40592 15904 40644 15910
rect 40592 15846 40644 15852
rect 40604 15473 40632 15846
rect 40590 15464 40646 15473
rect 40590 15399 40646 15408
rect 40592 15360 40644 15366
rect 40592 15302 40644 15308
rect 40604 14822 40632 15302
rect 40592 14816 40644 14822
rect 40592 14758 40644 14764
rect 40592 14340 40644 14346
rect 40592 14282 40644 14288
rect 40604 14113 40632 14282
rect 40590 14104 40646 14113
rect 40590 14039 40646 14048
rect 40696 13546 40724 18634
rect 40868 18216 40920 18222
rect 40868 18158 40920 18164
rect 40776 14816 40828 14822
rect 40776 14758 40828 14764
rect 40788 14482 40816 14758
rect 40776 14476 40828 14482
rect 40776 14418 40828 14424
rect 40788 14074 40816 14418
rect 40776 14068 40828 14074
rect 40776 14010 40828 14016
rect 40776 13864 40828 13870
rect 40776 13806 40828 13812
rect 40040 13262 40092 13268
rect 40328 13280 40540 13308
rect 40604 13518 40724 13546
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39960 12850 39988 13126
rect 39948 12844 40000 12850
rect 39948 12786 40000 12792
rect 39946 12744 40002 12753
rect 39946 12679 40002 12688
rect 39960 12646 39988 12679
rect 39948 12640 40000 12646
rect 39948 12582 40000 12588
rect 40052 12481 40080 13262
rect 40038 12472 40094 12481
rect 40038 12407 40094 12416
rect 40132 12096 40184 12102
rect 40130 12064 40132 12073
rect 40184 12064 40186 12073
rect 40130 11999 40186 12008
rect 40328 11762 40356 13280
rect 40604 13002 40632 13518
rect 40684 13456 40736 13462
rect 40684 13398 40736 13404
rect 40512 12974 40632 13002
rect 40512 12753 40540 12974
rect 40696 12850 40724 13398
rect 40788 13326 40816 13806
rect 40776 13320 40828 13326
rect 40776 13262 40828 13268
rect 40788 12850 40816 13262
rect 40684 12844 40736 12850
rect 40684 12786 40736 12792
rect 40776 12844 40828 12850
rect 40776 12786 40828 12792
rect 40498 12744 40554 12753
rect 40498 12679 40554 12688
rect 40500 12640 40552 12646
rect 40500 12582 40552 12588
rect 40512 11762 40540 12582
rect 40788 11914 40816 12786
rect 40880 12102 40908 18158
rect 40972 12918 41000 31078
rect 41144 23316 41196 23322
rect 41144 23258 41196 23264
rect 41156 20058 41184 23258
rect 41328 21956 41380 21962
rect 41328 21898 41380 21904
rect 41144 20052 41196 20058
rect 41144 19994 41196 20000
rect 41236 19508 41288 19514
rect 41064 19468 41236 19496
rect 41064 19310 41092 19468
rect 41236 19450 41288 19456
rect 41052 19304 41104 19310
rect 41236 19304 41288 19310
rect 41052 19246 41104 19252
rect 41234 19272 41236 19281
rect 41288 19272 41290 19281
rect 41064 19174 41092 19246
rect 41234 19207 41290 19216
rect 41052 19168 41104 19174
rect 41052 19110 41104 19116
rect 41236 19168 41288 19174
rect 41236 19110 41288 19116
rect 41248 18222 41276 19110
rect 41236 18216 41288 18222
rect 41236 18158 41288 18164
rect 41144 17876 41196 17882
rect 41144 17818 41196 17824
rect 41052 17808 41104 17814
rect 41052 17750 41104 17756
rect 41064 17066 41092 17750
rect 41156 17338 41184 17818
rect 41144 17332 41196 17338
rect 41144 17274 41196 17280
rect 41052 17060 41104 17066
rect 41052 17002 41104 17008
rect 41052 16652 41104 16658
rect 41248 16640 41276 18158
rect 41104 16612 41276 16640
rect 41052 16594 41104 16600
rect 41064 16250 41092 16594
rect 41340 16454 41368 21898
rect 41420 19916 41472 19922
rect 41420 19858 41472 19864
rect 41432 19378 41460 19858
rect 41420 19372 41472 19378
rect 41420 19314 41472 19320
rect 41420 17128 41472 17134
rect 41420 17070 41472 17076
rect 41432 16658 41460 17070
rect 41512 16992 41564 16998
rect 41512 16934 41564 16940
rect 41420 16652 41472 16658
rect 41420 16594 41472 16600
rect 41524 16522 41552 16934
rect 41512 16516 41564 16522
rect 41512 16458 41564 16464
rect 41144 16448 41196 16454
rect 41144 16390 41196 16396
rect 41328 16448 41380 16454
rect 41328 16390 41380 16396
rect 41052 16244 41104 16250
rect 41052 16186 41104 16192
rect 41052 15564 41104 15570
rect 41052 15506 41104 15512
rect 41064 14657 41092 15506
rect 41050 14648 41106 14657
rect 41050 14583 41106 14592
rect 41052 14340 41104 14346
rect 41052 14282 41104 14288
rect 41064 13938 41092 14282
rect 41052 13932 41104 13938
rect 41052 13874 41104 13880
rect 41052 13796 41104 13802
rect 41052 13738 41104 13744
rect 41064 13530 41092 13738
rect 41156 13569 41184 16390
rect 41512 16176 41564 16182
rect 41512 16118 41564 16124
rect 41328 15904 41380 15910
rect 41328 15846 41380 15852
rect 41340 15094 41368 15846
rect 41524 15502 41552 16118
rect 41512 15496 41564 15502
rect 41512 15438 41564 15444
rect 41328 15088 41380 15094
rect 41328 15030 41380 15036
rect 41418 14920 41474 14929
rect 41418 14855 41474 14864
rect 41432 14550 41460 14855
rect 41328 14544 41380 14550
rect 41328 14486 41380 14492
rect 41420 14544 41472 14550
rect 41420 14486 41472 14492
rect 41340 14414 41368 14486
rect 41524 14482 41552 15438
rect 41512 14476 41564 14482
rect 41512 14418 41564 14424
rect 41236 14408 41288 14414
rect 41236 14350 41288 14356
rect 41328 14408 41380 14414
rect 41328 14350 41380 14356
rect 41248 14006 41276 14350
rect 41616 14006 41644 32506
rect 41696 19508 41748 19514
rect 41696 19450 41748 19456
rect 41708 18290 41736 19450
rect 41880 19236 41932 19242
rect 41880 19178 41932 19184
rect 41892 18902 41920 19178
rect 41880 18896 41932 18902
rect 41880 18838 41932 18844
rect 41696 18284 41748 18290
rect 41696 18226 41748 18232
rect 41788 17604 41840 17610
rect 41788 17546 41840 17552
rect 41696 17536 41748 17542
rect 41696 17478 41748 17484
rect 41708 16250 41736 17478
rect 41800 16726 41828 17546
rect 41788 16720 41840 16726
rect 41788 16662 41840 16668
rect 41696 16244 41748 16250
rect 41696 16186 41748 16192
rect 41788 16040 41840 16046
rect 41788 15982 41840 15988
rect 41800 15706 41828 15982
rect 41788 15700 41840 15706
rect 41788 15642 41840 15648
rect 41800 15162 41828 15642
rect 41788 15156 41840 15162
rect 41788 15098 41840 15104
rect 41880 14408 41932 14414
rect 41880 14350 41932 14356
rect 41892 14074 41920 14350
rect 41880 14068 41932 14074
rect 41880 14010 41932 14016
rect 41236 14000 41288 14006
rect 41236 13942 41288 13948
rect 41604 14000 41656 14006
rect 41984 13954 42012 35866
rect 42064 21412 42116 21418
rect 42064 21354 42116 21360
rect 41604 13942 41656 13948
rect 41708 13926 42012 13954
rect 41328 13796 41380 13802
rect 41328 13738 41380 13744
rect 41142 13560 41198 13569
rect 41052 13524 41104 13530
rect 41142 13495 41198 13504
rect 41052 13466 41104 13472
rect 41052 13320 41104 13326
rect 41052 13262 41104 13268
rect 41144 13320 41196 13326
rect 41144 13262 41196 13268
rect 40960 12912 41012 12918
rect 40960 12854 41012 12860
rect 41064 12170 41092 13262
rect 41052 12164 41104 12170
rect 41052 12106 41104 12112
rect 40868 12096 40920 12102
rect 40868 12038 40920 12044
rect 40788 11886 41000 11914
rect 40684 11824 40736 11830
rect 40684 11766 40736 11772
rect 40132 11756 40184 11762
rect 40316 11756 40368 11762
rect 40184 11716 40264 11744
rect 40132 11698 40184 11704
rect 39948 10056 40000 10062
rect 39948 9998 40000 10004
rect 40040 10056 40092 10062
rect 40040 9998 40092 10004
rect 39856 9648 39908 9654
rect 39762 9616 39818 9625
rect 39856 9590 39908 9596
rect 39762 9551 39764 9560
rect 39816 9551 39818 9560
rect 39764 9522 39816 9528
rect 39856 9512 39908 9518
rect 39856 9454 39908 9460
rect 39672 9444 39724 9450
rect 39672 9386 39724 9392
rect 39684 9353 39712 9386
rect 39670 9344 39726 9353
rect 39670 9279 39726 9288
rect 39578 9208 39634 9217
rect 39578 9143 39634 9152
rect 39868 9058 39896 9454
rect 39592 9042 39896 9058
rect 39580 9036 39896 9042
rect 39632 9030 39896 9036
rect 39580 8978 39632 8984
rect 39764 8968 39816 8974
rect 39764 8910 39816 8916
rect 39580 8900 39632 8906
rect 39580 8842 39632 8848
rect 39592 8634 39620 8842
rect 39580 8628 39632 8634
rect 39580 8570 39632 8576
rect 39672 8560 39724 8566
rect 39670 8528 39672 8537
rect 39724 8528 39726 8537
rect 39670 8463 39726 8472
rect 39776 8344 39804 8910
rect 39856 8900 39908 8906
rect 39856 8842 39908 8848
rect 39684 8316 39804 8344
rect 39684 6361 39712 8316
rect 39762 8256 39818 8265
rect 39762 8191 39818 8200
rect 39776 7818 39804 8191
rect 39868 7954 39896 8842
rect 39856 7948 39908 7954
rect 39856 7890 39908 7896
rect 39764 7812 39816 7818
rect 39764 7754 39816 7760
rect 39670 6352 39726 6361
rect 39670 6287 39726 6296
rect 39580 5228 39632 5234
rect 39580 5170 39632 5176
rect 39592 3398 39620 5170
rect 39960 4690 39988 9998
rect 40052 9450 40080 9998
rect 40236 9908 40264 11716
rect 40316 11698 40368 11704
rect 40500 11756 40552 11762
rect 40500 11698 40552 11704
rect 40592 11688 40644 11694
rect 40512 11636 40592 11642
rect 40512 11630 40644 11636
rect 40512 11614 40632 11630
rect 40512 10470 40540 11614
rect 40696 11529 40724 11766
rect 40776 11688 40828 11694
rect 40776 11630 40828 11636
rect 40682 11520 40738 11529
rect 40682 11455 40738 11464
rect 40684 11280 40736 11286
rect 40684 11222 40736 11228
rect 40696 10996 40724 11222
rect 40788 11150 40816 11630
rect 40866 11384 40922 11393
rect 40866 11319 40922 11328
rect 40776 11144 40828 11150
rect 40776 11086 40828 11092
rect 40696 10968 40816 10996
rect 40592 10668 40644 10674
rect 40592 10610 40644 10616
rect 40316 10464 40368 10470
rect 40316 10406 40368 10412
rect 40500 10464 40552 10470
rect 40500 10406 40552 10412
rect 40328 10033 40356 10406
rect 40408 10192 40460 10198
rect 40408 10134 40460 10140
rect 40314 10024 40370 10033
rect 40314 9959 40370 9968
rect 40236 9880 40356 9908
rect 40222 9752 40278 9761
rect 40222 9687 40278 9696
rect 40040 9444 40092 9450
rect 40040 9386 40092 9392
rect 40052 8498 40080 9386
rect 40130 9344 40186 9353
rect 40130 9279 40186 9288
rect 40040 8492 40092 8498
rect 40040 8434 40092 8440
rect 40040 8356 40092 8362
rect 40040 8298 40092 8304
rect 40052 7993 40080 8298
rect 40144 8294 40172 9279
rect 40132 8288 40184 8294
rect 40132 8230 40184 8236
rect 40038 7984 40094 7993
rect 40038 7919 40094 7928
rect 40132 7880 40184 7886
rect 40132 7822 40184 7828
rect 40144 7410 40172 7822
rect 40132 7404 40184 7410
rect 40132 7346 40184 7352
rect 40040 6792 40092 6798
rect 40040 6734 40092 6740
rect 40052 6458 40080 6734
rect 40040 6452 40092 6458
rect 40040 6394 40092 6400
rect 40132 5160 40184 5166
rect 40132 5102 40184 5108
rect 39948 4684 40000 4690
rect 39948 4626 40000 4632
rect 40040 4684 40092 4690
rect 40040 4626 40092 4632
rect 39948 4140 40000 4146
rect 39948 4082 40000 4088
rect 39960 3942 39988 4082
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 39580 3392 39632 3398
rect 39580 3334 39632 3340
rect 39488 3188 39540 3194
rect 39488 3130 39540 3136
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 38856 2910 38976 2938
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 38672 2038 38700 2314
rect 38660 2032 38712 2038
rect 38660 1974 38712 1980
rect 38568 1420 38620 1426
rect 38568 1362 38620 1368
rect 38856 1170 38884 2910
rect 39132 2774 39160 2994
rect 38672 1142 38884 1170
rect 38948 2746 39160 2774
rect 38672 800 38700 1142
rect 38948 800 38976 2746
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 39224 800 39252 2314
rect 39488 1692 39540 1698
rect 39488 1634 39540 1640
rect 39500 800 39528 1634
rect 39776 800 39804 2994
rect 40052 800 40080 4626
rect 40144 3466 40172 5102
rect 40236 4826 40264 9687
rect 40328 9518 40356 9880
rect 40316 9512 40368 9518
rect 40316 9454 40368 9460
rect 40328 8498 40356 9454
rect 40420 8974 40448 10134
rect 40500 9580 40552 9586
rect 40500 9522 40552 9528
rect 40408 8968 40460 8974
rect 40408 8910 40460 8916
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 40420 7274 40448 8910
rect 40512 8537 40540 9522
rect 40604 9042 40632 10610
rect 40788 10554 40816 10968
rect 40880 10674 40908 11319
rect 40972 10810 41000 11886
rect 41156 11880 41184 13262
rect 41340 12850 41368 13738
rect 41512 13728 41564 13734
rect 41432 13688 41512 13716
rect 41432 13462 41460 13688
rect 41512 13670 41564 13676
rect 41602 13696 41658 13705
rect 41602 13631 41658 13640
rect 41420 13456 41472 13462
rect 41420 13398 41472 13404
rect 41512 13456 41564 13462
rect 41512 13398 41564 13404
rect 41420 13320 41472 13326
rect 41524 13308 41552 13398
rect 41472 13280 41552 13308
rect 41420 13262 41472 13268
rect 41420 13184 41472 13190
rect 41420 13126 41472 13132
rect 41328 12844 41380 12850
rect 41328 12786 41380 12792
rect 41234 12608 41290 12617
rect 41234 12543 41290 12552
rect 41064 11852 41184 11880
rect 40960 10804 41012 10810
rect 40960 10746 41012 10752
rect 40868 10668 40920 10674
rect 40868 10610 40920 10616
rect 40960 10668 41012 10674
rect 40960 10610 41012 10616
rect 40788 10526 40908 10554
rect 40776 10464 40828 10470
rect 40682 10432 40738 10441
rect 40776 10406 40828 10412
rect 40682 10367 40738 10376
rect 40696 10062 40724 10367
rect 40788 10062 40816 10406
rect 40684 10056 40736 10062
rect 40684 9998 40736 10004
rect 40776 10056 40828 10062
rect 40776 9998 40828 10004
rect 40788 9586 40816 9998
rect 40776 9580 40828 9586
rect 40776 9522 40828 9528
rect 40776 9376 40828 9382
rect 40776 9318 40828 9324
rect 40592 9036 40644 9042
rect 40592 8978 40644 8984
rect 40684 8968 40736 8974
rect 40684 8910 40736 8916
rect 40696 8838 40724 8910
rect 40684 8832 40736 8838
rect 40684 8774 40736 8780
rect 40592 8628 40644 8634
rect 40592 8570 40644 8576
rect 40498 8528 40554 8537
rect 40554 8492 40557 8498
rect 40498 8463 40505 8472
rect 40505 8434 40557 8440
rect 40408 7268 40460 7274
rect 40408 7210 40460 7216
rect 40604 6798 40632 8570
rect 40682 8392 40738 8401
rect 40682 8327 40738 8336
rect 40592 6792 40644 6798
rect 40592 6734 40644 6740
rect 40408 5704 40460 5710
rect 40408 5646 40460 5652
rect 40316 5296 40368 5302
rect 40316 5238 40368 5244
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 40132 3460 40184 3466
rect 40132 3402 40184 3408
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 40144 2514 40172 2790
rect 40222 2680 40278 2689
rect 40222 2615 40224 2624
rect 40276 2615 40278 2624
rect 40224 2586 40276 2592
rect 40132 2508 40184 2514
rect 40132 2450 40184 2456
rect 40328 800 40356 5238
rect 40420 4078 40448 5646
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40408 4072 40460 4078
rect 40408 4014 40460 4020
rect 40512 3670 40540 5170
rect 40592 5024 40644 5030
rect 40592 4966 40644 4972
rect 40604 4758 40632 4966
rect 40592 4752 40644 4758
rect 40592 4694 40644 4700
rect 40590 4040 40646 4049
rect 40590 3975 40646 3984
rect 40500 3664 40552 3670
rect 40500 3606 40552 3612
rect 40604 3194 40632 3975
rect 40696 3670 40724 8327
rect 40788 8090 40816 9318
rect 40880 8809 40908 10526
rect 40972 9722 41000 10610
rect 41064 9994 41092 11852
rect 41144 11756 41196 11762
rect 41144 11698 41196 11704
rect 41156 11218 41184 11698
rect 41144 11212 41196 11218
rect 41144 11154 41196 11160
rect 41144 10804 41196 10810
rect 41144 10746 41196 10752
rect 41052 9988 41104 9994
rect 41052 9930 41104 9936
rect 40960 9716 41012 9722
rect 40960 9658 41012 9664
rect 40960 9376 41012 9382
rect 40960 9318 41012 9324
rect 40866 8800 40922 8809
rect 40866 8735 40922 8744
rect 40868 8560 40920 8566
rect 40868 8502 40920 8508
rect 40880 8265 40908 8502
rect 40866 8256 40922 8265
rect 40866 8191 40922 8200
rect 40776 8084 40828 8090
rect 40776 8026 40828 8032
rect 40868 6792 40920 6798
rect 40868 6734 40920 6740
rect 40880 5710 40908 6734
rect 40868 5704 40920 5710
rect 40868 5646 40920 5652
rect 40776 5364 40828 5370
rect 40776 5306 40828 5312
rect 40684 3664 40736 3670
rect 40684 3606 40736 3612
rect 40592 3188 40644 3194
rect 40592 3130 40644 3136
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 40788 1494 40816 5306
rect 40880 4486 40908 5646
rect 40868 4480 40920 4486
rect 40868 4422 40920 4428
rect 40868 2848 40920 2854
rect 40868 2790 40920 2796
rect 40776 1488 40828 1494
rect 40776 1430 40828 1436
rect 40880 800 40908 2790
rect 40972 1358 41000 9318
rect 41156 8974 41184 10746
rect 41248 9382 41276 12543
rect 41340 10470 41368 12786
rect 41432 12782 41460 13126
rect 41420 12776 41472 12782
rect 41420 12718 41472 12724
rect 41512 12708 41564 12714
rect 41512 12650 41564 12656
rect 41524 12481 41552 12650
rect 41510 12472 41566 12481
rect 41420 12436 41472 12442
rect 41510 12407 41566 12416
rect 41420 12378 41472 12384
rect 41432 11830 41460 12378
rect 41420 11824 41472 11830
rect 41420 11766 41472 11772
rect 41616 10742 41644 13631
rect 41604 10736 41656 10742
rect 41604 10678 41656 10684
rect 41510 10568 41566 10577
rect 41510 10503 41566 10512
rect 41328 10464 41380 10470
rect 41328 10406 41380 10412
rect 41420 9920 41472 9926
rect 41420 9862 41472 9868
rect 41432 9586 41460 9862
rect 41420 9580 41472 9586
rect 41420 9522 41472 9528
rect 41236 9376 41288 9382
rect 41236 9318 41288 9324
rect 41420 9104 41472 9110
rect 41420 9046 41472 9052
rect 41328 9036 41380 9042
rect 41328 8978 41380 8984
rect 41144 8968 41196 8974
rect 41144 8910 41196 8916
rect 41234 8800 41290 8809
rect 41234 8735 41290 8744
rect 41248 8634 41276 8735
rect 41236 8628 41288 8634
rect 41236 8570 41288 8576
rect 41340 8498 41368 8978
rect 41328 8492 41380 8498
rect 41328 8434 41380 8440
rect 41234 7576 41290 7585
rect 41234 7511 41290 7520
rect 41052 4480 41104 4486
rect 41052 4422 41104 4428
rect 41064 3534 41092 4422
rect 41144 4004 41196 4010
rect 41144 3946 41196 3952
rect 41156 3534 41184 3946
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 41144 3528 41196 3534
rect 41144 3470 41196 3476
rect 41144 3188 41196 3194
rect 41144 3130 41196 3136
rect 40960 1352 41012 1358
rect 40960 1294 41012 1300
rect 41156 800 41184 3130
rect 41248 2378 41276 7511
rect 41340 4554 41368 8434
rect 41432 4740 41460 9046
rect 41524 5302 41552 10503
rect 41604 9512 41656 9518
rect 41604 9454 41656 9460
rect 41616 9042 41644 9454
rect 41604 9036 41656 9042
rect 41604 8978 41656 8984
rect 41708 8498 41736 13926
rect 41972 13320 42024 13326
rect 42076 13308 42104 21354
rect 42156 17332 42208 17338
rect 42156 17274 42208 17280
rect 42168 16114 42196 17274
rect 42156 16108 42208 16114
rect 42156 16050 42208 16056
rect 42154 13696 42210 13705
rect 42154 13631 42210 13640
rect 42168 13326 42196 13631
rect 42024 13280 42104 13308
rect 42156 13320 42208 13326
rect 41972 13262 42024 13268
rect 42156 13262 42208 13268
rect 41880 12844 41932 12850
rect 41880 12786 41932 12792
rect 41788 12640 41840 12646
rect 41788 12582 41840 12588
rect 41800 12238 41828 12582
rect 41788 12232 41840 12238
rect 41788 12174 41840 12180
rect 41892 11898 41920 12786
rect 42064 12776 42116 12782
rect 42064 12718 42116 12724
rect 42076 12481 42104 12718
rect 42062 12472 42118 12481
rect 42062 12407 42118 12416
rect 41880 11892 41932 11898
rect 41880 11834 41932 11840
rect 42076 10470 42104 12407
rect 41788 10464 41840 10470
rect 41788 10406 41840 10412
rect 42064 10464 42116 10470
rect 42064 10406 42116 10412
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 41696 8288 41748 8294
rect 41696 8230 41748 8236
rect 41708 7886 41736 8230
rect 41800 8090 41828 10406
rect 41880 9716 41932 9722
rect 41880 9658 41932 9664
rect 41788 8084 41840 8090
rect 41788 8026 41840 8032
rect 41696 7880 41748 7886
rect 41696 7822 41748 7828
rect 41604 7404 41656 7410
rect 41604 7346 41656 7352
rect 41788 7404 41840 7410
rect 41788 7346 41840 7352
rect 41616 6934 41644 7346
rect 41604 6928 41656 6934
rect 41604 6870 41656 6876
rect 41800 6746 41828 7346
rect 41708 6730 41828 6746
rect 41696 6724 41828 6730
rect 41748 6718 41828 6724
rect 41696 6666 41748 6672
rect 41800 6322 41828 6718
rect 41788 6316 41840 6322
rect 41788 6258 41840 6264
rect 41696 6180 41748 6186
rect 41696 6122 41748 6128
rect 41708 5914 41736 6122
rect 41696 5908 41748 5914
rect 41696 5850 41748 5856
rect 41604 5636 41656 5642
rect 41604 5578 41656 5584
rect 41512 5296 41564 5302
rect 41512 5238 41564 5244
rect 41512 4752 41564 4758
rect 41432 4712 41512 4740
rect 41512 4694 41564 4700
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 41340 3466 41368 4490
rect 41512 4072 41564 4078
rect 41512 4014 41564 4020
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 41326 2680 41382 2689
rect 41326 2615 41328 2624
rect 41380 2615 41382 2624
rect 41328 2586 41380 2592
rect 41432 2446 41460 3878
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41236 2372 41288 2378
rect 41236 2314 41288 2320
rect 41524 2122 41552 4014
rect 41616 2854 41644 5578
rect 41696 5228 41748 5234
rect 41696 5170 41748 5176
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41432 2094 41552 2122
rect 41432 800 41460 2094
rect 41708 800 41736 5170
rect 41892 3126 41920 9658
rect 42260 9450 42288 56102
rect 42904 42090 42932 61066
rect 45376 61056 45428 61062
rect 45376 60998 45428 61004
rect 46112 61056 46164 61062
rect 46112 60998 46164 61004
rect 44180 60512 44232 60518
rect 44180 60454 44232 60460
rect 43260 60104 43312 60110
rect 43260 60046 43312 60052
rect 43272 59770 43300 60046
rect 43260 59764 43312 59770
rect 43260 59706 43312 59712
rect 43272 59634 43300 59706
rect 43260 59628 43312 59634
rect 43260 59570 43312 59576
rect 44192 55282 44220 60454
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 45388 54534 45416 60998
rect 45376 54528 45428 54534
rect 45376 54470 45428 54476
rect 46124 53650 46152 60998
rect 46676 60790 46704 63294
rect 47214 63200 47270 64000
rect 47950 63322 48006 64000
rect 47950 63294 48268 63322
rect 47950 63200 48006 63294
rect 46756 61328 46808 61334
rect 46756 61270 46808 61276
rect 46664 60784 46716 60790
rect 46664 60726 46716 60732
rect 46768 56370 46796 61270
rect 47228 61198 47256 63200
rect 47216 61192 47268 61198
rect 48240 61180 48268 63294
rect 48686 63200 48742 64000
rect 49422 63322 49478 64000
rect 49422 63294 49648 63322
rect 49422 63200 49478 63294
rect 48700 61198 48728 63200
rect 48964 61328 49016 61334
rect 48964 61270 49016 61276
rect 48320 61192 48372 61198
rect 48240 61152 48320 61180
rect 47216 61134 47268 61140
rect 48320 61134 48372 61140
rect 48688 61192 48740 61198
rect 48688 61134 48740 61140
rect 46940 61124 46992 61130
rect 46940 61066 46992 61072
rect 46848 61056 46900 61062
rect 46848 60998 46900 61004
rect 46860 60858 46888 60998
rect 46848 60852 46900 60858
rect 46848 60794 46900 60800
rect 46952 60654 46980 61066
rect 47584 61056 47636 61062
rect 47584 60998 47636 61004
rect 46940 60648 46992 60654
rect 46940 60590 46992 60596
rect 46756 56364 46808 56370
rect 46756 56306 46808 56312
rect 46112 53644 46164 53650
rect 46112 53586 46164 53592
rect 45008 50312 45060 50318
rect 45008 50254 45060 50260
rect 44916 45824 44968 45830
rect 44916 45766 44968 45772
rect 42892 42084 42944 42090
rect 42892 42026 42944 42032
rect 44088 40452 44140 40458
rect 44088 40394 44140 40400
rect 43444 35284 43496 35290
rect 43444 35226 43496 35232
rect 42432 25764 42484 25770
rect 42432 25706 42484 25712
rect 42340 15020 42392 15026
rect 42340 14962 42392 14968
rect 42352 14618 42380 14962
rect 42340 14612 42392 14618
rect 42340 14554 42392 14560
rect 42338 14104 42394 14113
rect 42338 14039 42394 14048
rect 42352 11898 42380 14039
rect 42340 11892 42392 11898
rect 42340 11834 42392 11840
rect 42352 11762 42380 11834
rect 42340 11756 42392 11762
rect 42340 11698 42392 11704
rect 42340 11620 42392 11626
rect 42340 11562 42392 11568
rect 42352 10810 42380 11562
rect 42340 10804 42392 10810
rect 42340 10746 42392 10752
rect 42248 9444 42300 9450
rect 42248 9386 42300 9392
rect 42248 7948 42300 7954
rect 42248 7890 42300 7896
rect 42156 7880 42208 7886
rect 42156 7822 42208 7828
rect 42168 7478 42196 7822
rect 42260 7721 42288 7890
rect 42246 7712 42302 7721
rect 42246 7647 42302 7656
rect 42156 7472 42208 7478
rect 42156 7414 42208 7420
rect 42064 7268 42116 7274
rect 42064 7210 42116 7216
rect 42076 6866 42104 7210
rect 42064 6860 42116 6866
rect 42064 6802 42116 6808
rect 42338 5536 42394 5545
rect 42338 5471 42394 5480
rect 42352 4622 42380 5471
rect 42340 4616 42392 4622
rect 42340 4558 42392 4564
rect 42248 4208 42300 4214
rect 42248 4150 42300 4156
rect 41970 4040 42026 4049
rect 41970 3975 42026 3984
rect 41984 3738 42012 3975
rect 41972 3732 42024 3738
rect 41972 3674 42024 3680
rect 42156 3528 42208 3534
rect 42154 3496 42156 3505
rect 42208 3496 42210 3505
rect 42154 3431 42210 3440
rect 41880 3120 41932 3126
rect 41880 3062 41932 3068
rect 41970 3088 42026 3097
rect 41970 3023 42026 3032
rect 41984 800 42012 3023
rect 42260 800 42288 4150
rect 42444 3126 42472 25706
rect 42524 22772 42576 22778
rect 42524 22714 42576 22720
rect 42536 4146 42564 22714
rect 43456 22094 43484 35226
rect 43536 25696 43588 25702
rect 43536 25638 43588 25644
rect 43364 22066 43484 22094
rect 42984 19168 43036 19174
rect 42984 19110 43036 19116
rect 42996 18834 43024 19110
rect 42984 18828 43036 18834
rect 42984 18770 43036 18776
rect 43076 18692 43128 18698
rect 43076 18634 43128 18640
rect 42984 18624 43036 18630
rect 42984 18566 43036 18572
rect 42800 18284 42852 18290
rect 42800 18226 42852 18232
rect 42812 17882 42840 18226
rect 42892 18216 42944 18222
rect 42892 18158 42944 18164
rect 42800 17876 42852 17882
rect 42800 17818 42852 17824
rect 42904 17678 42932 18158
rect 42892 17672 42944 17678
rect 42892 17614 42944 17620
rect 42616 17604 42668 17610
rect 42616 17546 42668 17552
rect 42628 16590 42656 17546
rect 42616 16584 42668 16590
rect 42616 16526 42668 16532
rect 42628 14958 42656 16526
rect 42904 15706 42932 17614
rect 42996 17610 43024 18566
rect 42984 17604 43036 17610
rect 42984 17546 43036 17552
rect 42984 17128 43036 17134
rect 43088 17116 43116 18634
rect 43168 17604 43220 17610
rect 43168 17546 43220 17552
rect 43036 17088 43116 17116
rect 42984 17070 43036 17076
rect 42996 16250 43024 17070
rect 43180 16522 43208 17546
rect 43260 16992 43312 16998
rect 43260 16934 43312 16940
rect 43272 16658 43300 16934
rect 43260 16652 43312 16658
rect 43260 16594 43312 16600
rect 43168 16516 43220 16522
rect 43168 16458 43220 16464
rect 42984 16244 43036 16250
rect 42984 16186 43036 16192
rect 43168 15972 43220 15978
rect 43168 15914 43220 15920
rect 42892 15700 42944 15706
rect 42892 15642 42944 15648
rect 42706 15328 42762 15337
rect 42706 15263 42762 15272
rect 42616 14952 42668 14958
rect 42616 14894 42668 14900
rect 42720 14618 42748 15263
rect 42708 14612 42760 14618
rect 42708 14554 42760 14560
rect 42706 14512 42762 14521
rect 42706 14447 42762 14456
rect 42720 14414 42748 14447
rect 42708 14408 42760 14414
rect 42708 14350 42760 14356
rect 43180 12782 43208 15914
rect 43260 15360 43312 15366
rect 43260 15302 43312 15308
rect 43272 14414 43300 15302
rect 43260 14408 43312 14414
rect 43260 14350 43312 14356
rect 43076 12776 43128 12782
rect 43076 12718 43128 12724
rect 43168 12776 43220 12782
rect 43168 12718 43220 12724
rect 42892 12640 42944 12646
rect 42892 12582 42944 12588
rect 42708 12300 42760 12306
rect 42708 12242 42760 12248
rect 42720 11762 42748 12242
rect 42904 11830 42932 12582
rect 43088 11898 43116 12718
rect 43272 12481 43300 14350
rect 43364 14346 43392 22066
rect 43444 15904 43496 15910
rect 43444 15846 43496 15852
rect 43456 15026 43484 15846
rect 43444 15020 43496 15026
rect 43444 14962 43496 14968
rect 43352 14340 43404 14346
rect 43352 14282 43404 14288
rect 43350 14104 43406 14113
rect 43350 14039 43406 14048
rect 43364 13938 43392 14039
rect 43352 13932 43404 13938
rect 43352 13874 43404 13880
rect 43444 13456 43496 13462
rect 43444 13398 43496 13404
rect 43352 12776 43404 12782
rect 43352 12718 43404 12724
rect 43258 12472 43314 12481
rect 43258 12407 43314 12416
rect 42984 11892 43036 11898
rect 42984 11834 43036 11840
rect 43076 11892 43128 11898
rect 43076 11834 43128 11840
rect 42892 11824 42944 11830
rect 42892 11766 42944 11772
rect 42708 11756 42760 11762
rect 42708 11698 42760 11704
rect 42616 11552 42668 11558
rect 42616 11494 42668 11500
rect 42628 10713 42656 11494
rect 42614 10704 42670 10713
rect 42614 10639 42670 10648
rect 42720 10130 42748 11698
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 42708 10124 42760 10130
rect 42708 10066 42760 10072
rect 42720 9586 42748 10066
rect 42812 9994 42840 10610
rect 42892 10464 42944 10470
rect 42892 10406 42944 10412
rect 42800 9988 42852 9994
rect 42800 9930 42852 9936
rect 42904 9654 42932 10406
rect 42892 9648 42944 9654
rect 42892 9590 42944 9596
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 42614 9072 42670 9081
rect 42614 9007 42670 9016
rect 42628 8362 42656 9007
rect 42720 8974 42748 9522
rect 42708 8968 42760 8974
rect 42708 8910 42760 8916
rect 42616 8356 42668 8362
rect 42616 8298 42668 8304
rect 42720 7886 42748 8910
rect 42996 8906 43024 11834
rect 43088 11665 43116 11834
rect 43168 11824 43220 11830
rect 43168 11766 43220 11772
rect 43074 11656 43130 11665
rect 43074 11591 43130 11600
rect 43180 11150 43208 11766
rect 43272 11150 43300 12407
rect 43168 11144 43220 11150
rect 43168 11086 43220 11092
rect 43260 11144 43312 11150
rect 43260 11086 43312 11092
rect 43180 10130 43208 11086
rect 43260 10736 43312 10742
rect 43260 10678 43312 10684
rect 43168 10124 43220 10130
rect 43168 10066 43220 10072
rect 43272 9704 43300 10678
rect 43364 10606 43392 12718
rect 43456 11762 43484 13398
rect 43444 11756 43496 11762
rect 43444 11698 43496 11704
rect 43444 11076 43496 11082
rect 43444 11018 43496 11024
rect 43456 10742 43484 11018
rect 43444 10736 43496 10742
rect 43444 10678 43496 10684
rect 43352 10600 43404 10606
rect 43352 10542 43404 10548
rect 43364 10130 43392 10542
rect 43352 10124 43404 10130
rect 43352 10066 43404 10072
rect 43352 9716 43404 9722
rect 43272 9676 43352 9704
rect 43352 9658 43404 9664
rect 42984 8900 43036 8906
rect 42984 8842 43036 8848
rect 42996 8430 43024 8842
rect 42984 8424 43036 8430
rect 42984 8366 43036 8372
rect 42708 7880 42760 7886
rect 42708 7822 42760 7828
rect 42616 7540 42668 7546
rect 42668 7500 42748 7528
rect 42616 7482 42668 7488
rect 42720 7410 42748 7500
rect 42708 7404 42760 7410
rect 42708 7346 42760 7352
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 42800 7268 42852 7274
rect 42800 7210 42852 7216
rect 42812 7002 42840 7210
rect 42904 7206 42932 7346
rect 43260 7336 43312 7342
rect 43260 7278 43312 7284
rect 42892 7200 42944 7206
rect 42892 7142 42944 7148
rect 42800 6996 42852 7002
rect 42800 6938 42852 6944
rect 42904 5794 42932 7142
rect 43272 6798 43300 7278
rect 43260 6792 43312 6798
rect 43260 6734 43312 6740
rect 43272 6458 43300 6734
rect 43260 6452 43312 6458
rect 43260 6394 43312 6400
rect 42812 5766 42932 5794
rect 42812 5710 42840 5766
rect 42800 5704 42852 5710
rect 42800 5646 42852 5652
rect 42892 5704 42944 5710
rect 42892 5646 42944 5652
rect 42708 5024 42760 5030
rect 42708 4966 42760 4972
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 42628 3369 42656 3538
rect 42720 3534 42748 4966
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 42812 4010 42840 4558
rect 42800 4004 42852 4010
rect 42800 3946 42852 3952
rect 42812 3534 42840 3946
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42800 3528 42852 3534
rect 42800 3470 42852 3476
rect 42614 3360 42670 3369
rect 42614 3295 42670 3304
rect 42432 3120 42484 3126
rect 42432 3062 42484 3068
rect 42798 2680 42854 2689
rect 42798 2615 42800 2624
rect 42852 2615 42854 2624
rect 42800 2586 42852 2592
rect 42904 2530 42932 5646
rect 43364 5370 43392 9658
rect 43444 6792 43496 6798
rect 43444 6734 43496 6740
rect 43456 5574 43484 6734
rect 43444 5568 43496 5574
rect 43444 5510 43496 5516
rect 43548 5370 43576 25638
rect 44100 22094 44128 40394
rect 44824 35216 44876 35222
rect 44824 35158 44876 35164
rect 44364 31884 44416 31890
rect 44364 31826 44416 31832
rect 43916 22066 44128 22094
rect 43916 19378 43944 22066
rect 44272 20868 44324 20874
rect 44272 20810 44324 20816
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 43628 18760 43680 18766
rect 43628 18702 43680 18708
rect 43640 18426 43668 18702
rect 43628 18420 43680 18426
rect 43628 18362 43680 18368
rect 43628 17332 43680 17338
rect 43628 17274 43680 17280
rect 43640 16658 43668 17274
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 43628 16652 43680 16658
rect 43628 16594 43680 16600
rect 43628 15020 43680 15026
rect 43628 14962 43680 14968
rect 43640 14074 43668 14962
rect 43720 14884 43772 14890
rect 43720 14826 43772 14832
rect 43732 14278 43760 14826
rect 43824 14414 43852 17138
rect 43812 14408 43864 14414
rect 43812 14350 43864 14356
rect 43720 14272 43772 14278
rect 43720 14214 43772 14220
rect 43628 14068 43680 14074
rect 43628 14010 43680 14016
rect 43732 14006 43760 14214
rect 43824 14113 43852 14350
rect 43810 14104 43866 14113
rect 43810 14039 43866 14048
rect 43720 14000 43772 14006
rect 43720 13942 43772 13948
rect 43812 13864 43864 13870
rect 43812 13806 43864 13812
rect 43628 13388 43680 13394
rect 43628 13330 43680 13336
rect 43640 12442 43668 13330
rect 43628 12436 43680 12442
rect 43628 12378 43680 12384
rect 43720 11756 43772 11762
rect 43720 11698 43772 11704
rect 43628 11280 43680 11286
rect 43626 11248 43628 11257
rect 43680 11248 43682 11257
rect 43626 11183 43682 11192
rect 43628 11076 43680 11082
rect 43628 11018 43680 11024
rect 43640 10062 43668 11018
rect 43628 10056 43680 10062
rect 43628 9998 43680 10004
rect 43628 8492 43680 8498
rect 43628 8434 43680 8440
rect 43640 7546 43668 8434
rect 43628 7540 43680 7546
rect 43628 7482 43680 7488
rect 43732 5914 43760 11698
rect 43824 8430 43852 13806
rect 43812 8424 43864 8430
rect 43812 8366 43864 8372
rect 43916 7478 43944 19314
rect 44088 18896 44140 18902
rect 44088 18838 44140 18844
rect 43996 18760 44048 18766
rect 43996 18702 44048 18708
rect 44008 17202 44036 18702
rect 44100 17678 44128 18838
rect 44284 18698 44312 20810
rect 44272 18692 44324 18698
rect 44272 18634 44324 18640
rect 44284 18426 44312 18634
rect 44272 18420 44324 18426
rect 44272 18362 44324 18368
rect 44180 18216 44232 18222
rect 44180 18158 44232 18164
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 43996 17196 44048 17202
rect 43996 17138 44048 17144
rect 44192 17134 44220 18158
rect 44376 17882 44404 31826
rect 44732 30184 44784 30190
rect 44732 30126 44784 30132
rect 44744 22094 44772 30126
rect 44652 22066 44772 22094
rect 44364 17876 44416 17882
rect 44364 17818 44416 17824
rect 44376 17270 44404 17818
rect 44456 17604 44508 17610
rect 44456 17546 44508 17552
rect 44364 17264 44416 17270
rect 44364 17206 44416 17212
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 43996 16992 44048 16998
rect 43996 16934 44048 16940
rect 44008 16436 44036 16934
rect 44088 16448 44140 16454
rect 44008 16408 44088 16436
rect 44008 16114 44036 16408
rect 44088 16390 44140 16396
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 44008 13870 44036 16050
rect 44192 15910 44220 17070
rect 44364 16652 44416 16658
rect 44468 16640 44496 17546
rect 44416 16612 44496 16640
rect 44364 16594 44416 16600
rect 44272 16176 44324 16182
rect 44272 16118 44324 16124
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44088 15496 44140 15502
rect 44088 15438 44140 15444
rect 44100 15026 44128 15438
rect 44192 15026 44220 15846
rect 44284 15162 44312 16118
rect 44376 15434 44404 16594
rect 44548 16244 44600 16250
rect 44548 16186 44600 16192
rect 44560 15502 44588 16186
rect 44548 15496 44600 15502
rect 44548 15438 44600 15444
rect 44364 15428 44416 15434
rect 44364 15370 44416 15376
rect 44272 15156 44324 15162
rect 44272 15098 44324 15104
rect 44088 15020 44140 15026
rect 44088 14962 44140 14968
rect 44180 15020 44232 15026
rect 44180 14962 44232 14968
rect 44088 14544 44140 14550
rect 44088 14486 44140 14492
rect 44100 13938 44128 14486
rect 44180 14408 44232 14414
rect 44376 14396 44404 15370
rect 44456 15156 44508 15162
rect 44456 15098 44508 15104
rect 44468 14482 44496 15098
rect 44456 14476 44508 14482
rect 44456 14418 44508 14424
rect 44232 14368 44404 14396
rect 44180 14350 44232 14356
rect 44376 14362 44404 14368
rect 44376 14346 44496 14362
rect 44376 14340 44508 14346
rect 44376 14334 44456 14340
rect 44456 14282 44508 14288
rect 44364 14272 44416 14278
rect 44364 14214 44416 14220
rect 44088 13932 44140 13938
rect 44088 13874 44140 13880
rect 43996 13864 44048 13870
rect 44100 13841 44128 13874
rect 43996 13806 44048 13812
rect 44086 13832 44142 13841
rect 44086 13767 44142 13776
rect 44376 12434 44404 14214
rect 44376 12406 44496 12434
rect 44086 11248 44142 11257
rect 44086 11183 44142 11192
rect 44100 11150 44128 11183
rect 44088 11144 44140 11150
rect 44088 11086 44140 11092
rect 43996 9512 44048 9518
rect 43996 9454 44048 9460
rect 44008 9110 44036 9454
rect 44270 9208 44326 9217
rect 44270 9143 44326 9152
rect 43996 9104 44048 9110
rect 43996 9046 44048 9052
rect 43904 7472 43956 7478
rect 43904 7414 43956 7420
rect 43810 6896 43866 6905
rect 43810 6831 43866 6840
rect 43824 6798 43852 6831
rect 43812 6792 43864 6798
rect 43812 6734 43864 6740
rect 43720 5908 43772 5914
rect 43720 5850 43772 5856
rect 43720 5772 43772 5778
rect 43720 5714 43772 5720
rect 43732 5642 43760 5714
rect 43720 5636 43772 5642
rect 43720 5578 43772 5584
rect 43812 5568 43864 5574
rect 43812 5510 43864 5516
rect 43352 5364 43404 5370
rect 43352 5306 43404 5312
rect 43536 5364 43588 5370
rect 43536 5306 43588 5312
rect 43536 5228 43588 5234
rect 43536 5170 43588 5176
rect 43258 4720 43314 4729
rect 43258 4655 43260 4664
rect 43312 4655 43314 4664
rect 43260 4626 43312 4632
rect 43548 4622 43576 5170
rect 43536 4616 43588 4622
rect 43536 4558 43588 4564
rect 43718 4584 43774 4593
rect 43168 4548 43220 4554
rect 43718 4519 43720 4528
rect 43168 4490 43220 4496
rect 43772 4519 43774 4528
rect 43720 4490 43772 4496
rect 42982 4176 43038 4185
rect 42982 4111 43038 4120
rect 42996 4078 43024 4111
rect 42984 4072 43036 4078
rect 42984 4014 43036 4020
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 42812 2502 42932 2530
rect 42524 1216 42576 1222
rect 42524 1158 42576 1164
rect 42536 800 42564 1158
rect 42812 800 42840 2502
rect 43088 800 43116 3674
rect 43180 3602 43208 4490
rect 43260 4480 43312 4486
rect 43260 4422 43312 4428
rect 43272 4146 43300 4422
rect 43824 4162 43852 5510
rect 44008 5409 44036 9046
rect 44088 8900 44140 8906
rect 44088 8842 44140 8848
rect 44100 8498 44128 8842
rect 44088 8492 44140 8498
rect 44088 8434 44140 8440
rect 44180 8424 44232 8430
rect 44180 8366 44232 8372
rect 44192 8294 44220 8366
rect 44180 8288 44232 8294
rect 44180 8230 44232 8236
rect 44284 7818 44312 9143
rect 44272 7812 44324 7818
rect 44272 7754 44324 7760
rect 44180 7744 44232 7750
rect 44180 7686 44232 7692
rect 44192 7478 44220 7686
rect 44180 7472 44232 7478
rect 44180 7414 44232 7420
rect 44364 5636 44416 5642
rect 44364 5578 44416 5584
rect 43994 5400 44050 5409
rect 43994 5335 44050 5344
rect 43996 5024 44048 5030
rect 43996 4966 44048 4972
rect 44008 4690 44036 4966
rect 44272 4820 44324 4826
rect 44272 4762 44324 4768
rect 43996 4684 44048 4690
rect 43996 4626 44048 4632
rect 43904 4480 43956 4486
rect 43904 4422 43956 4428
rect 43732 4146 43852 4162
rect 43260 4140 43312 4146
rect 43260 4082 43312 4088
rect 43720 4140 43852 4146
rect 43772 4134 43852 4140
rect 43720 4082 43772 4088
rect 43536 4072 43588 4078
rect 43350 4040 43406 4049
rect 43536 4014 43588 4020
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43350 3975 43406 3984
rect 43168 3596 43220 3602
rect 43168 3538 43220 3544
rect 43364 3534 43392 3975
rect 43548 3942 43576 4014
rect 43536 3936 43588 3942
rect 43536 3878 43588 3884
rect 43628 3936 43680 3942
rect 43628 3878 43680 3884
rect 43534 3632 43590 3641
rect 43534 3567 43590 3576
rect 43548 3534 43576 3567
rect 43352 3528 43404 3534
rect 43352 3470 43404 3476
rect 43536 3528 43588 3534
rect 43536 3470 43588 3476
rect 43260 3460 43312 3466
rect 43260 3402 43312 3408
rect 43272 3058 43300 3402
rect 43640 3058 43668 3878
rect 43824 3534 43852 4014
rect 43812 3528 43864 3534
rect 43812 3470 43864 3476
rect 43824 3058 43852 3470
rect 43260 3052 43312 3058
rect 43260 2994 43312 3000
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 43534 2408 43590 2417
rect 43444 2372 43496 2378
rect 43534 2343 43590 2352
rect 43444 2314 43496 2320
rect 43456 2106 43484 2314
rect 43548 2310 43576 2343
rect 43536 2304 43588 2310
rect 43916 2292 43944 4422
rect 44284 2666 44312 4762
rect 44376 3097 44404 5578
rect 44468 4078 44496 12406
rect 44548 9376 44600 9382
rect 44548 9318 44600 9324
rect 44560 8974 44588 9318
rect 44548 8968 44600 8974
rect 44548 8910 44600 8916
rect 44546 7984 44602 7993
rect 44546 7919 44602 7928
rect 44560 4486 44588 7919
rect 44548 4480 44600 4486
rect 44548 4422 44600 4428
rect 44546 4176 44602 4185
rect 44546 4111 44548 4120
rect 44600 4111 44602 4120
rect 44548 4082 44600 4088
rect 44456 4072 44508 4078
rect 44456 4014 44508 4020
rect 44548 4004 44600 4010
rect 44548 3946 44600 3952
rect 44560 3602 44588 3946
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 44548 3460 44600 3466
rect 44548 3402 44600 3408
rect 44362 3088 44418 3097
rect 44362 3023 44418 3032
rect 44456 3052 44508 3058
rect 44456 2994 44508 3000
rect 44362 2952 44418 2961
rect 44362 2887 44418 2896
rect 43536 2246 43588 2252
rect 43640 2264 43944 2292
rect 44192 2638 44312 2666
rect 43444 2100 43496 2106
rect 43444 2042 43496 2048
rect 43352 1488 43404 1494
rect 43352 1430 43404 1436
rect 43364 800 43392 1430
rect 43640 800 43668 2264
rect 43904 2100 43956 2106
rect 43904 2042 43956 2048
rect 43916 800 43944 2042
rect 44192 800 44220 2638
rect 44376 2514 44404 2887
rect 44364 2508 44416 2514
rect 44364 2450 44416 2456
rect 44468 800 44496 2994
rect 44560 1222 44588 3402
rect 44652 3194 44680 22066
rect 44732 15020 44784 15026
rect 44732 14962 44784 14968
rect 44744 14074 44772 14962
rect 44836 14550 44864 35158
rect 44824 14544 44876 14550
rect 44824 14486 44876 14492
rect 44824 14272 44876 14278
rect 44824 14214 44876 14220
rect 44732 14068 44784 14074
rect 44732 14010 44784 14016
rect 44836 13938 44864 14214
rect 44824 13932 44876 13938
rect 44824 13874 44876 13880
rect 44928 9654 44956 45766
rect 45020 33318 45048 50254
rect 46296 47796 46348 47802
rect 46296 47738 46348 47744
rect 45836 38956 45888 38962
rect 45836 38898 45888 38904
rect 45100 34944 45152 34950
rect 45100 34886 45152 34892
rect 45008 33312 45060 33318
rect 45008 33254 45060 33260
rect 45112 20942 45140 34886
rect 45652 26376 45704 26382
rect 45652 26318 45704 26324
rect 45100 20936 45152 20942
rect 45100 20878 45152 20884
rect 45560 18760 45612 18766
rect 45560 18702 45612 18708
rect 45572 17882 45600 18702
rect 45560 17876 45612 17882
rect 45560 17818 45612 17824
rect 45560 17672 45612 17678
rect 45480 17632 45560 17660
rect 45480 16998 45508 17632
rect 45560 17614 45612 17620
rect 45664 17338 45692 26318
rect 45744 18624 45796 18630
rect 45744 18566 45796 18572
rect 45756 18358 45784 18566
rect 45744 18352 45796 18358
rect 45744 18294 45796 18300
rect 45652 17332 45704 17338
rect 45652 17274 45704 17280
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 45468 16992 45520 16998
rect 45468 16934 45520 16940
rect 45480 16182 45508 16934
rect 45572 16726 45600 17138
rect 45560 16720 45612 16726
rect 45560 16662 45612 16668
rect 45468 16176 45520 16182
rect 45468 16118 45520 16124
rect 45192 15496 45244 15502
rect 45192 15438 45244 15444
rect 45204 13530 45232 15438
rect 45480 15026 45508 16118
rect 45744 16108 45796 16114
rect 45744 16050 45796 16056
rect 45756 15706 45784 16050
rect 45744 15700 45796 15706
rect 45744 15642 45796 15648
rect 45468 15020 45520 15026
rect 45468 14962 45520 14968
rect 45468 14408 45520 14414
rect 45468 14350 45520 14356
rect 45192 13524 45244 13530
rect 45192 13466 45244 13472
rect 45480 10470 45508 14350
rect 45468 10464 45520 10470
rect 45468 10406 45520 10412
rect 45100 9988 45152 9994
rect 45100 9930 45152 9936
rect 44916 9648 44968 9654
rect 44916 9590 44968 9596
rect 45112 9518 45140 9930
rect 45192 9920 45244 9926
rect 45192 9862 45244 9868
rect 45100 9512 45152 9518
rect 45100 9454 45152 9460
rect 44732 9444 44784 9450
rect 44732 9386 44784 9392
rect 44744 4162 44772 9386
rect 44916 8084 44968 8090
rect 44916 8026 44968 8032
rect 44824 7404 44876 7410
rect 44824 7346 44876 7352
rect 44836 7206 44864 7346
rect 44824 7200 44876 7206
rect 44824 7142 44876 7148
rect 44836 5234 44864 7142
rect 44824 5228 44876 5234
rect 44824 5170 44876 5176
rect 44928 5166 44956 8026
rect 45112 6390 45140 9454
rect 45100 6384 45152 6390
rect 45100 6326 45152 6332
rect 45008 6248 45060 6254
rect 45008 6190 45060 6196
rect 45020 5370 45048 6190
rect 45008 5364 45060 5370
rect 45008 5306 45060 5312
rect 44916 5160 44968 5166
rect 44916 5102 44968 5108
rect 45008 5160 45060 5166
rect 45008 5102 45060 5108
rect 44928 4758 44956 5102
rect 44916 4752 44968 4758
rect 44916 4694 44968 4700
rect 44744 4134 44864 4162
rect 44732 4004 44784 4010
rect 44732 3946 44784 3952
rect 44640 3188 44692 3194
rect 44640 3130 44692 3136
rect 44548 1216 44600 1222
rect 44548 1158 44600 1164
rect 44744 800 44772 3946
rect 44836 2961 44864 4134
rect 45020 3534 45048 5102
rect 45100 4208 45152 4214
rect 45100 4150 45152 4156
rect 45112 3738 45140 4150
rect 45204 3738 45232 9862
rect 45480 7886 45508 10406
rect 45468 7880 45520 7886
rect 45468 7822 45520 7828
rect 45284 6724 45336 6730
rect 45284 6666 45336 6672
rect 45296 5914 45324 6666
rect 45284 5908 45336 5914
rect 45284 5850 45336 5856
rect 45376 5364 45428 5370
rect 45376 5306 45428 5312
rect 45284 5228 45336 5234
rect 45284 5170 45336 5176
rect 45296 4060 45324 5170
rect 45388 4570 45416 5306
rect 45480 4690 45508 7822
rect 45652 5228 45704 5234
rect 45652 5170 45704 5176
rect 45744 5228 45796 5234
rect 45744 5170 45796 5176
rect 45558 4720 45614 4729
rect 45468 4684 45520 4690
rect 45558 4655 45614 4664
rect 45468 4626 45520 4632
rect 45572 4622 45600 4655
rect 45560 4616 45612 4622
rect 45388 4554 45508 4570
rect 45560 4558 45612 4564
rect 45388 4548 45520 4554
rect 45388 4542 45468 4548
rect 45468 4490 45520 4496
rect 45376 4072 45428 4078
rect 45296 4032 45376 4060
rect 45376 4014 45428 4020
rect 45664 4010 45692 5170
rect 45756 4826 45784 5170
rect 45744 4820 45796 4826
rect 45744 4762 45796 4768
rect 45744 4208 45796 4214
rect 45744 4150 45796 4156
rect 45652 4004 45704 4010
rect 45652 3946 45704 3952
rect 45100 3732 45152 3738
rect 45100 3674 45152 3680
rect 45192 3732 45244 3738
rect 45192 3674 45244 3680
rect 45008 3528 45060 3534
rect 45008 3470 45060 3476
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 45204 3194 45232 3334
rect 45192 3188 45244 3194
rect 45192 3130 45244 3136
rect 45480 3126 45508 3402
rect 45468 3120 45520 3126
rect 45468 3062 45520 3068
rect 45284 2984 45336 2990
rect 44822 2952 44878 2961
rect 44822 2887 44878 2896
rect 45020 2932 45284 2938
rect 45020 2926 45336 2932
rect 45020 2910 45324 2926
rect 45020 800 45048 2910
rect 45284 2848 45336 2854
rect 45284 2790 45336 2796
rect 45296 800 45324 2790
rect 45560 2372 45612 2378
rect 45560 2314 45612 2320
rect 45572 800 45600 2314
rect 45756 2106 45784 4150
rect 45848 2650 45876 38898
rect 46204 36372 46256 36378
rect 46204 36314 46256 36320
rect 46020 20936 46072 20942
rect 46020 20878 46072 20884
rect 45928 18624 45980 18630
rect 45928 18566 45980 18572
rect 45940 18426 45968 18566
rect 45928 18420 45980 18426
rect 45928 18362 45980 18368
rect 45926 9616 45982 9625
rect 45926 9551 45982 9560
rect 45940 4282 45968 9551
rect 45928 4276 45980 4282
rect 45928 4218 45980 4224
rect 46032 3738 46060 20878
rect 46112 19304 46164 19310
rect 46112 19246 46164 19252
rect 46124 18834 46152 19246
rect 46112 18828 46164 18834
rect 46112 18770 46164 18776
rect 46216 18086 46244 36314
rect 46204 18080 46256 18086
rect 46204 18022 46256 18028
rect 46308 17542 46336 47738
rect 47400 32496 47452 32502
rect 47400 32438 47452 32444
rect 46940 31340 46992 31346
rect 46940 31282 46992 31288
rect 46480 31136 46532 31142
rect 46480 31078 46532 31084
rect 46388 30252 46440 30258
rect 46388 30194 46440 30200
rect 46296 17536 46348 17542
rect 46296 17478 46348 17484
rect 46204 16040 46256 16046
rect 46204 15982 46256 15988
rect 46216 15366 46244 15982
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 46204 12164 46256 12170
rect 46204 12106 46256 12112
rect 46216 11082 46244 12106
rect 46204 11076 46256 11082
rect 46204 11018 46256 11024
rect 46296 10804 46348 10810
rect 46296 10746 46348 10752
rect 46308 10538 46336 10746
rect 46296 10532 46348 10538
rect 46296 10474 46348 10480
rect 46020 3732 46072 3738
rect 46020 3674 46072 3680
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 45836 2372 45888 2378
rect 45836 2314 45888 2320
rect 45744 2100 45796 2106
rect 45744 2042 45796 2048
rect 45848 800 45876 2314
rect 46032 1698 46060 3470
rect 46400 3194 46428 30194
rect 46492 23322 46520 31078
rect 46756 24880 46808 24886
rect 46756 24822 46808 24828
rect 46480 23316 46532 23322
rect 46480 23258 46532 23264
rect 46768 18426 46796 24822
rect 46848 18692 46900 18698
rect 46848 18634 46900 18640
rect 46756 18420 46808 18426
rect 46756 18362 46808 18368
rect 46768 17610 46796 18362
rect 46860 18290 46888 18634
rect 46848 18284 46900 18290
rect 46848 18226 46900 18232
rect 46756 17604 46808 17610
rect 46756 17546 46808 17552
rect 46860 16658 46888 18226
rect 46848 16652 46900 16658
rect 46848 16594 46900 16600
rect 46756 16448 46808 16454
rect 46756 16390 46808 16396
rect 46480 16108 46532 16114
rect 46480 16050 46532 16056
rect 46492 15065 46520 16050
rect 46572 15904 46624 15910
rect 46572 15846 46624 15852
rect 46478 15056 46534 15065
rect 46478 14991 46534 15000
rect 46584 14346 46612 15846
rect 46664 15496 46716 15502
rect 46664 15438 46716 15444
rect 46676 15094 46704 15438
rect 46768 15434 46796 16390
rect 46860 16046 46888 16594
rect 46848 16040 46900 16046
rect 46848 15982 46900 15988
rect 46756 15428 46808 15434
rect 46756 15370 46808 15376
rect 46664 15088 46716 15094
rect 46664 15030 46716 15036
rect 46768 14618 46796 15370
rect 46756 14612 46808 14618
rect 46756 14554 46808 14560
rect 46756 14476 46808 14482
rect 46756 14418 46808 14424
rect 46572 14340 46624 14346
rect 46572 14282 46624 14288
rect 46768 13938 46796 14418
rect 46848 14272 46900 14278
rect 46848 14214 46900 14220
rect 46860 14006 46888 14214
rect 46848 14000 46900 14006
rect 46848 13942 46900 13948
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 46756 13932 46808 13938
rect 46756 13874 46808 13880
rect 46676 12986 46704 13874
rect 46664 12980 46716 12986
rect 46664 12922 46716 12928
rect 46754 11520 46810 11529
rect 46754 11455 46810 11464
rect 46768 4146 46796 11455
rect 46756 4140 46808 4146
rect 46756 4082 46808 4088
rect 46572 4004 46624 4010
rect 46572 3946 46624 3952
rect 46584 3505 46612 3946
rect 46570 3496 46626 3505
rect 46570 3431 46626 3440
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 46388 3188 46440 3194
rect 46388 3130 46440 3136
rect 46112 3052 46164 3058
rect 46112 2994 46164 3000
rect 46020 1692 46072 1698
rect 46020 1634 46072 1640
rect 46124 800 46152 2994
rect 46388 2440 46440 2446
rect 46388 2382 46440 2388
rect 46400 800 46428 2382
rect 46676 800 46704 3402
rect 46952 2650 46980 31282
rect 47032 18080 47084 18086
rect 47032 18022 47084 18028
rect 47044 3670 47072 18022
rect 47124 15496 47176 15502
rect 47124 15438 47176 15444
rect 47136 14822 47164 15438
rect 47216 15428 47268 15434
rect 47216 15370 47268 15376
rect 47124 14816 47176 14822
rect 47124 14758 47176 14764
rect 47228 10742 47256 15370
rect 47216 10736 47268 10742
rect 47216 10678 47268 10684
rect 47032 3664 47084 3670
rect 47032 3606 47084 3612
rect 47124 3460 47176 3466
rect 47124 3402 47176 3408
rect 47032 3052 47084 3058
rect 47032 2994 47084 3000
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 47044 1578 47072 2994
rect 46952 1550 47072 1578
rect 46952 800 46980 1550
rect 47136 1494 47164 3402
rect 47412 3194 47440 32438
rect 47596 24274 47624 60998
rect 48976 40934 49004 61270
rect 49620 61180 49648 63294
rect 50158 63200 50214 64000
rect 50894 63322 50950 64000
rect 50894 63294 51028 63322
rect 50894 63200 50950 63294
rect 49700 61192 49752 61198
rect 49620 61152 49700 61180
rect 49700 61134 49752 61140
rect 50068 61056 50120 61062
rect 50068 60998 50120 61004
rect 50080 55214 50108 60998
rect 50172 60790 50200 63200
rect 51000 61180 51028 63294
rect 51630 63200 51686 64000
rect 52366 63200 52422 64000
rect 53102 63322 53158 64000
rect 53838 63322 53894 64000
rect 54574 63322 54630 64000
rect 55310 63322 55366 64000
rect 53102 63294 53236 63322
rect 53102 63200 53158 63294
rect 51448 61736 51500 61742
rect 51448 61678 51500 61684
rect 51460 61402 51488 61678
rect 51448 61396 51500 61402
rect 51448 61338 51500 61344
rect 51644 61198 51672 63200
rect 51080 61192 51132 61198
rect 51000 61152 51080 61180
rect 51080 61134 51132 61140
rect 51632 61192 51684 61198
rect 51632 61134 51684 61140
rect 51816 61056 51868 61062
rect 51816 60998 51868 61004
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 50160 60784 50212 60790
rect 50160 60726 50212 60732
rect 50436 60512 50488 60518
rect 50436 60454 50488 60460
rect 50448 60042 50476 60454
rect 50436 60036 50488 60042
rect 50436 59978 50488 59984
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50080 55186 50200 55214
rect 48964 40928 49016 40934
rect 48964 40870 49016 40876
rect 47676 39092 47728 39098
rect 47676 39034 47728 39040
rect 47584 24268 47636 24274
rect 47584 24210 47636 24216
rect 47492 18352 47544 18358
rect 47492 18294 47544 18300
rect 47504 17678 47532 18294
rect 47492 17672 47544 17678
rect 47492 17614 47544 17620
rect 47504 15094 47532 17614
rect 47492 15088 47544 15094
rect 47492 15030 47544 15036
rect 47504 13938 47532 15030
rect 47492 13932 47544 13938
rect 47492 13874 47544 13880
rect 47688 6934 47716 39034
rect 49056 38344 49108 38350
rect 49056 38286 49108 38292
rect 47952 37800 48004 37806
rect 47952 37742 48004 37748
rect 47768 35080 47820 35086
rect 47768 35022 47820 35028
rect 47780 20874 47808 35022
rect 47768 20868 47820 20874
rect 47768 20810 47820 20816
rect 47860 19984 47912 19990
rect 47860 19926 47912 19932
rect 47768 19440 47820 19446
rect 47766 19408 47768 19417
rect 47820 19408 47822 19417
rect 47872 19378 47900 19926
rect 47766 19343 47822 19352
rect 47860 19372 47912 19378
rect 47860 19314 47912 19320
rect 47676 6928 47728 6934
rect 47676 6870 47728 6876
rect 47400 3188 47452 3194
rect 47400 3130 47452 3136
rect 47492 3120 47544 3126
rect 47492 3062 47544 3068
rect 47216 2372 47268 2378
rect 47216 2314 47268 2320
rect 47124 1488 47176 1494
rect 47124 1430 47176 1436
rect 47228 800 47256 2314
rect 47504 800 47532 3062
rect 47964 2650 47992 37742
rect 48964 37256 49016 37262
rect 48964 37198 49016 37204
rect 48780 29300 48832 29306
rect 48780 29242 48832 29248
rect 48136 20052 48188 20058
rect 48136 19994 48188 20000
rect 48148 19446 48176 19994
rect 48596 19848 48648 19854
rect 48596 19790 48648 19796
rect 48504 19712 48556 19718
rect 48504 19654 48556 19660
rect 48226 19544 48282 19553
rect 48226 19479 48228 19488
rect 48280 19479 48282 19488
rect 48228 19450 48280 19456
rect 48136 19440 48188 19446
rect 48188 19388 48452 19394
rect 48136 19382 48452 19388
rect 48044 19372 48096 19378
rect 48148 19366 48452 19382
rect 48044 19314 48096 19320
rect 48056 18902 48084 19314
rect 48136 19236 48188 19242
rect 48136 19178 48188 19184
rect 48148 19145 48176 19178
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48044 18896 48096 18902
rect 48044 18838 48096 18844
rect 48056 18698 48084 18838
rect 48228 18760 48280 18766
rect 48226 18728 48228 18737
rect 48280 18728 48282 18737
rect 48044 18692 48096 18698
rect 48044 18634 48096 18640
rect 48136 18692 48188 18698
rect 48226 18663 48282 18672
rect 48136 18634 48188 18640
rect 48056 17610 48084 18634
rect 48148 18426 48176 18634
rect 48136 18420 48188 18426
rect 48136 18362 48188 18368
rect 48240 18358 48268 18663
rect 48228 18352 48280 18358
rect 48228 18294 48280 18300
rect 48136 18216 48188 18222
rect 48136 18158 48188 18164
rect 48148 17746 48176 18158
rect 48136 17740 48188 17746
rect 48136 17682 48188 17688
rect 48044 17604 48096 17610
rect 48044 17546 48096 17552
rect 48056 15434 48084 17546
rect 48148 17134 48176 17682
rect 48424 17490 48452 19366
rect 48516 17610 48544 19654
rect 48608 19174 48636 19790
rect 48686 19544 48742 19553
rect 48686 19479 48742 19488
rect 48700 19446 48728 19479
rect 48688 19440 48740 19446
rect 48688 19382 48740 19388
rect 48596 19168 48648 19174
rect 48596 19110 48648 19116
rect 48594 18864 48650 18873
rect 48594 18799 48596 18808
rect 48648 18799 48650 18808
rect 48596 18770 48648 18776
rect 48688 18760 48740 18766
rect 48688 18702 48740 18708
rect 48700 18630 48728 18702
rect 48688 18624 48740 18630
rect 48688 18566 48740 18572
rect 48504 17604 48556 17610
rect 48504 17546 48556 17552
rect 48596 17604 48648 17610
rect 48596 17546 48648 17552
rect 48608 17490 48636 17546
rect 48424 17462 48636 17490
rect 48136 17128 48188 17134
rect 48136 17070 48188 17076
rect 48148 16658 48176 17070
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48148 15706 48176 16594
rect 48688 16516 48740 16522
rect 48688 16458 48740 16464
rect 48700 16250 48728 16458
rect 48688 16244 48740 16250
rect 48688 16186 48740 16192
rect 48136 15700 48188 15706
rect 48136 15642 48188 15648
rect 48044 15428 48096 15434
rect 48044 15370 48096 15376
rect 48228 15088 48280 15094
rect 48228 15030 48280 15036
rect 48136 14340 48188 14346
rect 48136 14282 48188 14288
rect 48148 14074 48176 14282
rect 48240 14074 48268 15030
rect 48136 14068 48188 14074
rect 48136 14010 48188 14016
rect 48228 14068 48280 14074
rect 48228 14010 48280 14016
rect 48792 7698 48820 29242
rect 48976 20058 49004 37198
rect 49068 24886 49096 38286
rect 50172 35290 50200 55186
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50896 44872 50948 44878
rect 50896 44814 50948 44820
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50804 43784 50856 43790
rect 50804 43726 50856 43732
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50160 35284 50212 35290
rect 50160 35226 50212 35232
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50712 34740 50764 34746
rect 50712 34682 50764 34688
rect 49332 33856 49384 33862
rect 49332 33798 49384 33804
rect 49056 24880 49108 24886
rect 49056 24822 49108 24828
rect 48964 20052 49016 20058
rect 48964 19994 49016 20000
rect 48872 19916 48924 19922
rect 48872 19858 48924 19864
rect 48884 19378 48912 19858
rect 48964 19508 49016 19514
rect 48964 19450 49016 19456
rect 48976 19417 49004 19450
rect 48962 19408 49018 19417
rect 48872 19372 48924 19378
rect 48962 19343 49018 19352
rect 49056 19372 49108 19378
rect 48872 19314 48924 19320
rect 49056 19314 49108 19320
rect 48884 16114 48912 19314
rect 49068 18970 49096 19314
rect 49148 19304 49200 19310
rect 49148 19246 49200 19252
rect 49056 18964 49108 18970
rect 49056 18906 49108 18912
rect 49160 18834 49188 19246
rect 49240 19168 49292 19174
rect 49240 19110 49292 19116
rect 49148 18828 49200 18834
rect 49148 18770 49200 18776
rect 49160 18737 49188 18770
rect 49146 18728 49202 18737
rect 49146 18663 49202 18672
rect 49252 18358 49280 19110
rect 49240 18352 49292 18358
rect 49240 18294 49292 18300
rect 49240 17536 49292 17542
rect 49240 17478 49292 17484
rect 49252 16114 49280 17478
rect 48872 16108 48924 16114
rect 48872 16050 48924 16056
rect 49240 16108 49292 16114
rect 49240 16050 49292 16056
rect 48884 15570 48912 16050
rect 48872 15564 48924 15570
rect 48872 15506 48924 15512
rect 48884 13938 48912 15506
rect 48872 13932 48924 13938
rect 48872 13874 48924 13880
rect 49240 13728 49292 13734
rect 49240 13670 49292 13676
rect 48964 13184 49016 13190
rect 48964 13126 49016 13132
rect 48976 10849 49004 13126
rect 48962 10840 49018 10849
rect 48962 10775 49018 10784
rect 48792 7670 49096 7698
rect 48596 6180 48648 6186
rect 48596 6122 48648 6128
rect 48228 4820 48280 4826
rect 48228 4762 48280 4768
rect 48240 4146 48268 4762
rect 48412 4480 48464 4486
rect 48412 4422 48464 4428
rect 48424 4146 48452 4422
rect 48228 4140 48280 4146
rect 48228 4082 48280 4088
rect 48412 4140 48464 4146
rect 48412 4082 48464 4088
rect 48608 3738 48636 6122
rect 48872 4208 48924 4214
rect 48872 4150 48924 4156
rect 48596 3732 48648 3738
rect 48596 3674 48648 3680
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 48042 3360 48098 3369
rect 48042 3295 48098 3304
rect 48056 3194 48084 3295
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 48148 3058 48176 3402
rect 48136 3052 48188 3058
rect 48136 2994 48188 3000
rect 48596 3052 48648 3058
rect 48596 2994 48648 3000
rect 48044 2984 48096 2990
rect 48044 2926 48096 2932
rect 47952 2644 48004 2650
rect 47952 2586 48004 2592
rect 48056 2496 48084 2926
rect 47780 2468 48084 2496
rect 47780 800 47808 2468
rect 48044 2372 48096 2378
rect 48044 2314 48096 2320
rect 48056 800 48084 2314
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 48332 800 48360 2246
rect 48608 800 48636 2994
rect 48884 800 48912 4150
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48976 2854 49004 2994
rect 49068 2854 49096 7670
rect 49252 4146 49280 13670
rect 49344 12434 49372 33798
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50160 24336 50212 24342
rect 50160 24278 50212 24284
rect 49884 18692 49936 18698
rect 49884 18634 49936 18640
rect 49424 18624 49476 18630
rect 49424 18566 49476 18572
rect 49436 18290 49464 18566
rect 49424 18284 49476 18290
rect 49424 18226 49476 18232
rect 49700 18080 49752 18086
rect 49700 18022 49752 18028
rect 49712 17270 49740 18022
rect 49896 17338 49924 18634
rect 49976 17604 50028 17610
rect 49976 17546 50028 17552
rect 49884 17332 49936 17338
rect 49884 17274 49936 17280
rect 49700 17264 49752 17270
rect 49700 17206 49752 17212
rect 49700 16448 49752 16454
rect 49700 16390 49752 16396
rect 49712 16182 49740 16390
rect 49988 16250 50016 17546
rect 49976 16244 50028 16250
rect 49976 16186 50028 16192
rect 49700 16176 49752 16182
rect 49700 16118 49752 16124
rect 49424 16040 49476 16046
rect 49424 15982 49476 15988
rect 49436 15502 49464 15982
rect 49424 15496 49476 15502
rect 49424 15438 49476 15444
rect 49792 15496 49844 15502
rect 49792 15438 49844 15444
rect 49804 14890 49832 15438
rect 49792 14884 49844 14890
rect 49792 14826 49844 14832
rect 49700 14816 49752 14822
rect 49700 14758 49752 14764
rect 49344 12406 49464 12434
rect 49240 4140 49292 4146
rect 49240 4082 49292 4088
rect 49330 3904 49386 3913
rect 49330 3839 49386 3848
rect 49344 3738 49372 3839
rect 49332 3732 49384 3738
rect 49332 3674 49384 3680
rect 49148 3528 49200 3534
rect 49148 3470 49200 3476
rect 48964 2848 49016 2854
rect 48964 2790 49016 2796
rect 49056 2848 49108 2854
rect 49056 2790 49108 2796
rect 49160 800 49188 3470
rect 49436 2650 49464 12406
rect 49712 10810 49740 14758
rect 50068 12708 50120 12714
rect 50068 12650 50120 12656
rect 49700 10804 49752 10810
rect 49700 10746 49752 10752
rect 49516 10736 49568 10742
rect 49516 10678 49568 10684
rect 49528 10266 49556 10678
rect 49516 10260 49568 10266
rect 49516 10202 49568 10208
rect 49698 8120 49754 8129
rect 49698 8055 49754 8064
rect 49712 7886 49740 8055
rect 49700 7880 49752 7886
rect 49700 7822 49752 7828
rect 50080 3738 50108 12650
rect 50068 3732 50120 3738
rect 50068 3674 50120 3680
rect 49700 3664 49752 3670
rect 49698 3632 49700 3641
rect 49752 3632 49754 3641
rect 49698 3567 49754 3576
rect 49516 3460 49568 3466
rect 49516 3402 49568 3408
rect 49424 2644 49476 2650
rect 49424 2586 49476 2592
rect 49528 1714 49556 3402
rect 49698 3224 49754 3233
rect 49698 3159 49754 3168
rect 49712 2854 49740 3159
rect 49884 3120 49936 3126
rect 49884 3062 49936 3068
rect 49700 2848 49752 2854
rect 49700 2790 49752 2796
rect 49436 1686 49556 1714
rect 49436 800 49464 1686
rect 49896 1578 49924 3062
rect 50172 2650 50200 24278
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50724 18698 50752 34682
rect 50712 18692 50764 18698
rect 50712 18634 50764 18640
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50816 16454 50844 43726
rect 50804 16448 50856 16454
rect 50804 16390 50856 16396
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50712 15360 50764 15366
rect 50712 15302 50764 15308
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50724 15094 50752 15302
rect 50712 15088 50764 15094
rect 50712 15030 50764 15036
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50804 13864 50856 13870
rect 50804 13806 50856 13812
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50618 11112 50674 11121
rect 50618 11047 50620 11056
rect 50672 11047 50674 11056
rect 50620 11018 50672 11024
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50620 4208 50672 4214
rect 50620 4150 50672 4156
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50252 3188 50304 3194
rect 50252 3130 50304 3136
rect 50160 2644 50212 2650
rect 50160 2586 50212 2592
rect 49976 2372 50028 2378
rect 49976 2314 50028 2320
rect 49712 1550 49924 1578
rect 49712 800 49740 1550
rect 49988 800 50016 2314
rect 50264 2292 50292 3130
rect 50172 2264 50292 2292
rect 50172 1714 50200 2264
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1986 50660 4150
rect 50816 4146 50844 13806
rect 50908 11830 50936 44814
rect 51724 41608 51776 41614
rect 51724 41550 51776 41556
rect 50988 28552 51040 28558
rect 50988 28494 51040 28500
rect 51000 14890 51028 28494
rect 51736 17882 51764 41550
rect 51724 17876 51776 17882
rect 51724 17818 51776 17824
rect 50988 14884 51040 14890
rect 50988 14826 51040 14832
rect 51080 13320 51132 13326
rect 51080 13262 51132 13268
rect 50896 11824 50948 11830
rect 50896 11766 50948 11772
rect 51092 7478 51120 13262
rect 51724 10464 51776 10470
rect 51724 10406 51776 10412
rect 51080 7472 51132 7478
rect 51080 7414 51132 7420
rect 51262 6760 51318 6769
rect 51262 6695 51318 6704
rect 50804 4140 50856 4146
rect 50804 4082 50856 4088
rect 50896 4004 50948 4010
rect 50896 3946 50948 3952
rect 50712 3528 50764 3534
rect 50712 3470 50764 3476
rect 50724 3194 50752 3470
rect 50804 3460 50856 3466
rect 50804 3402 50856 3408
rect 50712 3188 50764 3194
rect 50712 3130 50764 3136
rect 50540 1958 50660 1986
rect 50172 1686 50292 1714
rect 50264 800 50292 1686
rect 50540 800 50568 1958
rect 50816 800 50844 3402
rect 50908 2990 50936 3946
rect 51276 3194 51304 6695
rect 51356 4208 51408 4214
rect 51356 4150 51408 4156
rect 51264 3188 51316 3194
rect 51264 3130 51316 3136
rect 51172 3052 51224 3058
rect 51172 2994 51224 3000
rect 50896 2984 50948 2990
rect 50896 2926 50948 2932
rect 51184 1714 51212 2994
rect 51264 2304 51316 2310
rect 51264 2246 51316 2252
rect 51276 1970 51304 2246
rect 51264 1964 51316 1970
rect 51264 1906 51316 1912
rect 51092 1686 51212 1714
rect 51092 800 51120 1686
rect 51368 800 51396 4150
rect 51736 4146 51764 10406
rect 51828 10305 51856 60998
rect 52380 60874 52408 63200
rect 53208 61198 53236 63294
rect 53838 63294 54156 63322
rect 53838 63200 53894 63294
rect 54128 61198 54156 63294
rect 54574 63294 54708 63322
rect 54574 63200 54630 63294
rect 53196 61192 53248 61198
rect 53196 61134 53248 61140
rect 54116 61192 54168 61198
rect 54116 61134 54168 61140
rect 54300 61056 54352 61062
rect 54300 60998 54352 61004
rect 52380 60846 52500 60874
rect 52472 60790 52500 60846
rect 52460 60784 52512 60790
rect 52460 60726 52512 60732
rect 53104 60512 53156 60518
rect 53104 60454 53156 60460
rect 53116 59634 53144 60454
rect 53748 60172 53800 60178
rect 53748 60114 53800 60120
rect 53104 59628 53156 59634
rect 53104 59570 53156 59576
rect 52920 57996 52972 58002
rect 52920 57938 52972 57944
rect 52460 56976 52512 56982
rect 52460 56918 52512 56924
rect 52472 56166 52500 56918
rect 52460 56160 52512 56166
rect 52460 56102 52512 56108
rect 51908 49088 51960 49094
rect 51908 49030 51960 49036
rect 51920 12918 51948 49030
rect 52000 38004 52052 38010
rect 52000 37946 52052 37952
rect 51908 12912 51960 12918
rect 51908 12854 51960 12860
rect 52012 10606 52040 37946
rect 52828 36100 52880 36106
rect 52828 36042 52880 36048
rect 52472 11218 52776 11234
rect 52460 11212 52788 11218
rect 52512 11206 52736 11212
rect 52460 11154 52512 11160
rect 52736 11154 52788 11160
rect 52840 11150 52868 36042
rect 52932 35894 52960 57938
rect 53656 36780 53708 36786
rect 53656 36722 53708 36728
rect 53472 36168 53524 36174
rect 53472 36110 53524 36116
rect 52932 35866 53144 35894
rect 52828 11144 52880 11150
rect 53012 11144 53064 11150
rect 52828 11086 52880 11092
rect 53010 11112 53012 11121
rect 53064 11112 53066 11121
rect 52000 10600 52052 10606
rect 52000 10542 52052 10548
rect 51814 10296 51870 10305
rect 51814 10231 51870 10240
rect 52644 8628 52696 8634
rect 52644 8570 52696 8576
rect 52000 4616 52052 4622
rect 52000 4558 52052 4564
rect 51724 4140 51776 4146
rect 51724 4082 51776 4088
rect 51540 3936 51592 3942
rect 51540 3878 51592 3884
rect 51552 3602 51580 3878
rect 52012 3738 52040 4558
rect 52460 4208 52512 4214
rect 52460 4150 52512 4156
rect 52000 3732 52052 3738
rect 52000 3674 52052 3680
rect 51540 3596 51592 3602
rect 51540 3538 51592 3544
rect 52000 3528 52052 3534
rect 52000 3470 52052 3476
rect 51632 3460 51684 3466
rect 51632 3402 51684 3408
rect 51644 800 51672 3402
rect 51816 3392 51868 3398
rect 51816 3334 51868 3340
rect 51828 3194 51856 3334
rect 51816 3188 51868 3194
rect 51816 3130 51868 3136
rect 52012 2774 52040 3470
rect 51920 2746 52040 2774
rect 51920 800 51948 2746
rect 52184 2372 52236 2378
rect 52184 2314 52236 2320
rect 52196 800 52224 2314
rect 52472 800 52500 4150
rect 52656 3738 52684 8570
rect 52840 4593 52868 11086
rect 53116 11082 53144 35866
rect 53010 11047 53066 11056
rect 53104 11076 53156 11082
rect 53104 11018 53156 11024
rect 53288 10736 53340 10742
rect 53288 10678 53340 10684
rect 53196 5228 53248 5234
rect 53196 5170 53248 5176
rect 52826 4584 52882 4593
rect 52826 4519 52882 4528
rect 53104 4208 53156 4214
rect 53104 4150 53156 4156
rect 52644 3732 52696 3738
rect 52644 3674 52696 3680
rect 52736 3460 52788 3466
rect 52736 3402 52788 3408
rect 52748 800 52776 3402
rect 53116 2394 53144 4150
rect 53208 4146 53236 5170
rect 53300 4146 53328 10678
rect 53484 4282 53512 36110
rect 53668 36106 53696 36722
rect 53760 36174 53788 60114
rect 54312 43450 54340 60998
rect 54680 60722 54708 63294
rect 55310 63294 55536 63322
rect 55310 63200 55366 63294
rect 55402 61568 55458 61577
rect 55402 61503 55458 61512
rect 55416 60722 55444 61503
rect 55508 61198 55536 63294
rect 56046 63200 56102 64000
rect 56782 63322 56838 64000
rect 56782 63294 56916 63322
rect 56782 63200 56838 63294
rect 56060 61198 56088 63200
rect 56414 62656 56470 62665
rect 56414 62591 56470 62600
rect 56138 62112 56194 62121
rect 56138 62047 56194 62056
rect 55496 61192 55548 61198
rect 55496 61134 55548 61140
rect 56048 61192 56100 61198
rect 56048 61134 56100 61140
rect 56152 60722 56180 62047
rect 54668 60716 54720 60722
rect 54668 60658 54720 60664
rect 55404 60716 55456 60722
rect 55404 60658 55456 60664
rect 56140 60716 56192 60722
rect 56140 60658 56192 60664
rect 54852 60512 54904 60518
rect 54852 60454 54904 60460
rect 55588 60512 55640 60518
rect 55588 60454 55640 60460
rect 56324 60512 56376 60518
rect 56324 60454 56376 60460
rect 54576 49156 54628 49162
rect 54576 49098 54628 49104
rect 54300 43444 54352 43450
rect 54300 43386 54352 43392
rect 54024 37732 54076 37738
rect 54024 37674 54076 37680
rect 54036 36378 54064 37674
rect 54588 36718 54616 49098
rect 54864 46374 54892 60454
rect 55600 59430 55628 60454
rect 56232 60240 56284 60246
rect 56232 60182 56284 60188
rect 56244 59770 56272 60182
rect 56232 59764 56284 59770
rect 56232 59706 56284 59712
rect 56336 59498 56364 60454
rect 56428 59702 56456 62591
rect 56506 61024 56562 61033
rect 56506 60959 56562 60968
rect 56520 60110 56548 60959
rect 56888 60722 56916 63294
rect 57518 63200 57574 64000
rect 58254 63322 58310 64000
rect 57992 63294 58310 63322
rect 57532 61198 57560 63200
rect 57520 61192 57572 61198
rect 57520 61134 57572 61140
rect 56876 60716 56928 60722
rect 56876 60658 56928 60664
rect 57060 60512 57112 60518
rect 57060 60454 57112 60460
rect 57242 60480 57298 60489
rect 56508 60104 56560 60110
rect 56508 60046 56560 60052
rect 56600 59968 56652 59974
rect 56600 59910 56652 59916
rect 56416 59696 56468 59702
rect 56416 59638 56468 59644
rect 56324 59492 56376 59498
rect 56324 59434 56376 59440
rect 55588 59424 55640 59430
rect 55588 59366 55640 59372
rect 56508 58336 56560 58342
rect 56508 58278 56560 58284
rect 56520 56914 56548 58278
rect 56508 56908 56560 56914
rect 56508 56850 56560 56856
rect 54852 46368 54904 46374
rect 54852 46310 54904 46316
rect 56612 36786 56640 59910
rect 57072 44946 57100 60454
rect 57242 60415 57298 60424
rect 57256 60110 57284 60415
rect 57992 60110 58020 63294
rect 58254 63200 58310 63294
rect 58990 63200 59046 64000
rect 58348 61124 58400 61130
rect 58348 61066 58400 61072
rect 58072 60716 58124 60722
rect 58072 60658 58124 60664
rect 57244 60104 57296 60110
rect 57244 60046 57296 60052
rect 57980 60104 58032 60110
rect 57980 60046 58032 60052
rect 58084 59945 58112 60658
rect 58256 60308 58308 60314
rect 58256 60250 58308 60256
rect 58070 59936 58126 59945
rect 58070 59871 58126 59880
rect 58268 59770 58296 60250
rect 58256 59764 58308 59770
rect 58256 59706 58308 59712
rect 58164 59628 58216 59634
rect 58164 59570 58216 59576
rect 57152 59424 57204 59430
rect 58176 59401 58204 59570
rect 57152 59366 57204 59372
rect 58162 59392 58218 59401
rect 57164 59022 57192 59366
rect 58162 59327 58218 59336
rect 58360 59158 58388 61066
rect 58440 60036 58492 60042
rect 58440 59978 58492 59984
rect 58348 59152 58400 59158
rect 58348 59094 58400 59100
rect 57152 59016 57204 59022
rect 57152 58958 57204 58964
rect 57888 59016 57940 59022
rect 57888 58958 57940 58964
rect 57336 58880 57388 58886
rect 57336 58822 57388 58828
rect 57348 58682 57376 58822
rect 57336 58676 57388 58682
rect 57336 58618 57388 58624
rect 57900 58313 57928 58958
rect 58162 58848 58218 58857
rect 58162 58783 58218 58792
rect 58176 58614 58204 58783
rect 58164 58608 58216 58614
rect 58164 58550 58216 58556
rect 57886 58304 57942 58313
rect 57886 58239 57942 58248
rect 57980 57860 58032 57866
rect 57980 57802 58032 57808
rect 57992 57769 58020 57802
rect 57978 57760 58034 57769
rect 57978 57695 58034 57704
rect 57886 57216 57942 57225
rect 57886 57151 57942 57160
rect 57900 56846 57928 57151
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 58072 56772 58124 56778
rect 58072 56714 58124 56720
rect 58084 53145 58112 56714
rect 58162 56672 58218 56681
rect 58162 56607 58218 56616
rect 58176 56438 58204 56607
rect 58164 56432 58216 56438
rect 58164 56374 58216 56380
rect 58346 56128 58402 56137
rect 58346 56063 58402 56072
rect 58360 55962 58388 56063
rect 58348 55956 58400 55962
rect 58348 55898 58400 55904
rect 58348 54664 58400 54670
rect 58348 54606 58400 54612
rect 58360 54505 58388 54606
rect 58346 54496 58402 54505
rect 58346 54431 58402 54440
rect 58070 53136 58126 53145
rect 58070 53071 58126 53080
rect 58348 52896 58400 52902
rect 58346 52864 58348 52873
rect 58400 52864 58402 52873
rect 58346 52799 58402 52808
rect 58348 51400 58400 51406
rect 58348 51342 58400 51348
rect 58360 51241 58388 51342
rect 58346 51232 58402 51241
rect 58346 51167 58402 51176
rect 57888 50176 57940 50182
rect 57888 50118 57940 50124
rect 57900 49609 57928 50118
rect 57886 49600 57942 49609
rect 57886 49535 57942 49544
rect 57980 49156 58032 49162
rect 57980 49098 58032 49104
rect 57992 49065 58020 49098
rect 57978 49056 58034 49065
rect 57978 48991 58034 49000
rect 57244 48068 57296 48074
rect 57244 48010 57296 48016
rect 57980 48068 58032 48074
rect 57980 48010 58032 48016
rect 57256 47977 57284 48010
rect 57242 47968 57298 47977
rect 57242 47903 57298 47912
rect 57992 47433 58020 48010
rect 58072 48000 58124 48006
rect 58072 47942 58124 47948
rect 58084 47802 58112 47942
rect 58072 47796 58124 47802
rect 58072 47738 58124 47744
rect 57978 47424 58034 47433
rect 57978 47359 58034 47368
rect 57520 47048 57572 47054
rect 57520 46990 57572 46996
rect 57060 44940 57112 44946
rect 57060 44882 57112 44888
rect 57244 44804 57296 44810
rect 57244 44746 57296 44752
rect 57256 44713 57284 44746
rect 57242 44704 57298 44713
rect 57242 44639 57298 44648
rect 57060 42628 57112 42634
rect 57060 42570 57112 42576
rect 57072 42537 57100 42570
rect 57152 42560 57204 42566
rect 57058 42528 57114 42537
rect 57152 42502 57204 42508
rect 57058 42463 57114 42472
rect 56968 40520 57020 40526
rect 56968 40462 57020 40468
rect 56980 40361 57008 40462
rect 56966 40352 57022 40361
rect 56966 40287 57022 40296
rect 57060 39364 57112 39370
rect 57060 39306 57112 39312
rect 57072 39273 57100 39306
rect 57058 39264 57114 39273
rect 57058 39199 57114 39208
rect 56600 36780 56652 36786
rect 56600 36722 56652 36728
rect 54576 36712 54628 36718
rect 54576 36654 54628 36660
rect 54024 36372 54076 36378
rect 54024 36314 54076 36320
rect 54588 36174 54616 36654
rect 55128 36644 55180 36650
rect 55128 36586 55180 36592
rect 53748 36168 53800 36174
rect 53748 36110 53800 36116
rect 54576 36168 54628 36174
rect 54576 36110 54628 36116
rect 53656 36100 53708 36106
rect 53656 36042 53708 36048
rect 55140 33266 55168 36586
rect 57164 33930 57192 42502
rect 57244 41540 57296 41546
rect 57244 41482 57296 41488
rect 57256 41449 57284 41482
rect 57242 41440 57298 41449
rect 57242 41375 57298 41384
rect 57152 33924 57204 33930
rect 57152 33866 57204 33872
rect 55140 33238 55352 33266
rect 53840 32428 53892 32434
rect 53840 32370 53892 32376
rect 53472 4276 53524 4282
rect 53472 4218 53524 4224
rect 53196 4140 53248 4146
rect 53196 4082 53248 4088
rect 53288 4140 53340 4146
rect 53288 4082 53340 4088
rect 53378 4040 53434 4049
rect 53378 3975 53434 3984
rect 53392 2990 53420 3975
rect 53472 3392 53524 3398
rect 53472 3334 53524 3340
rect 53656 3392 53708 3398
rect 53656 3334 53708 3340
rect 53380 2984 53432 2990
rect 53380 2926 53432 2932
rect 53024 2366 53144 2394
rect 53288 2372 53340 2378
rect 53024 800 53052 2366
rect 53288 2314 53340 2320
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 53116 1902 53144 2246
rect 53104 1896 53156 1902
rect 53104 1838 53156 1844
rect 53300 800 53328 2314
rect 53484 1766 53512 3334
rect 53668 3126 53696 3334
rect 53852 3194 53880 32370
rect 54760 28416 54812 28422
rect 54760 28358 54812 28364
rect 54024 24200 54076 24206
rect 54024 24142 54076 24148
rect 53932 7336 53984 7342
rect 53932 7278 53984 7284
rect 53944 5846 53972 7278
rect 53932 5840 53984 5846
rect 53932 5782 53984 5788
rect 53932 4548 53984 4554
rect 53932 4490 53984 4496
rect 53944 3466 53972 4490
rect 53932 3460 53984 3466
rect 53932 3402 53984 3408
rect 53840 3188 53892 3194
rect 53840 3130 53892 3136
rect 53656 3120 53708 3126
rect 53656 3062 53708 3068
rect 53564 3052 53616 3058
rect 53564 2994 53616 3000
rect 53840 3052 53892 3058
rect 53840 2994 53892 3000
rect 53472 1760 53524 1766
rect 53472 1702 53524 1708
rect 53576 800 53604 2994
rect 53852 800 53880 2994
rect 54036 2650 54064 24142
rect 54208 11280 54260 11286
rect 54208 11222 54260 11228
rect 54220 4826 54248 11222
rect 54484 11212 54536 11218
rect 54484 11154 54536 11160
rect 54208 4820 54260 4826
rect 54208 4762 54260 4768
rect 54116 4140 54168 4146
rect 54116 4082 54168 4088
rect 54024 2644 54076 2650
rect 54024 2586 54076 2592
rect 54128 800 54156 4082
rect 54300 4072 54352 4078
rect 54300 4014 54352 4020
rect 54312 2774 54340 4014
rect 54312 2746 54432 2774
rect 54404 800 54432 2746
rect 28632 740 28684 746
rect 28632 682 28684 688
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54114 0 54170 800
rect 54390 0 54446 800
rect 54496 105 54524 11154
rect 54772 3194 54800 28358
rect 55220 24132 55272 24138
rect 55220 24074 55272 24080
rect 55232 7546 55260 24074
rect 55220 7540 55272 7546
rect 55220 7482 55272 7488
rect 55218 6216 55274 6225
rect 55218 6151 55220 6160
rect 55272 6151 55274 6160
rect 55220 6122 55272 6128
rect 55324 4010 55352 33238
rect 57060 32836 57112 32842
rect 57060 32778 57112 32784
rect 57072 32745 57100 32778
rect 57152 32768 57204 32774
rect 57058 32736 57114 32745
rect 57152 32710 57204 32716
rect 57058 32671 57114 32680
rect 57164 31210 57192 32710
rect 57152 31204 57204 31210
rect 57152 31146 57204 31152
rect 57060 29572 57112 29578
rect 57060 29514 57112 29520
rect 57072 29481 57100 29514
rect 57058 29472 57114 29481
rect 57058 29407 57114 29416
rect 55680 26920 55732 26926
rect 55680 26862 55732 26868
rect 55404 9512 55456 9518
rect 55404 9454 55456 9460
rect 55416 8945 55444 9454
rect 55402 8936 55458 8945
rect 55402 8871 55458 8880
rect 55404 7540 55456 7546
rect 55404 7482 55456 7488
rect 55312 4004 55364 4010
rect 55312 3946 55364 3952
rect 54760 3188 54812 3194
rect 54760 3130 54812 3136
rect 54944 3052 54996 3058
rect 54944 2994 54996 3000
rect 54668 2440 54720 2446
rect 54668 2382 54720 2388
rect 54680 800 54708 2382
rect 54956 800 54984 2994
rect 55416 2514 55444 7482
rect 55692 3126 55720 26862
rect 57060 26308 57112 26314
rect 57060 26250 57112 26256
rect 57072 26217 57100 26250
rect 57058 26208 57114 26217
rect 57058 26143 57114 26152
rect 55864 22024 55916 22030
rect 55864 21966 55916 21972
rect 55876 15026 55904 21966
rect 57060 16516 57112 16522
rect 57060 16458 57112 16464
rect 57072 16425 57100 16458
rect 57058 16416 57114 16425
rect 57058 16351 57114 16360
rect 56508 15496 56560 15502
rect 56508 15438 56560 15444
rect 55864 15020 55916 15026
rect 55864 14962 55916 14968
rect 56520 14618 56548 15438
rect 56508 14612 56560 14618
rect 56508 14554 56560 14560
rect 57244 14068 57296 14074
rect 57244 14010 57296 14016
rect 57060 13252 57112 13258
rect 57060 13194 57112 13200
rect 57072 13161 57100 13194
rect 57058 13152 57114 13161
rect 57058 13087 57114 13096
rect 56876 10804 56928 10810
rect 56876 10746 56928 10752
rect 56888 10130 56916 10746
rect 57256 10674 57284 14010
rect 57532 13394 57560 46990
rect 57888 46912 57940 46918
rect 57888 46854 57940 46860
rect 57900 46345 57928 46854
rect 57886 46336 57942 46345
rect 57886 46271 57942 46280
rect 57980 45892 58032 45898
rect 57980 45834 58032 45840
rect 57992 45801 58020 45834
rect 57978 45792 58034 45801
rect 57978 45727 58034 45736
rect 57888 44804 57940 44810
rect 57888 44746 57940 44752
rect 57900 44169 57928 44746
rect 58256 44736 58308 44742
rect 58256 44678 58308 44684
rect 57886 44160 57942 44169
rect 57886 44095 57942 44104
rect 58164 43716 58216 43722
rect 58164 43658 58216 43664
rect 58176 43081 58204 43658
rect 58162 43072 58218 43081
rect 58162 43007 58218 43016
rect 57980 42628 58032 42634
rect 57980 42570 58032 42576
rect 57992 41993 58020 42570
rect 57978 41984 58034 41993
rect 57978 41919 58034 41928
rect 57888 41540 57940 41546
rect 57888 41482 57940 41488
rect 57900 40905 57928 41482
rect 57886 40896 57942 40905
rect 57886 40831 57942 40840
rect 57796 40520 57848 40526
rect 57796 40462 57848 40468
rect 57808 34746 57836 40462
rect 57888 40384 57940 40390
rect 57888 40326 57940 40332
rect 57900 39817 57928 40326
rect 57886 39808 57942 39817
rect 57886 39743 57942 39752
rect 57980 39364 58032 39370
rect 57980 39306 58032 39312
rect 57992 38729 58020 39306
rect 58072 39296 58124 39302
rect 58072 39238 58124 39244
rect 58084 39098 58112 39238
rect 58072 39092 58124 39098
rect 58072 39034 58124 39040
rect 57978 38720 58034 38729
rect 57978 38655 58034 38664
rect 58164 38276 58216 38282
rect 58164 38218 58216 38224
rect 58176 38185 58204 38218
rect 58162 38176 58218 38185
rect 58162 38111 58218 38120
rect 58268 38010 58296 44678
rect 58256 38004 58308 38010
rect 58256 37946 58308 37952
rect 58072 37868 58124 37874
rect 58072 37810 58124 37816
rect 58084 37641 58112 37810
rect 58256 37664 58308 37670
rect 58070 37632 58126 37641
rect 58256 37606 58308 37612
rect 58070 37567 58126 37576
rect 58164 37188 58216 37194
rect 58164 37130 58216 37136
rect 58176 36553 58204 37130
rect 58162 36544 58218 36553
rect 58162 36479 58218 36488
rect 57980 36100 58032 36106
rect 57980 36042 58032 36048
rect 57992 36009 58020 36042
rect 57978 36000 58034 36009
rect 57978 35935 58034 35944
rect 58164 35012 58216 35018
rect 58164 34954 58216 34960
rect 58176 34921 58204 34954
rect 58162 34912 58218 34921
rect 58162 34847 58218 34856
rect 57796 34740 57848 34746
rect 57796 34682 57848 34688
rect 57980 34740 58032 34746
rect 57980 34682 58032 34688
rect 57888 34604 57940 34610
rect 57888 34546 57940 34552
rect 57900 34377 57928 34546
rect 57886 34368 57942 34377
rect 57886 34303 57942 34312
rect 57704 32904 57756 32910
rect 57704 32846 57756 32852
rect 57612 23112 57664 23118
rect 57612 23054 57664 23060
rect 57624 14958 57652 23054
rect 57716 18426 57744 32846
rect 57796 31884 57848 31890
rect 57796 31826 57848 31832
rect 57808 31657 57836 31826
rect 57794 31648 57850 31657
rect 57794 31583 57850 31592
rect 57796 29640 57848 29646
rect 57796 29582 57848 29588
rect 57704 18420 57756 18426
rect 57704 18362 57756 18368
rect 57808 15978 57836 29582
rect 57992 20398 58020 34682
rect 58162 33280 58218 33289
rect 58162 33215 58218 33224
rect 58176 32978 58204 33215
rect 58164 32972 58216 32978
rect 58164 32914 58216 32920
rect 58072 31340 58124 31346
rect 58072 31282 58124 31288
rect 58084 31113 58112 31282
rect 58070 31104 58126 31113
rect 58070 31039 58126 31048
rect 58162 30016 58218 30025
rect 58162 29951 58218 29960
rect 58176 29714 58204 29951
rect 58164 29708 58216 29714
rect 58164 29650 58216 29656
rect 58164 28484 58216 28490
rect 58164 28426 58216 28432
rect 58176 28393 58204 28426
rect 58162 28384 58218 28393
rect 58162 28319 58218 28328
rect 58072 28076 58124 28082
rect 58072 28018 58124 28024
rect 58084 27849 58112 28018
rect 58070 27840 58126 27849
rect 58070 27775 58126 27784
rect 58162 26752 58218 26761
rect 58162 26687 58218 26696
rect 58176 26450 58204 26687
rect 58164 26444 58216 26450
rect 58164 26386 58216 26392
rect 58164 25220 58216 25226
rect 58164 25162 58216 25168
rect 58176 25129 58204 25162
rect 58162 25120 58218 25129
rect 58162 25055 58218 25064
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 58084 24585 58112 24754
rect 58070 24576 58126 24585
rect 58070 24511 58126 24520
rect 58162 23488 58218 23497
rect 58162 23423 58218 23432
rect 58176 23186 58204 23423
rect 58164 23180 58216 23186
rect 58164 23122 58216 23128
rect 58070 22944 58126 22953
rect 58070 22879 58126 22888
rect 58084 22642 58112 22879
rect 58072 22636 58124 22642
rect 58072 22578 58124 22584
rect 58164 21956 58216 21962
rect 58164 21898 58216 21904
rect 58176 21865 58204 21898
rect 58162 21856 58218 21865
rect 58162 21791 58218 21800
rect 58072 21548 58124 21554
rect 58072 21490 58124 21496
rect 58084 21321 58112 21490
rect 58070 21312 58126 21321
rect 58070 21247 58126 21256
rect 57980 20392 58032 20398
rect 57980 20334 58032 20340
rect 58162 20224 58218 20233
rect 58162 20159 58218 20168
rect 58176 19922 58204 20159
rect 58164 19916 58216 19922
rect 58164 19858 58216 19864
rect 58070 19680 58126 19689
rect 58070 19615 58126 19624
rect 58084 19378 58112 19615
rect 58268 19530 58296 37606
rect 58348 36100 58400 36106
rect 58348 36042 58400 36048
rect 58360 20806 58388 36042
rect 58452 31958 58480 59978
rect 59004 59430 59032 63200
rect 58992 59424 59044 59430
rect 58992 59366 59044 59372
rect 58532 58948 58584 58954
rect 58532 58890 58584 58896
rect 58440 31952 58492 31958
rect 58440 31894 58492 31900
rect 58544 26897 58572 58890
rect 58624 42628 58676 42634
rect 58624 42570 58676 42576
rect 58636 35222 58664 42570
rect 58624 35216 58676 35222
rect 58624 35158 58676 35164
rect 58530 26888 58586 26897
rect 58530 26823 58586 26832
rect 58348 20800 58400 20806
rect 58348 20742 58400 20748
rect 58176 19502 58296 19530
rect 58176 19446 58204 19502
rect 58164 19440 58216 19446
rect 58164 19382 58216 19388
rect 58072 19372 58124 19378
rect 58072 19314 58124 19320
rect 58256 19236 58308 19242
rect 58256 19178 58308 19184
rect 57886 18864 57942 18873
rect 57886 18799 57942 18808
rect 57900 18766 57928 18799
rect 57888 18760 57940 18766
rect 57888 18702 57940 18708
rect 58164 18692 58216 18698
rect 58164 18634 58216 18640
rect 58176 18601 58204 18634
rect 58162 18592 58218 18601
rect 58162 18527 58218 18536
rect 58268 18426 58296 19178
rect 58256 18420 58308 18426
rect 58256 18362 58308 18368
rect 58072 18284 58124 18290
rect 58072 18226 58124 18232
rect 58084 18057 58112 18226
rect 58070 18048 58126 18057
rect 58070 17983 58126 17992
rect 58162 16960 58218 16969
rect 58162 16895 58218 16904
rect 58176 16590 58204 16895
rect 58164 16584 58216 16590
rect 58164 16526 58216 16532
rect 57796 15972 57848 15978
rect 57796 15914 57848 15920
rect 58164 15428 58216 15434
rect 58164 15370 58216 15376
rect 58176 15337 58204 15370
rect 58162 15328 58218 15337
rect 58162 15263 58218 15272
rect 57612 14952 57664 14958
rect 57612 14894 57664 14900
rect 57978 14784 58034 14793
rect 57978 14719 58034 14728
rect 57992 14414 58020 14719
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 58070 14376 58126 14385
rect 58070 14311 58126 14320
rect 58084 14278 58112 14311
rect 58072 14272 58124 14278
rect 58072 14214 58124 14220
rect 58162 13696 58218 13705
rect 58162 13631 58218 13640
rect 58176 13394 58204 13631
rect 57520 13388 57572 13394
rect 57520 13330 57572 13336
rect 58164 13388 58216 13394
rect 58164 13330 58216 13336
rect 57520 12232 57572 12238
rect 57520 12174 57572 12180
rect 57532 10674 57560 12174
rect 58164 12164 58216 12170
rect 58164 12106 58216 12112
rect 58176 12073 58204 12106
rect 58162 12064 58218 12073
rect 58162 11999 58218 12008
rect 58072 11756 58124 11762
rect 58072 11698 58124 11704
rect 58084 11529 58112 11698
rect 58070 11520 58126 11529
rect 58070 11455 58126 11464
rect 57888 11008 57940 11014
rect 57888 10950 57940 10956
rect 57244 10668 57296 10674
rect 57244 10610 57296 10616
rect 57520 10668 57572 10674
rect 57520 10610 57572 10616
rect 56876 10124 56928 10130
rect 56876 10066 56928 10072
rect 56784 9988 56836 9994
rect 56784 9930 56836 9936
rect 56692 9580 56744 9586
rect 56692 9522 56744 9528
rect 56600 8832 56652 8838
rect 56600 8774 56652 8780
rect 56612 7818 56640 8774
rect 56140 7812 56192 7818
rect 56140 7754 56192 7760
rect 56600 7812 56652 7818
rect 56600 7754 56652 7760
rect 56152 7478 56180 7754
rect 56140 7472 56192 7478
rect 56140 7414 56192 7420
rect 56048 6724 56100 6730
rect 56048 6666 56100 6672
rect 56060 6322 56088 6666
rect 56152 6458 56180 7414
rect 56140 6452 56192 6458
rect 56140 6394 56192 6400
rect 56048 6316 56100 6322
rect 56048 6258 56100 6264
rect 56152 6254 56180 6394
rect 56704 6322 56732 9522
rect 56796 9450 56824 9930
rect 56784 9444 56836 9450
rect 56784 9386 56836 9392
rect 56888 7954 56916 10066
rect 57256 9058 57284 10610
rect 57336 10464 57388 10470
rect 57336 10406 57388 10412
rect 57348 9722 57376 10406
rect 57532 10266 57560 10610
rect 57900 10441 57928 10950
rect 58256 10532 58308 10538
rect 58256 10474 58308 10480
rect 57886 10432 57942 10441
rect 57886 10367 57942 10376
rect 57520 10260 57572 10266
rect 57520 10202 57572 10208
rect 58070 9888 58126 9897
rect 58070 9823 58126 9832
rect 57336 9716 57388 9722
rect 57336 9658 57388 9664
rect 58084 9586 58112 9823
rect 58268 9722 58296 10474
rect 58256 9716 58308 9722
rect 58256 9658 58308 9664
rect 58072 9580 58124 9586
rect 58072 9522 58124 9528
rect 57164 9030 57284 9058
rect 57164 8974 57192 9030
rect 57152 8968 57204 8974
rect 57152 8910 57204 8916
rect 57152 8492 57204 8498
rect 57152 8434 57204 8440
rect 57164 8265 57192 8434
rect 57150 8256 57206 8265
rect 57150 8191 57206 8200
rect 56876 7948 56928 7954
rect 56876 7890 56928 7896
rect 56784 7200 56836 7206
rect 56784 7142 56836 7148
rect 56796 6798 56824 7142
rect 56888 6866 56916 7890
rect 57256 7546 57284 9030
rect 58256 8968 58308 8974
rect 58256 8910 58308 8916
rect 58164 8900 58216 8906
rect 58164 8842 58216 8848
rect 58176 8809 58204 8842
rect 58162 8800 58218 8809
rect 58162 8735 58218 8744
rect 58268 8090 58296 8910
rect 58256 8084 58308 8090
rect 58256 8026 58308 8032
rect 57244 7540 57296 7546
rect 57244 7482 57296 7488
rect 57256 7426 57284 7482
rect 57164 7398 57284 7426
rect 58256 7404 58308 7410
rect 56876 6860 56928 6866
rect 56876 6802 56928 6808
rect 56784 6792 56836 6798
rect 56784 6734 56836 6740
rect 56692 6316 56744 6322
rect 56692 6258 56744 6264
rect 56140 6248 56192 6254
rect 56140 6190 56192 6196
rect 55772 6112 55824 6118
rect 55772 6054 55824 6060
rect 55784 5710 55812 6054
rect 55772 5704 55824 5710
rect 55772 5646 55824 5652
rect 56704 4826 56732 6258
rect 56888 5778 56916 6802
rect 56876 5772 56928 5778
rect 56876 5714 56928 5720
rect 56692 4820 56744 4826
rect 56692 4762 56744 4768
rect 56888 3602 56916 5714
rect 57164 5234 57192 7398
rect 58256 7346 58308 7352
rect 57336 7336 57388 7342
rect 57336 7278 57388 7284
rect 57348 7177 57376 7278
rect 57334 7168 57390 7177
rect 57334 7103 57390 7112
rect 58268 7002 58296 7346
rect 58256 6996 58308 7002
rect 58256 6938 58308 6944
rect 58070 6624 58126 6633
rect 58070 6559 58126 6568
rect 57244 6384 57296 6390
rect 57244 6326 57296 6332
rect 57256 5370 57284 6326
rect 58084 6322 58112 6559
rect 58072 6316 58124 6322
rect 58072 6258 58124 6264
rect 58348 5636 58400 5642
rect 58348 5578 58400 5584
rect 57336 5568 57388 5574
rect 57336 5510 57388 5516
rect 58162 5536 58218 5545
rect 57244 5364 57296 5370
rect 57244 5306 57296 5312
rect 57348 5234 57376 5510
rect 58162 5471 58218 5480
rect 57152 5228 57204 5234
rect 57152 5170 57204 5176
rect 57336 5228 57388 5234
rect 57336 5170 57388 5176
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 57348 4622 57376 5170
rect 58084 5001 58112 5170
rect 58070 4992 58126 5001
rect 58070 4927 58126 4936
rect 58176 4690 58204 5471
rect 58164 4684 58216 4690
rect 58164 4626 58216 4632
rect 57336 4616 57388 4622
rect 57336 4558 57388 4564
rect 57244 4548 57296 4554
rect 57244 4490 57296 4496
rect 56876 3596 56928 3602
rect 56876 3538 56928 3544
rect 56232 3460 56284 3466
rect 56232 3402 56284 3408
rect 55680 3120 55732 3126
rect 55680 3062 55732 3068
rect 55772 2984 55824 2990
rect 55772 2926 55824 2932
rect 55404 2508 55456 2514
rect 55404 2450 55456 2456
rect 55496 2304 55548 2310
rect 55496 2246 55548 2252
rect 55508 800 55536 2246
rect 55784 800 55812 2926
rect 56244 2281 56272 3402
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56230 2272 56286 2281
rect 56230 2207 56286 2216
rect 56428 1834 56456 2382
rect 56416 1828 56468 1834
rect 56416 1770 56468 1776
rect 57256 1737 57284 4490
rect 57888 4208 57940 4214
rect 57888 4150 57940 4156
rect 57900 3913 57928 4150
rect 58360 4146 58388 5578
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 58348 4140 58400 4146
rect 58348 4082 58400 4088
rect 57886 3904 57942 3913
rect 57886 3839 57942 3848
rect 57886 2816 57942 2825
rect 57886 2751 57942 2760
rect 57900 2446 57928 2751
rect 57992 2650 58020 4082
rect 58256 4072 58308 4078
rect 58256 4014 58308 4020
rect 58162 3360 58218 3369
rect 58162 3295 58218 3304
rect 58176 3126 58204 3295
rect 58268 3194 58296 4014
rect 58256 3188 58308 3194
rect 58256 3130 58308 3136
rect 58164 3120 58216 3126
rect 58164 3062 58216 3068
rect 57980 2644 58032 2650
rect 57980 2586 58032 2592
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 57242 1728 57298 1737
rect 57242 1663 57298 1672
rect 56506 1184 56562 1193
rect 56506 1119 56562 1128
rect 54482 96 54538 105
rect 54482 31 54538 40
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56520 105 56548 1119
rect 56506 96 56562 105
rect 56506 31 56562 40
<< via2 >>
rect 1674 61784 1730 61840
rect 1582 60424 1638 60480
rect 1674 59744 1730 59800
rect 2778 61140 2780 61160
rect 2780 61140 2832 61160
rect 2832 61140 2834 61160
rect 2778 61104 2834 61140
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 1582 59064 1638 59120
rect 1582 58384 1638 58440
rect 1582 57704 1638 57760
rect 1582 57024 1638 57080
rect 1582 56344 1638 56400
rect 1674 55684 1730 55720
rect 1674 55664 1676 55684
rect 1676 55664 1728 55684
rect 1728 55664 1730 55684
rect 1582 54984 1638 55040
rect 1674 54304 1730 54360
rect 1582 53624 1638 53680
rect 1674 52944 1730 53000
rect 1582 52264 1638 52320
rect 1674 51584 1730 51640
rect 1674 50904 1730 50960
rect 1674 50244 1730 50280
rect 1674 50224 1676 50244
rect 1676 50224 1728 50244
rect 1728 50224 1730 50244
rect 1582 49544 1638 49600
rect 1674 48864 1730 48920
rect 1674 48184 1730 48240
rect 1674 47504 1730 47560
rect 1858 52556 1914 52592
rect 1858 52536 1860 52556
rect 1860 52536 1912 52556
rect 1912 52536 1914 52556
rect 1858 47504 1914 47560
rect 1582 46824 1638 46880
rect 1582 46144 1638 46200
rect 1674 45464 1730 45520
rect 1582 44820 1584 44840
rect 1584 44820 1636 44840
rect 1636 44820 1638 44840
rect 1582 44784 1638 44820
rect 1674 44104 1730 44160
rect 1674 43424 1730 43480
rect 1582 42744 1638 42800
rect 1674 42064 1730 42120
rect 1674 41384 1730 41440
rect 1674 40704 1730 40760
rect 1674 40024 1730 40080
rect 1674 39364 1730 39400
rect 1674 39344 1676 39364
rect 1676 39344 1728 39364
rect 1728 39344 1730 39364
rect 1674 38664 1730 38720
rect 1674 37984 1730 38040
rect 1674 37304 1730 37360
rect 1674 35944 1730 36000
rect 1674 35264 1730 35320
rect 1674 34584 1730 34640
rect 1674 33924 1730 33960
rect 1674 33904 1676 33924
rect 1676 33904 1728 33924
rect 1728 33904 1730 33924
rect 1674 33224 1730 33280
rect 1674 32544 1730 32600
rect 1674 31864 1730 31920
rect 1674 31184 1730 31240
rect 1674 30504 1730 30560
rect 1766 29824 1822 29880
rect 1858 29144 1914 29200
rect 1858 28484 1914 28520
rect 1858 28464 1860 28484
rect 1860 28464 1912 28484
rect 1912 28464 1914 28484
rect 1766 27784 1822 27840
rect 1858 27104 1914 27160
rect 1766 26424 1822 26480
rect 1766 25780 1768 25800
rect 1768 25780 1820 25800
rect 1820 25780 1822 25800
rect 1766 25744 1822 25780
rect 1858 25064 1914 25120
rect 1766 24384 1822 24440
rect 1858 23704 1914 23760
rect 1858 23044 1914 23080
rect 1858 23024 1860 23044
rect 1860 23024 1912 23044
rect 1912 23024 1914 23044
rect 1766 22344 1822 22400
rect 1858 21664 1914 21720
rect 1766 20984 1822 21040
rect 1766 20340 1768 20360
rect 1768 20340 1820 20360
rect 1820 20340 1822 20360
rect 1766 20304 1822 20340
rect 1858 19624 1914 19680
rect 1858 18944 1914 19000
rect 1858 18264 1914 18320
rect 1858 17604 1914 17640
rect 1858 17584 1860 17604
rect 1860 17584 1912 17604
rect 1912 17584 1914 17604
rect 1766 16904 1822 16960
rect 1858 16224 1914 16280
rect 1766 15544 1822 15600
rect 1766 14900 1768 14920
rect 1768 14900 1820 14920
rect 1820 14900 1822 14920
rect 1766 14864 1822 14900
rect 1858 14184 1914 14240
rect 1766 13504 1822 13560
rect 1858 12824 1914 12880
rect 1858 12180 1860 12200
rect 1860 12180 1912 12200
rect 1912 12180 1914 12200
rect 1858 12144 1914 12180
rect 1766 11464 1822 11520
rect 1858 10784 1914 10840
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4802 51720 4858 51776
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 3054 36624 3110 36680
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 6826 59628 6882 59664
rect 6826 59608 6828 59628
rect 6828 59608 6880 59628
rect 6880 59608 6882 59628
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 2410 14900 2412 14920
rect 2412 14900 2464 14920
rect 2464 14900 2466 14920
rect 2410 14864 2466 14900
rect 2410 14320 2466 14376
rect 1766 10104 1822 10160
rect 1582 9580 1638 9616
rect 1582 9560 1584 9580
rect 1584 9560 1636 9580
rect 1636 9560 1638 9580
rect 1766 9460 1768 9480
rect 1768 9460 1820 9480
rect 1820 9460 1822 9480
rect 1766 9424 1822 9460
rect 1858 8744 1914 8800
rect 1766 8064 1822 8120
rect 1858 7384 1914 7440
rect 1858 6724 1914 6760
rect 1858 6704 1860 6724
rect 1860 6704 1912 6724
rect 1912 6704 1914 6724
rect 1766 6024 1822 6080
rect 1858 5344 1914 5400
rect 1766 4664 1822 4720
rect 1766 4020 1768 4040
rect 1768 4020 1820 4040
rect 1820 4020 1822 4040
rect 1766 3984 1822 4020
rect 1858 3304 1914 3360
rect 1766 2624 1822 2680
rect 1858 1944 1914 2000
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3146 5072 3202 5128
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3698 856 3754 912
rect 5170 3168 5226 3224
rect 6734 2896 6790 2952
rect 7470 3304 7526 3360
rect 8666 4800 8722 4856
rect 12898 60696 12954 60752
rect 15198 50224 15254 50280
rect 10506 26832 10562 26888
rect 10230 13776 10286 13832
rect 9402 7248 9458 7304
rect 8758 2488 8814 2544
rect 9310 4936 9366 4992
rect 9586 4820 9642 4856
rect 9586 4800 9588 4820
rect 9588 4800 9640 4820
rect 9640 4800 9642 4820
rect 9218 4256 9274 4312
rect 9126 4120 9182 4176
rect 8942 1944 8998 2000
rect 9494 3304 9550 3360
rect 9862 2916 9918 2952
rect 9862 2896 9864 2916
rect 9864 2896 9916 2916
rect 9916 2896 9918 2916
rect 10322 7792 10378 7848
rect 10598 12824 10654 12880
rect 11242 15020 11298 15056
rect 11242 15000 11244 15020
rect 11244 15000 11296 15020
rect 11296 15000 11298 15020
rect 11794 14728 11850 14784
rect 11426 13504 11482 13560
rect 10782 12280 10838 12336
rect 10690 11872 10746 11928
rect 10598 4528 10654 4584
rect 11886 12688 11942 12744
rect 11702 12144 11758 12200
rect 11610 11328 11666 11384
rect 13266 14184 13322 14240
rect 12346 13232 12402 13288
rect 12622 12980 12678 13016
rect 12622 12960 12624 12980
rect 12624 12960 12676 12980
rect 12676 12960 12678 12980
rect 12438 12688 12494 12744
rect 11886 8200 11942 8256
rect 11518 3168 11574 3224
rect 12990 13132 12992 13152
rect 12992 13132 13044 13152
rect 13044 13132 13046 13152
rect 12990 13096 13046 13132
rect 13542 13640 13598 13696
rect 13542 13096 13598 13152
rect 12806 12008 12862 12064
rect 12622 10784 12678 10840
rect 12162 5208 12218 5264
rect 12070 3168 12126 3224
rect 12530 3848 12586 3904
rect 12438 3440 12494 3496
rect 12070 2624 12126 2680
rect 11794 2352 11850 2408
rect 12622 2624 12678 2680
rect 13082 7792 13138 7848
rect 12990 4120 13046 4176
rect 13358 11192 13414 11248
rect 13266 11056 13322 11112
rect 14186 11736 14242 11792
rect 13634 9016 13690 9072
rect 14462 17992 14518 18048
rect 14370 13640 14426 13696
rect 14554 10920 14610 10976
rect 14922 15408 14978 15464
rect 15014 15000 15070 15056
rect 14738 12960 14794 13016
rect 14830 12688 14886 12744
rect 14462 9288 14518 9344
rect 13726 7656 13782 7712
rect 13910 7112 13966 7168
rect 13266 2624 13322 2680
rect 14002 6976 14058 7032
rect 14094 5228 14150 5264
rect 14094 5208 14096 5228
rect 14096 5208 14148 5228
rect 14148 5208 14150 5228
rect 15106 12280 15162 12336
rect 15014 11872 15070 11928
rect 15474 12416 15530 12472
rect 15198 11600 15254 11656
rect 15658 12980 15714 13016
rect 15842 14220 15844 14240
rect 15844 14220 15896 14240
rect 15896 14220 15898 14240
rect 15842 14184 15898 14220
rect 15658 12960 15660 12980
rect 15660 12960 15712 12980
rect 15712 12960 15714 12980
rect 15658 12552 15714 12608
rect 15106 10104 15162 10160
rect 14738 7656 14794 7712
rect 14278 2760 14334 2816
rect 14554 1400 14610 1456
rect 14922 6432 14978 6488
rect 15750 12280 15806 12336
rect 16026 13404 16028 13424
rect 16028 13404 16080 13424
rect 16080 13404 16082 13424
rect 16026 13368 16082 13404
rect 15934 11464 15990 11520
rect 15750 10512 15806 10568
rect 16762 17720 16818 17776
rect 16210 13640 16266 13696
rect 16118 12280 16174 12336
rect 15842 9696 15898 9752
rect 16118 9832 16174 9888
rect 15474 5616 15530 5672
rect 15290 3576 15346 3632
rect 15106 992 15162 1048
rect 15658 7384 15714 7440
rect 16210 8900 16266 8936
rect 16210 8880 16212 8900
rect 16212 8880 16264 8900
rect 16264 8880 16266 8900
rect 16302 8744 16358 8800
rect 15658 1128 15714 1184
rect 15842 2896 15898 2952
rect 16854 12008 16910 12064
rect 17222 24248 17278 24304
rect 17130 17856 17186 17912
rect 18510 59372 18512 59392
rect 18512 59372 18564 59392
rect 18564 59372 18566 59392
rect 18510 59336 18566 59372
rect 17682 50360 17738 50416
rect 17958 36624 18014 36680
rect 17590 19080 17646 19136
rect 17406 17176 17462 17232
rect 16946 11328 17002 11384
rect 16670 11056 16726 11112
rect 17038 11192 17094 11248
rect 16854 10240 16910 10296
rect 16946 10104 17002 10160
rect 17406 13504 17462 13560
rect 17498 12824 17554 12880
rect 17314 11192 17370 11248
rect 17590 11464 17646 11520
rect 17406 11056 17462 11112
rect 17222 10920 17278 10976
rect 16946 9424 17002 9480
rect 16578 3068 16580 3088
rect 16580 3068 16632 3088
rect 16632 3068 16634 3088
rect 16578 3032 16634 3068
rect 17222 6704 17278 6760
rect 17498 10104 17554 10160
rect 17406 9288 17462 9344
rect 17406 9172 17462 9208
rect 17406 9152 17408 9172
rect 17408 9152 17460 9172
rect 17460 9152 17462 9172
rect 18050 19796 18052 19816
rect 18052 19796 18104 19816
rect 18104 19796 18106 19816
rect 18050 19760 18106 19796
rect 17866 13912 17922 13968
rect 18050 13796 18106 13832
rect 18050 13776 18052 13796
rect 18052 13776 18104 13796
rect 18104 13776 18106 13796
rect 18050 12280 18106 12336
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19154 36644 19210 36680
rect 19154 36624 19156 36644
rect 19156 36624 19208 36644
rect 19208 36624 19210 36644
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19522 37868 19578 37904
rect 19522 37848 19524 37868
rect 19524 37848 19576 37868
rect 19576 37848 19578 37868
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19706 35012 19762 35048
rect 19706 34992 19708 35012
rect 19708 34992 19760 35012
rect 19760 34992 19762 35012
rect 21178 60052 21180 60072
rect 21180 60052 21232 60072
rect 21232 60052 21234 60072
rect 21178 60016 21234 60052
rect 21086 58792 21142 58848
rect 20166 34992 20222 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 20074 30640 20130 30696
rect 19430 24112 19486 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 18234 12844 18290 12880
rect 18234 12824 18236 12844
rect 18236 12824 18288 12844
rect 18288 12824 18290 12844
rect 18326 10920 18382 10976
rect 18602 12724 18604 12744
rect 18604 12724 18656 12744
rect 18656 12724 18658 12744
rect 18602 12688 18658 12724
rect 18970 19080 19026 19136
rect 18878 16904 18934 16960
rect 18602 10784 18658 10840
rect 17958 8880 18014 8936
rect 17682 8472 17738 8528
rect 17498 6160 17554 6216
rect 17590 5888 17646 5944
rect 17590 5752 17646 5808
rect 16946 4156 16948 4176
rect 16948 4156 17000 4176
rect 17000 4156 17002 4176
rect 16946 4120 17002 4156
rect 17130 3984 17186 4040
rect 17130 2352 17186 2408
rect 17222 1536 17278 1592
rect 17498 1264 17554 1320
rect 18694 9832 18750 9888
rect 18418 9696 18474 9752
rect 18510 9288 18566 9344
rect 18234 8336 18290 8392
rect 18418 7928 18474 7984
rect 18418 6840 18474 6896
rect 18326 6568 18382 6624
rect 18234 6296 18290 6352
rect 18142 5208 18198 5264
rect 18418 4936 18474 4992
rect 17958 2352 18014 2408
rect 18050 1672 18106 1728
rect 18878 11348 18934 11384
rect 18878 11328 18880 11348
rect 18880 11328 18932 11348
rect 18932 11328 18934 11348
rect 19246 14184 19302 14240
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19982 15544 20038 15600
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18878 9696 18934 9752
rect 18786 9152 18842 9208
rect 18602 8064 18658 8120
rect 18786 7656 18842 7712
rect 18786 5072 18842 5128
rect 18510 3984 18566 4040
rect 18510 3712 18566 3768
rect 18602 3168 18658 3224
rect 18694 2624 18750 2680
rect 19062 8880 19118 8936
rect 18970 8744 19026 8800
rect 19062 8336 19118 8392
rect 19246 10648 19302 10704
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19430 9968 19486 10024
rect 19798 10004 19800 10024
rect 19800 10004 19852 10024
rect 19852 10004 19854 10024
rect 19798 9968 19854 10004
rect 19338 8336 19394 8392
rect 19154 8064 19210 8120
rect 19154 7656 19210 7712
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19798 9424 19854 9480
rect 19706 8900 19762 8936
rect 19706 8880 19708 8900
rect 19708 8880 19760 8900
rect 19760 8880 19762 8900
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19982 8608 20038 8664
rect 19982 8336 20038 8392
rect 19798 7928 19854 7984
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7520 19486 7576
rect 19982 7520 20038 7576
rect 19062 6568 19118 6624
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19338 6452 19394 6488
rect 19338 6432 19340 6452
rect 19340 6432 19392 6452
rect 19392 6432 19394 6452
rect 19246 6316 19302 6352
rect 19246 6296 19248 6316
rect 19248 6296 19300 6316
rect 19300 6296 19302 6316
rect 20534 15272 20590 15328
rect 20350 14456 20406 14512
rect 20350 11736 20406 11792
rect 20350 10920 20406 10976
rect 20442 10784 20498 10840
rect 20810 13132 20812 13152
rect 20812 13132 20864 13152
rect 20864 13132 20866 13152
rect 20810 13096 20866 13132
rect 20442 9832 20498 9888
rect 20810 11736 20866 11792
rect 20810 11464 20866 11520
rect 20810 10920 20866 10976
rect 22098 59336 22154 59392
rect 22650 59744 22706 59800
rect 22558 59472 22614 59528
rect 21454 22072 21510 22128
rect 20718 9696 20774 9752
rect 20626 9424 20682 9480
rect 20626 9152 20682 9208
rect 20258 8336 20314 8392
rect 20258 7948 20314 7984
rect 20258 7928 20260 7948
rect 20260 7928 20312 7948
rect 20312 7928 20314 7948
rect 20258 6840 20314 6896
rect 20442 8744 20498 8800
rect 20534 8064 20590 8120
rect 21086 8608 21142 8664
rect 20810 7828 20812 7848
rect 20812 7828 20864 7848
rect 20864 7828 20866 7848
rect 20810 7792 20866 7828
rect 20902 7540 20958 7576
rect 20902 7520 20904 7540
rect 20904 7520 20956 7540
rect 20956 7520 20958 7540
rect 20718 6840 20774 6896
rect 20442 6296 20498 6352
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19338 5072 19394 5128
rect 19982 4392 20038 4448
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20166 5480 20222 5536
rect 19430 4020 19432 4040
rect 19432 4020 19484 4040
rect 19484 4020 19486 4040
rect 19430 3984 19486 4020
rect 19614 3712 19670 3768
rect 20258 5344 20314 5400
rect 20350 5072 20406 5128
rect 20442 4256 20498 4312
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19430 3168 19486 3224
rect 20074 3168 20130 3224
rect 19798 2896 19854 2952
rect 19982 2932 19984 2952
rect 19984 2932 20036 2952
rect 20036 2932 20038 2952
rect 19982 2896 20038 2932
rect 20074 2760 20130 2816
rect 19982 2488 20038 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20718 4256 20774 4312
rect 20626 3712 20682 3768
rect 20902 3340 20904 3360
rect 20904 3340 20956 3360
rect 20956 3340 20958 3360
rect 20902 3304 20958 3340
rect 20718 2760 20774 2816
rect 20902 2760 20958 2816
rect 20626 2624 20682 2680
rect 20442 1808 20498 1864
rect 20902 2624 20958 2680
rect 21270 11056 21326 11112
rect 22098 38528 22154 38584
rect 22098 34604 22154 34640
rect 22098 34584 22100 34604
rect 22100 34584 22152 34604
rect 22152 34584 22154 34604
rect 23202 38528 23258 38584
rect 22190 34448 22246 34504
rect 22650 35944 22706 36000
rect 23018 34992 23074 35048
rect 22558 28464 22614 28520
rect 21638 19488 21694 19544
rect 21730 17584 21786 17640
rect 21546 12960 21602 13016
rect 21638 12824 21694 12880
rect 22098 19760 22154 19816
rect 22006 19292 22062 19348
rect 22190 19488 22246 19544
rect 22742 22616 22798 22672
rect 22374 19080 22430 19136
rect 22006 15408 22062 15464
rect 22098 14864 22154 14920
rect 21546 10920 21602 10976
rect 21454 7520 21510 7576
rect 21270 3576 21326 3632
rect 21546 7112 21602 7168
rect 21546 4256 21602 4312
rect 21914 11464 21970 11520
rect 21914 11076 21970 11112
rect 21914 11056 21916 11076
rect 21916 11056 21968 11076
rect 21968 11056 21970 11076
rect 21914 10648 21970 10704
rect 21914 7928 21970 7984
rect 22190 11092 22192 11112
rect 22192 11092 22244 11112
rect 22244 11092 22246 11112
rect 22190 11056 22246 11092
rect 22190 10668 22246 10704
rect 22190 10648 22192 10668
rect 22192 10648 22244 10668
rect 22244 10648 22246 10668
rect 22374 10648 22430 10704
rect 22098 8780 22100 8800
rect 22100 8780 22152 8800
rect 22152 8780 22154 8800
rect 22098 8744 22154 8780
rect 22006 7520 22062 7576
rect 22742 19488 22798 19544
rect 22650 19352 22706 19408
rect 22742 17992 22798 18048
rect 22374 8744 22430 8800
rect 22282 7656 22338 7712
rect 22098 6704 22154 6760
rect 21914 6060 21916 6080
rect 21916 6060 21968 6080
rect 21968 6060 21970 6080
rect 21914 6024 21970 6060
rect 22098 6024 22154 6080
rect 21914 3848 21970 3904
rect 21822 3712 21878 3768
rect 22558 8336 22614 8392
rect 22558 8064 22614 8120
rect 22466 6840 22522 6896
rect 22466 6432 22522 6488
rect 22834 13232 22890 13288
rect 22926 9288 22982 9344
rect 23110 7792 23166 7848
rect 22466 4392 22522 4448
rect 22190 3460 22246 3496
rect 22190 3440 22192 3460
rect 22192 3440 22244 3460
rect 22244 3440 22246 3460
rect 22834 5888 22890 5944
rect 22834 5228 22890 5264
rect 22834 5208 22836 5228
rect 22836 5208 22888 5228
rect 22888 5208 22890 5228
rect 22098 3032 22154 3088
rect 22006 2624 22062 2680
rect 22742 3984 22798 4040
rect 23018 6704 23074 6760
rect 23478 34992 23534 35048
rect 23846 59880 23902 59936
rect 23846 34584 23902 34640
rect 23570 14864 23626 14920
rect 23570 12416 23626 12472
rect 23294 8744 23350 8800
rect 23294 8336 23350 8392
rect 23478 6840 23534 6896
rect 23294 6316 23350 6352
rect 23294 6296 23296 6316
rect 23296 6296 23348 6316
rect 23348 6296 23350 6316
rect 23110 4256 23166 4312
rect 23386 6024 23442 6080
rect 23938 30096 23994 30152
rect 23846 23432 23902 23488
rect 23754 19216 23810 19272
rect 23754 13504 23810 13560
rect 23846 11192 23902 11248
rect 23662 10920 23718 10976
rect 23662 10004 23664 10024
rect 23664 10004 23716 10024
rect 23716 10004 23718 10024
rect 23662 9968 23718 10004
rect 23662 9288 23718 9344
rect 23754 8608 23810 8664
rect 23754 8492 23810 8528
rect 23754 8472 23756 8492
rect 23756 8472 23808 8492
rect 23808 8472 23810 8492
rect 23662 5480 23718 5536
rect 24674 59880 24730 59936
rect 25870 59744 25926 59800
rect 25778 59492 25834 59528
rect 25778 59472 25780 59492
rect 25780 59472 25832 59492
rect 25832 59472 25834 59492
rect 24582 41540 24638 41576
rect 24582 41520 24584 41540
rect 24584 41520 24636 41540
rect 24636 41520 24638 41540
rect 25134 30252 25190 30288
rect 25134 30232 25136 30252
rect 25136 30232 25188 30252
rect 25188 30232 25190 30252
rect 25594 37848 25650 37904
rect 26054 37848 26110 37904
rect 27250 59880 27306 59936
rect 26882 58792 26938 58848
rect 26422 47640 26478 47696
rect 25686 30232 25742 30288
rect 26330 30116 26386 30152
rect 26330 30096 26332 30116
rect 26332 30096 26384 30116
rect 26384 30096 26386 30116
rect 24766 19896 24822 19952
rect 24582 19780 24638 19816
rect 24582 19760 24584 19780
rect 24584 19760 24636 19780
rect 24636 19760 24638 19780
rect 24766 19352 24822 19408
rect 24306 18264 24362 18320
rect 24582 17756 24584 17776
rect 24584 17756 24636 17776
rect 24636 17756 24638 17776
rect 24582 17720 24638 17756
rect 24030 14320 24086 14376
rect 24122 14048 24178 14104
rect 24030 12844 24086 12880
rect 24030 12824 24032 12844
rect 24032 12824 24084 12844
rect 24084 12824 24086 12844
rect 24030 10684 24032 10704
rect 24032 10684 24084 10704
rect 24084 10684 24086 10704
rect 24030 10648 24086 10684
rect 24122 10240 24178 10296
rect 24582 12008 24638 12064
rect 24214 8744 24270 8800
rect 24398 8472 24454 8528
rect 23478 5072 23534 5128
rect 23110 3440 23166 3496
rect 22926 3052 22982 3088
rect 22926 3032 22928 3052
rect 22928 3032 22980 3052
rect 22980 3032 22982 3052
rect 23110 2760 23166 2816
rect 23018 2624 23074 2680
rect 23938 3168 23994 3224
rect 25226 19896 25282 19952
rect 24674 9968 24730 10024
rect 24674 9832 24730 9888
rect 25134 7948 25190 7984
rect 25686 19760 25742 19816
rect 25502 14356 25504 14376
rect 25504 14356 25556 14376
rect 25556 14356 25558 14376
rect 25502 14320 25558 14356
rect 25778 14456 25834 14512
rect 25594 11464 25650 11520
rect 25134 7928 25136 7948
rect 25136 7928 25188 7948
rect 25188 7928 25190 7948
rect 24490 5888 24546 5944
rect 24306 5480 24362 5536
rect 24950 6568 25006 6624
rect 24122 3168 24178 3224
rect 24398 3848 24454 3904
rect 24398 3576 24454 3632
rect 24950 3576 25006 3632
rect 25134 3576 25190 3632
rect 25778 12008 25834 12064
rect 26054 18164 26056 18184
rect 26056 18164 26108 18184
rect 26108 18164 26110 18184
rect 26054 18128 26110 18164
rect 26882 24792 26938 24848
rect 26422 17720 26478 17776
rect 26514 13096 26570 13152
rect 25962 10920 26018 10976
rect 25778 9424 25834 9480
rect 26054 9152 26110 9208
rect 26422 9696 26478 9752
rect 25778 7284 25780 7304
rect 25780 7284 25832 7304
rect 25832 7284 25834 7304
rect 25778 7248 25834 7284
rect 25594 5480 25650 5536
rect 26698 10784 26754 10840
rect 26698 9968 26754 10024
rect 26422 4120 26478 4176
rect 25502 3712 25558 3768
rect 25778 3596 25834 3632
rect 25778 3576 25780 3596
rect 25780 3576 25832 3596
rect 25832 3576 25834 3596
rect 25134 1808 25190 1864
rect 24674 720 24730 776
rect 25410 1536 25466 1592
rect 25686 1400 25742 1456
rect 27158 26968 27214 27024
rect 27434 21936 27490 21992
rect 28538 60016 28594 60072
rect 28998 60052 29000 60072
rect 29000 60052 29052 60072
rect 29052 60052 29054 60072
rect 28998 60016 29054 60052
rect 29734 60308 29790 60344
rect 29734 60288 29736 60308
rect 29736 60288 29788 60308
rect 29788 60288 29790 60308
rect 29642 60172 29698 60208
rect 29642 60152 29644 60172
rect 29644 60152 29696 60172
rect 29696 60152 29698 60172
rect 28446 22752 28502 22808
rect 26974 12552 27030 12608
rect 26974 8628 27030 8664
rect 27526 18300 27528 18320
rect 27528 18300 27580 18320
rect 27580 18300 27582 18320
rect 27526 18264 27582 18300
rect 27434 18164 27436 18184
rect 27436 18164 27488 18184
rect 27488 18164 27490 18184
rect 27434 18128 27490 18164
rect 27618 16360 27674 16416
rect 27894 17740 27950 17776
rect 27894 17720 27896 17740
rect 27896 17720 27948 17740
rect 27948 17720 27950 17740
rect 27250 13776 27306 13832
rect 27526 13132 27528 13152
rect 27528 13132 27580 13152
rect 27580 13132 27582 13152
rect 27526 13096 27582 13132
rect 27158 12552 27214 12608
rect 27802 12552 27858 12608
rect 26974 8608 26976 8628
rect 26976 8608 27028 8628
rect 27028 8608 27030 8628
rect 27434 9016 27490 9072
rect 27618 10240 27674 10296
rect 27526 7112 27582 7168
rect 27526 6840 27582 6896
rect 27342 5908 27398 5944
rect 27342 5888 27344 5908
rect 27344 5888 27396 5908
rect 27396 5888 27398 5908
rect 27894 9696 27950 9752
rect 29274 19080 29330 19136
rect 28998 17720 29054 17776
rect 28538 14320 28594 14376
rect 28998 15544 29054 15600
rect 27986 7692 27988 7712
rect 27988 7692 28040 7712
rect 28040 7692 28042 7712
rect 27986 7656 28042 7692
rect 27802 5480 27858 5536
rect 27066 1672 27122 1728
rect 27986 4256 28042 4312
rect 28170 4528 28226 4584
rect 28354 4664 28410 4720
rect 28814 10376 28870 10432
rect 28906 9424 28962 9480
rect 28906 8336 28962 8392
rect 28906 5344 28962 5400
rect 28630 4700 28632 4720
rect 28632 4700 28684 4720
rect 28684 4700 28686 4720
rect 28630 4664 28686 4700
rect 28814 4800 28870 4856
rect 28630 3848 28686 3904
rect 27802 992 27858 1048
rect 28538 3032 28594 3088
rect 28998 3576 29054 3632
rect 29458 9152 29514 9208
rect 29458 9016 29514 9072
rect 29182 6332 29184 6352
rect 29184 6332 29236 6352
rect 29236 6332 29238 6352
rect 29182 6296 29238 6332
rect 31574 61124 31630 61160
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 31574 61104 31576 61124
rect 31576 61104 31628 61124
rect 31628 61104 31630 61124
rect 30010 60308 30066 60344
rect 30010 60288 30012 60308
rect 30012 60288 30064 60308
rect 30064 60288 30066 60308
rect 30010 60152 30066 60208
rect 30194 60052 30196 60072
rect 30196 60052 30248 60072
rect 30248 60052 30250 60072
rect 30194 60016 30250 60052
rect 30286 18672 30342 18728
rect 30010 15952 30066 16008
rect 29734 13096 29790 13152
rect 30194 15000 30250 15056
rect 30102 13504 30158 13560
rect 30010 13096 30066 13152
rect 30378 15680 30434 15736
rect 30102 12144 30158 12200
rect 29918 11464 29974 11520
rect 29918 11056 29974 11112
rect 29642 9016 29698 9072
rect 29366 4528 29422 4584
rect 29090 1264 29146 1320
rect 29458 4120 29514 4176
rect 29458 4020 29460 4040
rect 29460 4020 29512 4040
rect 29512 4020 29514 4040
rect 29458 3984 29514 4020
rect 30010 10784 30066 10840
rect 29918 9288 29974 9344
rect 29734 6840 29790 6896
rect 30102 9696 30158 9752
rect 30102 9288 30158 9344
rect 30102 8200 30158 8256
rect 31022 26288 31078 26344
rect 31206 17076 31208 17096
rect 31208 17076 31260 17096
rect 31260 17076 31262 17096
rect 31206 17040 31262 17076
rect 31114 16396 31116 16416
rect 31116 16396 31168 16416
rect 31168 16396 31170 16416
rect 31114 16360 31170 16396
rect 30746 14728 30802 14784
rect 30286 7656 30342 7712
rect 30102 6160 30158 6216
rect 30010 5888 30066 5944
rect 30286 5752 30342 5808
rect 30010 3984 30066 4040
rect 30746 9152 30802 9208
rect 32126 16224 32182 16280
rect 32218 15136 32274 15192
rect 31298 10804 31354 10840
rect 31298 10784 31300 10804
rect 31300 10784 31352 10804
rect 31352 10784 31354 10804
rect 30654 5888 30710 5944
rect 30654 5516 30656 5536
rect 30656 5516 30708 5536
rect 30708 5516 30710 5536
rect 30654 5480 30710 5516
rect 30470 4120 30526 4176
rect 30102 2896 30158 2952
rect 31206 9580 31262 9616
rect 31206 9560 31208 9580
rect 31208 9560 31260 9580
rect 31260 9560 31262 9580
rect 31114 7656 31170 7712
rect 31114 6840 31170 6896
rect 31206 6568 31262 6624
rect 31022 6024 31078 6080
rect 31022 5752 31078 5808
rect 31850 10124 31906 10160
rect 31850 10104 31852 10124
rect 31852 10104 31904 10124
rect 31904 10104 31906 10124
rect 31574 9580 31630 9616
rect 31574 9560 31576 9580
rect 31576 9560 31628 9580
rect 31628 9560 31630 9580
rect 31574 8744 31630 8800
rect 31758 9152 31814 9208
rect 31666 8064 31722 8120
rect 31942 8336 31998 8392
rect 31390 5108 31392 5128
rect 31392 5108 31444 5128
rect 31444 5108 31446 5128
rect 31390 5072 31446 5108
rect 30562 2488 30618 2544
rect 30286 1944 30342 2000
rect 31666 5480 31722 5536
rect 31850 5480 31906 5536
rect 31850 5344 31906 5400
rect 32402 13232 32458 13288
rect 33322 56652 33324 56672
rect 33324 56652 33376 56672
rect 33376 56652 33378 56672
rect 33322 56616 33378 56652
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34518 42880 34574 42936
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 32586 13096 32642 13152
rect 32494 12860 32496 12880
rect 32496 12860 32548 12880
rect 32548 12860 32550 12880
rect 32494 12824 32550 12860
rect 33138 12960 33194 13016
rect 33046 12824 33102 12880
rect 32678 12588 32680 12608
rect 32680 12588 32732 12608
rect 32732 12588 32734 12608
rect 32678 12552 32734 12588
rect 32770 12416 32826 12472
rect 32586 10668 32642 10704
rect 32586 10648 32588 10668
rect 32588 10648 32640 10668
rect 32640 10648 32642 10668
rect 32126 8472 32182 8528
rect 32402 7248 32458 7304
rect 32862 11464 32918 11520
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 35530 60016 35586 60072
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 33690 17040 33746 17096
rect 33782 14592 33838 14648
rect 34058 15680 34114 15736
rect 34058 14864 34114 14920
rect 33966 14592 34022 14648
rect 33598 12552 33654 12608
rect 32862 10376 32918 10432
rect 32678 9716 32734 9752
rect 32678 9696 32680 9716
rect 32680 9696 32732 9716
rect 32732 9696 32734 9716
rect 32678 6840 32734 6896
rect 32954 9560 33010 9616
rect 32954 8880 33010 8936
rect 32586 6432 32642 6488
rect 31758 4120 31814 4176
rect 32402 5888 32458 5944
rect 32402 5616 32458 5672
rect 32402 5208 32458 5264
rect 32770 4936 32826 4992
rect 32678 4664 32734 4720
rect 33506 12144 33562 12200
rect 33322 11092 33324 11112
rect 33324 11092 33376 11112
rect 33376 11092 33378 11112
rect 33322 11056 33378 11092
rect 33506 9696 33562 9752
rect 33414 9288 33470 9344
rect 33322 9016 33378 9072
rect 33690 10920 33746 10976
rect 34058 11328 34114 11384
rect 34058 10376 34114 10432
rect 33966 10240 34022 10296
rect 33230 6840 33286 6896
rect 33322 6024 33378 6080
rect 33230 5616 33286 5672
rect 32310 3168 32366 3224
rect 32954 4548 33010 4584
rect 32954 4528 32956 4548
rect 32956 4528 33008 4548
rect 33008 4528 33010 4548
rect 33230 3612 33232 3632
rect 33232 3612 33284 3632
rect 33284 3612 33286 3632
rect 33230 3576 33286 3612
rect 34058 9832 34114 9888
rect 34058 9580 34114 9616
rect 34058 9560 34060 9580
rect 34060 9560 34112 9580
rect 34112 9560 34114 9580
rect 34426 19216 34482 19272
rect 34242 14048 34298 14104
rect 34518 14048 34574 14104
rect 34334 11872 34390 11928
rect 34242 11056 34298 11112
rect 34518 12416 34574 12472
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35070 19508 35126 19544
rect 35070 19488 35072 19508
rect 35072 19488 35124 19508
rect 35124 19488 35126 19508
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34886 18808 34942 18864
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34886 17720 34942 17776
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35806 19488 35862 19544
rect 35714 16652 35770 16688
rect 35714 16632 35716 16652
rect 35716 16632 35768 16652
rect 35768 16632 35770 16652
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35070 15136 35126 15192
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34702 13912 34758 13968
rect 34886 13932 34942 13968
rect 34886 13912 34888 13932
rect 34888 13912 34940 13932
rect 34940 13912 34942 13932
rect 35530 14900 35532 14920
rect 35532 14900 35584 14920
rect 35584 14900 35586 14920
rect 35530 14864 35586 14900
rect 35806 15544 35862 15600
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35438 13640 35494 13696
rect 34978 13096 35034 13152
rect 34702 11464 34758 11520
rect 34610 11328 34666 11384
rect 35530 12824 35586 12880
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34886 12144 34942 12200
rect 35622 12300 35678 12336
rect 35622 12280 35624 12300
rect 35624 12280 35676 12300
rect 35676 12280 35678 12300
rect 36910 42644 36912 42664
rect 36912 42644 36964 42664
rect 36964 42644 36966 42664
rect 36910 42608 36966 42644
rect 36266 18808 36322 18864
rect 35806 13132 35808 13152
rect 35808 13132 35860 13152
rect 35860 13132 35862 13152
rect 35806 13096 35862 13132
rect 35162 11872 35218 11928
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35530 11056 35586 11112
rect 34334 10240 34390 10296
rect 34242 9596 34244 9616
rect 34244 9596 34296 9616
rect 34296 9596 34298 9616
rect 34242 9560 34298 9596
rect 33966 9288 34022 9344
rect 33874 8200 33930 8256
rect 33966 7520 34022 7576
rect 33598 5888 33654 5944
rect 33598 5752 33654 5808
rect 34242 8608 34298 8664
rect 34702 10376 34758 10432
rect 34610 9288 34666 9344
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34794 10240 34850 10296
rect 35254 9832 35310 9888
rect 34978 9560 35034 9616
rect 34794 9288 34850 9344
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34518 8608 34574 8664
rect 34610 8200 34666 8256
rect 34886 8472 34942 8528
rect 35254 8608 35310 8664
rect 35530 10376 35586 10432
rect 35806 11056 35862 11112
rect 36082 11464 36138 11520
rect 36266 11756 36322 11792
rect 36266 11736 36268 11756
rect 36268 11736 36320 11756
rect 36320 11736 36322 11756
rect 36266 11328 36322 11384
rect 36174 11056 36230 11112
rect 35714 10240 35770 10296
rect 35438 9832 35494 9888
rect 35622 9324 35624 9344
rect 35624 9324 35676 9344
rect 35676 9324 35678 9344
rect 35622 9288 35678 9324
rect 35346 8472 35402 8528
rect 34150 7112 34206 7168
rect 33966 5752 34022 5808
rect 33506 4140 33562 4176
rect 33506 4120 33508 4140
rect 33508 4120 33560 4140
rect 33560 4120 33562 4140
rect 33322 856 33378 912
rect 34150 3168 34206 3224
rect 34610 6976 34666 7032
rect 34702 6840 34758 6896
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35254 7404 35310 7440
rect 35254 7384 35256 7404
rect 35256 7384 35308 7404
rect 35308 7384 35310 7404
rect 35806 9580 35862 9616
rect 35806 9560 35808 9580
rect 35808 9560 35860 9580
rect 35860 9560 35862 9580
rect 36082 10920 36138 10976
rect 35990 9832 36046 9888
rect 36174 9832 36230 9888
rect 36082 9424 36138 9480
rect 35990 9288 36046 9344
rect 35346 7112 35402 7168
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35806 8064 35862 8120
rect 36450 12960 36506 13016
rect 36634 15000 36690 15056
rect 36634 14592 36690 14648
rect 36910 15952 36966 16008
rect 36910 14048 36966 14104
rect 36818 13368 36874 13424
rect 36634 11192 36690 11248
rect 36634 10920 36690 10976
rect 36542 9152 36598 9208
rect 36910 9832 36966 9888
rect 35806 7112 35862 7168
rect 34886 6876 34888 6896
rect 34888 6876 34940 6896
rect 34940 6876 34942 6896
rect 34886 6840 34942 6876
rect 35530 6840 35586 6896
rect 34610 6024 34666 6080
rect 34518 5888 34574 5944
rect 34426 4664 34482 4720
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35530 6024 35586 6080
rect 35438 5344 35494 5400
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35530 4684 35586 4720
rect 35530 4664 35532 4684
rect 35532 4664 35584 4684
rect 35584 4664 35586 4684
rect 36358 8200 36414 8256
rect 36358 7248 36414 7304
rect 36174 6568 36230 6624
rect 36174 5616 36230 5672
rect 35898 5108 35900 5128
rect 35900 5108 35952 5128
rect 35952 5108 35954 5128
rect 35898 5072 35954 5108
rect 36542 7112 36598 7168
rect 36266 4800 36322 4856
rect 35898 4120 35954 4176
rect 35438 3304 35494 3360
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35714 3848 35770 3904
rect 35898 3732 35954 3768
rect 36266 4256 36322 4312
rect 35898 3712 35900 3732
rect 35900 3712 35952 3732
rect 35952 3712 35954 3732
rect 36910 8508 36912 8528
rect 36912 8508 36964 8528
rect 36964 8508 36966 8528
rect 36910 8472 36966 8508
rect 37186 16632 37242 16688
rect 37186 13912 37242 13968
rect 37554 16632 37610 16688
rect 38014 20712 38070 20768
rect 37738 15952 37794 16008
rect 37738 15444 37740 15464
rect 37740 15444 37792 15464
rect 37792 15444 37794 15464
rect 37738 15408 37794 15444
rect 37554 14612 37610 14648
rect 37554 14592 37556 14612
rect 37556 14592 37608 14612
rect 37608 14592 37610 14612
rect 37094 13504 37150 13560
rect 37646 13776 37702 13832
rect 37738 13640 37794 13696
rect 37738 13268 37740 13288
rect 37740 13268 37792 13288
rect 37792 13268 37794 13288
rect 37738 13232 37794 13268
rect 37370 11348 37426 11384
rect 37370 11328 37372 11348
rect 37372 11328 37424 11348
rect 37424 11328 37426 11348
rect 37186 9288 37242 9344
rect 37002 6604 37004 6624
rect 37004 6604 37056 6624
rect 37056 6604 37058 6624
rect 37002 6568 37058 6604
rect 37554 12144 37610 12200
rect 37554 10104 37610 10160
rect 38106 17720 38162 17776
rect 38198 13776 38254 13832
rect 38106 10920 38162 10976
rect 38106 10376 38162 10432
rect 37278 8200 37334 8256
rect 36910 6024 36966 6080
rect 36818 5208 36874 5264
rect 36726 3984 36782 4040
rect 36910 3576 36966 3632
rect 38014 9696 38070 9752
rect 37646 6976 37702 7032
rect 37554 6840 37610 6896
rect 37370 6160 37426 6216
rect 36082 1128 36138 1184
rect 38198 8200 38254 8256
rect 38842 15428 38898 15464
rect 38842 15408 38844 15428
rect 38844 15408 38896 15428
rect 38896 15408 38898 15428
rect 38842 15156 38898 15192
rect 38842 15136 38844 15156
rect 38844 15136 38896 15156
rect 38896 15136 38898 15156
rect 38750 15000 38806 15056
rect 38750 14048 38806 14104
rect 38566 12824 38622 12880
rect 38566 11464 38622 11520
rect 38658 10920 38714 10976
rect 38750 10240 38806 10296
rect 38382 9560 38438 9616
rect 38658 9424 38714 9480
rect 38566 8200 38622 8256
rect 38474 7928 38530 7984
rect 38934 9696 38990 9752
rect 38750 7928 38806 7984
rect 38474 7112 38530 7168
rect 37830 4800 37886 4856
rect 38198 6568 38254 6624
rect 37462 3168 37518 3224
rect 38014 3848 38070 3904
rect 38934 8608 38990 8664
rect 38842 7248 38898 7304
rect 39210 17584 39266 17640
rect 39118 14864 39174 14920
rect 39394 14220 39396 14240
rect 39396 14220 39448 14240
rect 39448 14220 39450 14240
rect 39394 14184 39450 14220
rect 39118 7828 39120 7848
rect 39120 7828 39172 7848
rect 39172 7828 39174 7848
rect 39118 7792 39174 7828
rect 39210 7384 39266 7440
rect 39118 7248 39174 7304
rect 38382 4664 38438 4720
rect 39026 3984 39082 4040
rect 39302 3440 39358 3496
rect 39762 59608 39818 59664
rect 39854 18944 39910 19000
rect 40406 57976 40462 58032
rect 42614 59336 42670 59392
rect 42706 57296 42762 57352
rect 40314 15136 40370 15192
rect 39578 9696 39634 9752
rect 40130 14592 40186 14648
rect 40314 13640 40370 13696
rect 40682 19252 40684 19272
rect 40684 19252 40736 19272
rect 40736 19252 40738 19272
rect 40682 19216 40738 19252
rect 40590 19080 40646 19136
rect 40590 15408 40646 15464
rect 40590 14048 40646 14104
rect 39946 12688 40002 12744
rect 40038 12416 40094 12472
rect 40130 12044 40132 12064
rect 40132 12044 40184 12064
rect 40184 12044 40186 12064
rect 40130 12008 40186 12044
rect 40498 12688 40554 12744
rect 41234 19252 41236 19272
rect 41236 19252 41288 19272
rect 41288 19252 41290 19272
rect 41234 19216 41290 19252
rect 41050 14592 41106 14648
rect 41418 14864 41474 14920
rect 41142 13504 41198 13560
rect 39762 9580 39818 9616
rect 39762 9560 39764 9580
rect 39764 9560 39816 9580
rect 39816 9560 39818 9580
rect 39670 9288 39726 9344
rect 39578 9152 39634 9208
rect 39670 8508 39672 8528
rect 39672 8508 39724 8528
rect 39724 8508 39726 8528
rect 39670 8472 39726 8508
rect 39762 8200 39818 8256
rect 39670 6296 39726 6352
rect 40682 11464 40738 11520
rect 40866 11328 40922 11384
rect 40314 9968 40370 10024
rect 40222 9696 40278 9752
rect 40130 9288 40186 9344
rect 40038 7928 40094 7984
rect 41602 13640 41658 13696
rect 41234 12552 41290 12608
rect 40682 10376 40738 10432
rect 40498 8492 40554 8528
rect 40498 8472 40505 8492
rect 40505 8472 40554 8492
rect 40682 8336 40738 8392
rect 40222 2644 40278 2680
rect 40222 2624 40224 2644
rect 40224 2624 40276 2644
rect 40276 2624 40278 2644
rect 40590 3984 40646 4040
rect 40866 8744 40922 8800
rect 40866 8200 40922 8256
rect 41510 12416 41566 12472
rect 41510 10512 41566 10568
rect 41234 8744 41290 8800
rect 41234 7520 41290 7576
rect 42154 13640 42210 13696
rect 42062 12416 42118 12472
rect 41326 2644 41382 2680
rect 41326 2624 41328 2644
rect 41328 2624 41380 2644
rect 41380 2624 41382 2644
rect 42338 14048 42394 14104
rect 42246 7656 42302 7712
rect 42338 5480 42394 5536
rect 41970 3984 42026 4040
rect 42154 3476 42156 3496
rect 42156 3476 42208 3496
rect 42208 3476 42210 3496
rect 42154 3440 42210 3476
rect 41970 3032 42026 3088
rect 42706 15272 42762 15328
rect 42706 14456 42762 14512
rect 43350 14048 43406 14104
rect 43258 12416 43314 12472
rect 42614 10648 42670 10704
rect 42614 9016 42670 9072
rect 43074 11600 43130 11656
rect 42614 3304 42670 3360
rect 42798 2644 42854 2680
rect 42798 2624 42800 2644
rect 42800 2624 42852 2644
rect 42852 2624 42854 2644
rect 43810 14048 43866 14104
rect 43626 11228 43628 11248
rect 43628 11228 43680 11248
rect 43680 11228 43682 11248
rect 43626 11192 43682 11228
rect 44086 13776 44142 13832
rect 44086 11192 44142 11248
rect 44270 9152 44326 9208
rect 43810 6840 43866 6896
rect 43258 4684 43314 4720
rect 43258 4664 43260 4684
rect 43260 4664 43312 4684
rect 43312 4664 43314 4684
rect 43718 4548 43774 4584
rect 43718 4528 43720 4548
rect 43720 4528 43772 4548
rect 43772 4528 43774 4548
rect 42982 4120 43038 4176
rect 43994 5344 44050 5400
rect 43350 3984 43406 4040
rect 43534 3576 43590 3632
rect 43534 2352 43590 2408
rect 44546 7928 44602 7984
rect 44546 4140 44602 4176
rect 44546 4120 44548 4140
rect 44548 4120 44600 4140
rect 44600 4120 44602 4140
rect 44362 3032 44418 3088
rect 44362 2896 44418 2952
rect 45558 4664 45614 4720
rect 44822 2896 44878 2952
rect 45926 9560 45982 9616
rect 46478 15000 46534 15056
rect 46754 11464 46810 11520
rect 46570 3440 46626 3496
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 47766 19388 47768 19408
rect 47768 19388 47820 19408
rect 47820 19388 47822 19408
rect 47766 19352 47822 19388
rect 48226 19508 48282 19544
rect 48226 19488 48228 19508
rect 48228 19488 48280 19508
rect 48280 19488 48282 19508
rect 48134 19080 48190 19136
rect 48226 18708 48228 18728
rect 48228 18708 48280 18728
rect 48280 18708 48282 18728
rect 48226 18672 48282 18708
rect 48686 19488 48742 19544
rect 48594 18828 48650 18864
rect 48594 18808 48596 18828
rect 48596 18808 48648 18828
rect 48648 18808 48650 18828
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 48962 19352 49018 19408
rect 49146 18672 49202 18728
rect 48962 10784 49018 10840
rect 48042 3304 48098 3360
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 49330 3848 49386 3904
rect 49698 8064 49754 8120
rect 49698 3612 49700 3632
rect 49700 3612 49752 3632
rect 49752 3612 49754 3632
rect 49698 3576 49754 3612
rect 49698 3168 49754 3224
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50618 11076 50674 11112
rect 50618 11056 50620 11076
rect 50620 11056 50672 11076
rect 50672 11056 50674 11076
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 51262 6704 51318 6760
rect 53010 11092 53012 11112
rect 53012 11092 53064 11112
rect 53064 11092 53066 11112
rect 51814 10240 51870 10296
rect 53010 11056 53066 11092
rect 52826 4528 52882 4584
rect 55402 61512 55458 61568
rect 56414 62600 56470 62656
rect 56138 62056 56194 62112
rect 56506 60968 56562 61024
rect 57242 60424 57298 60480
rect 58070 59880 58126 59936
rect 58162 59336 58218 59392
rect 58162 58792 58218 58848
rect 57886 58248 57942 58304
rect 57978 57704 58034 57760
rect 57886 57160 57942 57216
rect 58162 56616 58218 56672
rect 58346 56072 58402 56128
rect 58346 54440 58402 54496
rect 58070 53080 58126 53136
rect 58346 52844 58348 52864
rect 58348 52844 58400 52864
rect 58400 52844 58402 52864
rect 58346 52808 58402 52844
rect 58346 51176 58402 51232
rect 57886 49544 57942 49600
rect 57978 49000 58034 49056
rect 57242 47912 57298 47968
rect 57978 47368 58034 47424
rect 57242 44648 57298 44704
rect 57058 42472 57114 42528
rect 56966 40296 57022 40352
rect 57058 39208 57114 39264
rect 57242 41384 57298 41440
rect 53378 3984 53434 4040
rect 55218 6180 55274 6216
rect 55218 6160 55220 6180
rect 55220 6160 55272 6180
rect 55272 6160 55274 6180
rect 57058 32680 57114 32736
rect 57058 29416 57114 29472
rect 55402 8880 55458 8936
rect 57058 26152 57114 26208
rect 57058 16360 57114 16416
rect 57058 13096 57114 13152
rect 57886 46280 57942 46336
rect 57978 45736 58034 45792
rect 57886 44104 57942 44160
rect 58162 43016 58218 43072
rect 57978 41928 58034 41984
rect 57886 40840 57942 40896
rect 57886 39752 57942 39808
rect 57978 38664 58034 38720
rect 58162 38120 58218 38176
rect 58070 37576 58126 37632
rect 58162 36488 58218 36544
rect 57978 35944 58034 36000
rect 58162 34856 58218 34912
rect 57886 34312 57942 34368
rect 57794 31592 57850 31648
rect 58162 33224 58218 33280
rect 58070 31048 58126 31104
rect 58162 29960 58218 30016
rect 58162 28328 58218 28384
rect 58070 27784 58126 27840
rect 58162 26696 58218 26752
rect 58162 25064 58218 25120
rect 58070 24520 58126 24576
rect 58162 23432 58218 23488
rect 58070 22888 58126 22944
rect 58162 21800 58218 21856
rect 58070 21256 58126 21312
rect 58162 20168 58218 20224
rect 58070 19624 58126 19680
rect 58530 26832 58586 26888
rect 57886 18808 57942 18864
rect 58162 18536 58218 18592
rect 58070 17992 58126 18048
rect 58162 16904 58218 16960
rect 58162 15272 58218 15328
rect 57978 14728 58034 14784
rect 58070 14320 58126 14376
rect 58162 13640 58218 13696
rect 58162 12008 58218 12064
rect 58070 11464 58126 11520
rect 57886 10376 57942 10432
rect 58070 9832 58126 9888
rect 57150 8200 57206 8256
rect 58162 8744 58218 8800
rect 57334 7112 57390 7168
rect 58070 6568 58126 6624
rect 58162 5480 58218 5536
rect 58070 4936 58126 4992
rect 56230 2216 56286 2272
rect 57886 3848 57942 3904
rect 57886 2760 57942 2816
rect 58162 3304 58218 3360
rect 57242 1672 57298 1728
rect 56506 1128 56562 1184
rect 54482 40 54538 96
rect 56506 40 56562 96
<< metal3 >>
rect 56409 62658 56475 62661
rect 59200 62658 60000 62688
rect 56409 62656 60000 62658
rect 56409 62600 56414 62656
rect 56470 62600 60000 62656
rect 56409 62598 60000 62600
rect 56409 62595 56475 62598
rect 59200 62568 60000 62598
rect 56133 62114 56199 62117
rect 59200 62114 60000 62144
rect 56133 62112 60000 62114
rect 56133 62056 56138 62112
rect 56194 62056 60000 62112
rect 56133 62054 60000 62056
rect 56133 62051 56199 62054
rect 59200 62024 60000 62054
rect 0 61842 800 61872
rect 1669 61842 1735 61845
rect 0 61840 1735 61842
rect 0 61784 1674 61840
rect 1730 61784 1735 61840
rect 0 61782 1735 61784
rect 0 61752 800 61782
rect 1669 61779 1735 61782
rect 55397 61570 55463 61573
rect 59200 61570 60000 61600
rect 55397 61568 60000 61570
rect 55397 61512 55402 61568
rect 55458 61512 60000 61568
rect 55397 61510 60000 61512
rect 55397 61507 55463 61510
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 59200 61480 60000 61510
rect 34930 61439 35246 61440
rect 0 61162 800 61192
rect 2773 61162 2839 61165
rect 0 61160 2839 61162
rect 0 61104 2778 61160
rect 2834 61104 2839 61160
rect 0 61102 2839 61104
rect 0 61072 800 61102
rect 2773 61099 2839 61102
rect 31569 61162 31635 61165
rect 39246 61162 39252 61164
rect 31569 61160 39252 61162
rect 31569 61104 31574 61160
rect 31630 61104 39252 61160
rect 31569 61102 39252 61104
rect 31569 61099 31635 61102
rect 39246 61100 39252 61102
rect 39316 61100 39322 61164
rect 56501 61026 56567 61029
rect 59200 61026 60000 61056
rect 56501 61024 60000 61026
rect 56501 60968 56506 61024
rect 56562 60968 60000 61024
rect 56501 60966 60000 60968
rect 56501 60963 56567 60966
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 59200 60936 60000 60966
rect 50290 60895 50606 60896
rect 12893 60756 12959 60757
rect 12893 60752 12940 60756
rect 13004 60754 13010 60756
rect 12893 60696 12898 60752
rect 12893 60692 12940 60696
rect 13004 60694 13050 60754
rect 13004 60692 13010 60694
rect 12893 60691 12959 60692
rect 0 60482 800 60512
rect 1577 60482 1643 60485
rect 0 60480 1643 60482
rect 0 60424 1582 60480
rect 1638 60424 1643 60480
rect 0 60422 1643 60424
rect 0 60392 800 60422
rect 1577 60419 1643 60422
rect 57237 60482 57303 60485
rect 59200 60482 60000 60512
rect 57237 60480 60000 60482
rect 57237 60424 57242 60480
rect 57298 60424 60000 60480
rect 57237 60422 60000 60424
rect 57237 60419 57303 60422
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 59200 60392 60000 60422
rect 34930 60351 35246 60352
rect 29729 60346 29795 60349
rect 30005 60346 30071 60349
rect 29729 60344 30071 60346
rect 29729 60288 29734 60344
rect 29790 60288 30010 60344
rect 30066 60288 30071 60344
rect 29729 60286 30071 60288
rect 29729 60283 29795 60286
rect 30005 60283 30071 60286
rect 29637 60210 29703 60213
rect 30005 60210 30071 60213
rect 29637 60208 30071 60210
rect 29637 60152 29642 60208
rect 29698 60152 30010 60208
rect 30066 60152 30071 60208
rect 29637 60150 30071 60152
rect 29637 60147 29703 60150
rect 30005 60147 30071 60150
rect 21173 60074 21239 60077
rect 28533 60074 28599 60077
rect 21173 60072 28599 60074
rect 21173 60016 21178 60072
rect 21234 60016 28538 60072
rect 28594 60016 28599 60072
rect 21173 60014 28599 60016
rect 21173 60011 21239 60014
rect 28533 60011 28599 60014
rect 28993 60074 29059 60077
rect 30189 60074 30255 60077
rect 35525 60074 35591 60077
rect 28993 60072 35591 60074
rect 28993 60016 28998 60072
rect 29054 60016 30194 60072
rect 30250 60016 35530 60072
rect 35586 60016 35591 60072
rect 28993 60014 35591 60016
rect 28993 60011 29059 60014
rect 30189 60011 30255 60014
rect 35525 60011 35591 60014
rect 23841 59938 23907 59941
rect 24669 59938 24735 59941
rect 27245 59938 27311 59941
rect 23841 59936 27311 59938
rect 23841 59880 23846 59936
rect 23902 59880 24674 59936
rect 24730 59880 27250 59936
rect 27306 59880 27311 59936
rect 23841 59878 27311 59880
rect 23841 59875 23907 59878
rect 24669 59875 24735 59878
rect 27245 59875 27311 59878
rect 58065 59938 58131 59941
rect 59200 59938 60000 59968
rect 58065 59936 60000 59938
rect 58065 59880 58070 59936
rect 58126 59880 60000 59936
rect 58065 59878 60000 59880
rect 58065 59875 58131 59878
rect 19570 59872 19886 59873
rect 0 59802 800 59832
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 59200 59848 60000 59878
rect 50290 59807 50606 59808
rect 1669 59802 1735 59805
rect 0 59800 1735 59802
rect 0 59744 1674 59800
rect 1730 59744 1735 59800
rect 0 59742 1735 59744
rect 0 59712 800 59742
rect 1669 59739 1735 59742
rect 22645 59802 22711 59805
rect 25865 59802 25931 59805
rect 22645 59800 25931 59802
rect 22645 59744 22650 59800
rect 22706 59744 25870 59800
rect 25926 59744 25931 59800
rect 22645 59742 25931 59744
rect 22645 59739 22711 59742
rect 25865 59739 25931 59742
rect 6821 59666 6887 59669
rect 39757 59666 39823 59669
rect 6821 59664 39823 59666
rect 6821 59608 6826 59664
rect 6882 59608 39762 59664
rect 39818 59608 39823 59664
rect 6821 59606 39823 59608
rect 6821 59603 6887 59606
rect 39757 59603 39823 59606
rect 22553 59530 22619 59533
rect 25773 59530 25839 59533
rect 22553 59528 25839 59530
rect 22553 59472 22558 59528
rect 22614 59472 25778 59528
rect 25834 59472 25839 59528
rect 22553 59470 25839 59472
rect 22553 59467 22619 59470
rect 25773 59467 25839 59470
rect 18505 59396 18571 59397
rect 18454 59332 18460 59396
rect 18524 59394 18571 59396
rect 22093 59394 22159 59397
rect 23054 59394 23060 59396
rect 18524 59392 18616 59394
rect 18566 59336 18616 59392
rect 18524 59334 18616 59336
rect 22093 59392 23060 59394
rect 22093 59336 22098 59392
rect 22154 59336 23060 59392
rect 22093 59334 23060 59336
rect 18524 59332 18571 59334
rect 18505 59331 18571 59332
rect 22093 59331 22159 59334
rect 23054 59332 23060 59334
rect 23124 59332 23130 59396
rect 42374 59332 42380 59396
rect 42444 59394 42450 59396
rect 42609 59394 42675 59397
rect 42444 59392 42675 59394
rect 42444 59336 42614 59392
rect 42670 59336 42675 59392
rect 42444 59334 42675 59336
rect 42444 59332 42450 59334
rect 42609 59331 42675 59334
rect 58157 59394 58223 59397
rect 59200 59394 60000 59424
rect 58157 59392 60000 59394
rect 58157 59336 58162 59392
rect 58218 59336 60000 59392
rect 58157 59334 60000 59336
rect 58157 59331 58223 59334
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 59200 59304 60000 59334
rect 34930 59263 35246 59264
rect 0 59122 800 59152
rect 1577 59122 1643 59125
rect 0 59120 1643 59122
rect 0 59064 1582 59120
rect 1638 59064 1643 59120
rect 0 59062 1643 59064
rect 0 59032 800 59062
rect 1577 59059 1643 59062
rect 21081 58850 21147 58853
rect 21950 58850 21956 58852
rect 21081 58848 21956 58850
rect 21081 58792 21086 58848
rect 21142 58792 21956 58848
rect 21081 58790 21956 58792
rect 21081 58787 21147 58790
rect 21950 58788 21956 58790
rect 22020 58850 22026 58852
rect 26877 58850 26943 58853
rect 22020 58848 26943 58850
rect 22020 58792 26882 58848
rect 26938 58792 26943 58848
rect 22020 58790 26943 58792
rect 22020 58788 22026 58790
rect 26877 58787 26943 58790
rect 58157 58850 58223 58853
rect 59200 58850 60000 58880
rect 58157 58848 60000 58850
rect 58157 58792 58162 58848
rect 58218 58792 60000 58848
rect 58157 58790 60000 58792
rect 58157 58787 58223 58790
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 59200 58760 60000 58790
rect 50290 58719 50606 58720
rect 0 58442 800 58472
rect 1577 58442 1643 58445
rect 0 58440 1643 58442
rect 0 58384 1582 58440
rect 1638 58384 1643 58440
rect 0 58382 1643 58384
rect 0 58352 800 58382
rect 1577 58379 1643 58382
rect 57881 58306 57947 58309
rect 59200 58306 60000 58336
rect 57881 58304 60000 58306
rect 57881 58248 57886 58304
rect 57942 58248 60000 58304
rect 57881 58246 60000 58248
rect 57881 58243 57947 58246
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 59200 58216 60000 58246
rect 34930 58175 35246 58176
rect 40401 58036 40467 58037
rect 40350 58034 40356 58036
rect 40310 57974 40356 58034
rect 40420 58032 40467 58036
rect 40462 57976 40467 58032
rect 40350 57972 40356 57974
rect 40420 57972 40467 57976
rect 40401 57971 40467 57972
rect 0 57762 800 57792
rect 1577 57762 1643 57765
rect 0 57760 1643 57762
rect 0 57704 1582 57760
rect 1638 57704 1643 57760
rect 0 57702 1643 57704
rect 0 57672 800 57702
rect 1577 57699 1643 57702
rect 57973 57762 58039 57765
rect 59200 57762 60000 57792
rect 57973 57760 60000 57762
rect 57973 57704 57978 57760
rect 58034 57704 60000 57760
rect 57973 57702 60000 57704
rect 57973 57699 58039 57702
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 59200 57672 60000 57702
rect 50290 57631 50606 57632
rect 42701 57354 42767 57357
rect 43478 57354 43484 57356
rect 42701 57352 43484 57354
rect 42701 57296 42706 57352
rect 42762 57296 43484 57352
rect 42701 57294 43484 57296
rect 42701 57291 42767 57294
rect 43478 57292 43484 57294
rect 43548 57292 43554 57356
rect 57881 57218 57947 57221
rect 59200 57218 60000 57248
rect 57881 57216 60000 57218
rect 57881 57160 57886 57216
rect 57942 57160 60000 57216
rect 57881 57158 60000 57160
rect 57881 57155 57947 57158
rect 4210 57152 4526 57153
rect 0 57082 800 57112
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 60000 57158
rect 34930 57087 35246 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 800 57022
rect 1577 57019 1643 57022
rect 33317 56674 33383 56677
rect 33910 56674 33916 56676
rect 33317 56672 33916 56674
rect 33317 56616 33322 56672
rect 33378 56616 33916 56672
rect 33317 56614 33916 56616
rect 33317 56611 33383 56614
rect 33910 56612 33916 56614
rect 33980 56612 33986 56676
rect 58157 56674 58223 56677
rect 59200 56674 60000 56704
rect 58157 56672 60000 56674
rect 58157 56616 58162 56672
rect 58218 56616 60000 56672
rect 58157 56614 60000 56616
rect 58157 56611 58223 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 59200 56584 60000 56614
rect 50290 56543 50606 56544
rect 0 56402 800 56432
rect 1577 56402 1643 56405
rect 0 56400 1643 56402
rect 0 56344 1582 56400
rect 1638 56344 1643 56400
rect 0 56342 1643 56344
rect 0 56312 800 56342
rect 1577 56339 1643 56342
rect 58341 56130 58407 56133
rect 59200 56130 60000 56160
rect 58341 56128 60000 56130
rect 58341 56072 58346 56128
rect 58402 56072 60000 56128
rect 58341 56070 60000 56072
rect 58341 56067 58407 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 59200 56040 60000 56070
rect 34930 55999 35246 56000
rect 0 55722 800 55752
rect 1669 55722 1735 55725
rect 0 55720 1735 55722
rect 0 55664 1674 55720
rect 1730 55664 1735 55720
rect 0 55662 1735 55664
rect 0 55632 800 55662
rect 1669 55659 1735 55662
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 59200 55496 60000 55616
rect 50290 55455 50606 55456
rect 0 55042 800 55072
rect 1577 55042 1643 55045
rect 0 55040 1643 55042
rect 0 54984 1582 55040
rect 1638 54984 1643 55040
rect 0 54982 1643 54984
rect 0 54952 800 54982
rect 1577 54979 1643 54982
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 59200 54952 60000 55072
rect 34930 54911 35246 54912
rect 58341 54498 58407 54501
rect 59200 54498 60000 54528
rect 58341 54496 60000 54498
rect 58341 54440 58346 54496
rect 58402 54440 60000 54496
rect 58341 54438 60000 54440
rect 58341 54435 58407 54438
rect 19570 54432 19886 54433
rect 0 54362 800 54392
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 59200 54408 60000 54438
rect 50290 54367 50606 54368
rect 1669 54362 1735 54365
rect 0 54360 1735 54362
rect 0 54304 1674 54360
rect 1730 54304 1735 54360
rect 0 54302 1735 54304
rect 0 54272 800 54302
rect 1669 54299 1735 54302
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 59200 53864 60000 53984
rect 34930 53823 35246 53824
rect 0 53682 800 53712
rect 1577 53682 1643 53685
rect 0 53680 1643 53682
rect 0 53624 1582 53680
rect 1638 53624 1643 53680
rect 0 53622 1643 53624
rect 0 53592 800 53622
rect 1577 53619 1643 53622
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 59200 53320 60000 53440
rect 50290 53279 50606 53280
rect 36118 53076 36124 53140
rect 36188 53138 36194 53140
rect 58065 53138 58131 53141
rect 36188 53136 58131 53138
rect 36188 53080 58070 53136
rect 58126 53080 58131 53136
rect 36188 53078 58131 53080
rect 36188 53076 36194 53078
rect 58065 53075 58131 53078
rect 0 53002 800 53032
rect 1669 53002 1735 53005
rect 0 53000 1735 53002
rect 0 52944 1674 53000
rect 1730 52944 1735 53000
rect 0 52942 1735 52944
rect 0 52912 800 52942
rect 1669 52939 1735 52942
rect 58341 52866 58407 52869
rect 59200 52866 60000 52896
rect 58341 52864 60000 52866
rect 58341 52808 58346 52864
rect 58402 52808 60000 52864
rect 58341 52806 60000 52808
rect 58341 52803 58407 52806
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 59200 52776 60000 52806
rect 34930 52735 35246 52736
rect 1853 52594 1919 52597
rect 31150 52594 31156 52596
rect 1853 52592 31156 52594
rect 1853 52536 1858 52592
rect 1914 52536 31156 52592
rect 1853 52534 31156 52536
rect 1853 52531 1919 52534
rect 31150 52532 31156 52534
rect 31220 52532 31226 52596
rect 0 52322 800 52352
rect 1577 52322 1643 52325
rect 0 52320 1643 52322
rect 0 52264 1582 52320
rect 1638 52264 1643 52320
rect 0 52262 1643 52264
rect 0 52232 800 52262
rect 1577 52259 1643 52262
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 59200 52232 60000 52352
rect 50290 52191 50606 52192
rect 4797 51778 4863 51781
rect 32806 51778 32812 51780
rect 4797 51776 32812 51778
rect 4797 51720 4802 51776
rect 4858 51720 32812 51776
rect 4797 51718 32812 51720
rect 4797 51715 4863 51718
rect 32806 51716 32812 51718
rect 32876 51716 32882 51780
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51808
rect 34930 51647 35246 51648
rect 1669 51642 1735 51645
rect 0 51640 1735 51642
rect 0 51584 1674 51640
rect 1730 51584 1735 51640
rect 0 51582 1735 51584
rect 0 51552 800 51582
rect 1669 51579 1735 51582
rect 58341 51234 58407 51237
rect 59200 51234 60000 51264
rect 58341 51232 60000 51234
rect 58341 51176 58346 51232
rect 58402 51176 60000 51232
rect 58341 51174 60000 51176
rect 58341 51171 58407 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 59200 51144 60000 51174
rect 50290 51103 50606 51104
rect 0 50962 800 50992
rect 1669 50962 1735 50965
rect 0 50960 1735 50962
rect 0 50904 1674 50960
rect 1730 50904 1735 50960
rect 0 50902 1735 50904
rect 0 50872 800 50902
rect 1669 50899 1735 50902
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 59200 50600 60000 50720
rect 34930 50559 35246 50560
rect 17677 50418 17743 50421
rect 36854 50418 36860 50420
rect 17677 50416 36860 50418
rect 17677 50360 17682 50416
rect 17738 50360 36860 50416
rect 17677 50358 36860 50360
rect 17677 50355 17743 50358
rect 36854 50356 36860 50358
rect 36924 50356 36930 50420
rect 0 50282 800 50312
rect 1669 50282 1735 50285
rect 0 50280 1735 50282
rect 0 50224 1674 50280
rect 1730 50224 1735 50280
rect 0 50222 1735 50224
rect 0 50192 800 50222
rect 1669 50219 1735 50222
rect 15193 50282 15259 50285
rect 38510 50282 38516 50284
rect 15193 50280 38516 50282
rect 15193 50224 15198 50280
rect 15254 50224 38516 50280
rect 15193 50222 38516 50224
rect 15193 50219 15259 50222
rect 38510 50220 38516 50222
rect 38580 50220 38586 50284
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 59200 50056 60000 50176
rect 50290 50015 50606 50016
rect 0 49602 800 49632
rect 1577 49602 1643 49605
rect 0 49600 1643 49602
rect 0 49544 1582 49600
rect 1638 49544 1643 49600
rect 0 49542 1643 49544
rect 0 49512 800 49542
rect 1577 49539 1643 49542
rect 57881 49602 57947 49605
rect 59200 49602 60000 49632
rect 57881 49600 60000 49602
rect 57881 49544 57886 49600
rect 57942 49544 60000 49600
rect 57881 49542 60000 49544
rect 57881 49539 57947 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 59200 49512 60000 49542
rect 34930 49471 35246 49472
rect 57973 49058 58039 49061
rect 59200 49058 60000 49088
rect 57973 49056 60000 49058
rect 57973 49000 57978 49056
rect 58034 49000 60000 49056
rect 57973 48998 60000 49000
rect 57973 48995 58039 48998
rect 19570 48992 19886 48993
rect 0 48922 800 48952
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 59200 48968 60000 48998
rect 50290 48927 50606 48928
rect 1669 48922 1735 48925
rect 0 48920 1735 48922
rect 0 48864 1674 48920
rect 1730 48864 1735 48920
rect 0 48862 1735 48864
rect 0 48832 800 48862
rect 1669 48859 1735 48862
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 59200 48424 60000 48544
rect 34930 48383 35246 48384
rect 0 48242 800 48272
rect 1669 48242 1735 48245
rect 0 48240 1735 48242
rect 0 48184 1674 48240
rect 1730 48184 1735 48240
rect 0 48182 1735 48184
rect 0 48152 800 48182
rect 1669 48179 1735 48182
rect 57237 47970 57303 47973
rect 59200 47970 60000 48000
rect 57237 47968 60000 47970
rect 57237 47912 57242 47968
rect 57298 47912 60000 47968
rect 57237 47910 60000 47912
rect 57237 47907 57303 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 59200 47880 60000 47910
rect 50290 47839 50606 47840
rect 26417 47698 26483 47701
rect 41822 47698 41828 47700
rect 26417 47696 41828 47698
rect 26417 47640 26422 47696
rect 26478 47640 41828 47696
rect 26417 47638 41828 47640
rect 26417 47635 26483 47638
rect 41822 47636 41828 47638
rect 41892 47636 41898 47700
rect 0 47562 800 47592
rect 1669 47562 1735 47565
rect 0 47560 1735 47562
rect 0 47504 1674 47560
rect 1730 47504 1735 47560
rect 0 47502 1735 47504
rect 0 47472 800 47502
rect 1669 47499 1735 47502
rect 1853 47562 1919 47565
rect 30230 47562 30236 47564
rect 1853 47560 30236 47562
rect 1853 47504 1858 47560
rect 1914 47504 30236 47560
rect 1853 47502 30236 47504
rect 1853 47499 1919 47502
rect 30230 47500 30236 47502
rect 30300 47500 30306 47564
rect 57973 47426 58039 47429
rect 59200 47426 60000 47456
rect 57973 47424 60000 47426
rect 57973 47368 57978 47424
rect 58034 47368 60000 47424
rect 57973 47366 60000 47368
rect 57973 47363 58039 47366
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 59200 47336 60000 47366
rect 34930 47295 35246 47296
rect 0 46882 800 46912
rect 1577 46882 1643 46885
rect 0 46880 1643 46882
rect 0 46824 1582 46880
rect 1638 46824 1643 46880
rect 0 46822 1643 46824
rect 0 46792 800 46822
rect 1577 46819 1643 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 59200 46792 60000 46912
rect 50290 46751 50606 46752
rect 57881 46338 57947 46341
rect 59200 46338 60000 46368
rect 57881 46336 60000 46338
rect 57881 46280 57886 46336
rect 57942 46280 60000 46336
rect 57881 46278 60000 46280
rect 57881 46275 57947 46278
rect 4210 46272 4526 46273
rect 0 46202 800 46232
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 1577 46202 1643 46205
rect 0 46200 1643 46202
rect 0 46144 1582 46200
rect 1638 46144 1643 46200
rect 0 46142 1643 46144
rect 0 46112 800 46142
rect 1577 46139 1643 46142
rect 57973 45794 58039 45797
rect 59200 45794 60000 45824
rect 57973 45792 60000 45794
rect 57973 45736 57978 45792
rect 58034 45736 60000 45792
rect 57973 45734 60000 45736
rect 57973 45731 58039 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 59200 45704 60000 45734
rect 50290 45663 50606 45664
rect 0 45522 800 45552
rect 1669 45522 1735 45525
rect 0 45520 1735 45522
rect 0 45464 1674 45520
rect 1730 45464 1735 45520
rect 0 45462 1735 45464
rect 0 45432 800 45462
rect 1669 45459 1735 45462
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 59200 45160 60000 45280
rect 34930 45119 35246 45120
rect 0 44842 800 44872
rect 1577 44842 1643 44845
rect 0 44840 1643 44842
rect 0 44784 1582 44840
rect 1638 44784 1643 44840
rect 0 44782 1643 44784
rect 0 44752 800 44782
rect 1577 44779 1643 44782
rect 57237 44706 57303 44709
rect 59200 44706 60000 44736
rect 57237 44704 60000 44706
rect 57237 44648 57242 44704
rect 57298 44648 60000 44704
rect 57237 44646 60000 44648
rect 57237 44643 57303 44646
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 59200 44616 60000 44646
rect 50290 44575 50606 44576
rect 0 44162 800 44192
rect 1669 44162 1735 44165
rect 0 44160 1735 44162
rect 0 44104 1674 44160
rect 1730 44104 1735 44160
rect 0 44102 1735 44104
rect 0 44072 800 44102
rect 1669 44099 1735 44102
rect 57881 44162 57947 44165
rect 59200 44162 60000 44192
rect 57881 44160 60000 44162
rect 57881 44104 57886 44160
rect 57942 44104 60000 44160
rect 57881 44102 60000 44104
rect 57881 44099 57947 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 59200 44072 60000 44102
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 59200 43528 60000 43648
rect 50290 43487 50606 43488
rect 1669 43482 1735 43485
rect 0 43480 1735 43482
rect 0 43424 1674 43480
rect 1730 43424 1735 43480
rect 0 43422 1735 43424
rect 0 43392 800 43422
rect 1669 43419 1735 43422
rect 58157 43074 58223 43077
rect 59200 43074 60000 43104
rect 58157 43072 60000 43074
rect 58157 43016 58162 43072
rect 58218 43016 60000 43072
rect 58157 43014 60000 43016
rect 58157 43011 58223 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 59200 42984 60000 43014
rect 34930 42943 35246 42944
rect 34513 42938 34579 42941
rect 34646 42938 34652 42940
rect 34513 42936 34652 42938
rect 34513 42880 34518 42936
rect 34574 42880 34652 42936
rect 34513 42878 34652 42880
rect 34513 42875 34579 42878
rect 34646 42876 34652 42878
rect 34716 42876 34722 42940
rect 0 42802 800 42832
rect 1577 42802 1643 42805
rect 0 42800 1643 42802
rect 0 42744 1582 42800
rect 1638 42744 1643 42800
rect 0 42742 1643 42744
rect 0 42712 800 42742
rect 1577 42739 1643 42742
rect 36905 42666 36971 42669
rect 42926 42666 42932 42668
rect 36905 42664 42932 42666
rect 36905 42608 36910 42664
rect 36966 42608 42932 42664
rect 36905 42606 42932 42608
rect 36905 42603 36971 42606
rect 42926 42604 42932 42606
rect 42996 42604 43002 42668
rect 57053 42530 57119 42533
rect 59200 42530 60000 42560
rect 57053 42528 60000 42530
rect 57053 42472 57058 42528
rect 57114 42472 60000 42528
rect 57053 42470 60000 42472
rect 57053 42467 57119 42470
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 59200 42440 60000 42470
rect 50290 42399 50606 42400
rect 0 42122 800 42152
rect 1669 42122 1735 42125
rect 0 42120 1735 42122
rect 0 42064 1674 42120
rect 1730 42064 1735 42120
rect 0 42062 1735 42064
rect 0 42032 800 42062
rect 1669 42059 1735 42062
rect 57973 41986 58039 41989
rect 59200 41986 60000 42016
rect 57973 41984 60000 41986
rect 57973 41928 57978 41984
rect 58034 41928 60000 41984
rect 57973 41926 60000 41928
rect 57973 41923 58039 41926
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 59200 41896 60000 41926
rect 34930 41855 35246 41856
rect 24577 41578 24643 41581
rect 29862 41578 29868 41580
rect 24577 41576 29868 41578
rect 24577 41520 24582 41576
rect 24638 41520 29868 41576
rect 24577 41518 29868 41520
rect 24577 41515 24643 41518
rect 29862 41516 29868 41518
rect 29932 41516 29938 41580
rect 0 41442 800 41472
rect 1669 41442 1735 41445
rect 0 41440 1735 41442
rect 0 41384 1674 41440
rect 1730 41384 1735 41440
rect 0 41382 1735 41384
rect 0 41352 800 41382
rect 1669 41379 1735 41382
rect 57237 41442 57303 41445
rect 59200 41442 60000 41472
rect 57237 41440 60000 41442
rect 57237 41384 57242 41440
rect 57298 41384 60000 41440
rect 57237 41382 60000 41384
rect 57237 41379 57303 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 59200 41352 60000 41382
rect 50290 41311 50606 41312
rect 57881 40898 57947 40901
rect 59200 40898 60000 40928
rect 57881 40896 60000 40898
rect 57881 40840 57886 40896
rect 57942 40840 60000 40896
rect 57881 40838 60000 40840
rect 57881 40835 57947 40838
rect 4210 40832 4526 40833
rect 0 40762 800 40792
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 1669 40762 1735 40765
rect 0 40760 1735 40762
rect 0 40704 1674 40760
rect 1730 40704 1735 40760
rect 0 40702 1735 40704
rect 0 40672 800 40702
rect 1669 40699 1735 40702
rect 56961 40354 57027 40357
rect 59200 40354 60000 40384
rect 56961 40352 60000 40354
rect 56961 40296 56966 40352
rect 57022 40296 60000 40352
rect 56961 40294 60000 40296
rect 56961 40291 57027 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 59200 40264 60000 40294
rect 50290 40223 50606 40224
rect 0 40082 800 40112
rect 1669 40082 1735 40085
rect 0 40080 1735 40082
rect 0 40024 1674 40080
rect 1730 40024 1735 40080
rect 0 40022 1735 40024
rect 0 39992 800 40022
rect 1669 40019 1735 40022
rect 57881 39810 57947 39813
rect 59200 39810 60000 39840
rect 57881 39808 60000 39810
rect 57881 39752 57886 39808
rect 57942 39752 60000 39808
rect 57881 39750 60000 39752
rect 57881 39747 57947 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 59200 39720 60000 39750
rect 34930 39679 35246 39680
rect 0 39402 800 39432
rect 1669 39402 1735 39405
rect 0 39400 1735 39402
rect 0 39344 1674 39400
rect 1730 39344 1735 39400
rect 0 39342 1735 39344
rect 0 39312 800 39342
rect 1669 39339 1735 39342
rect 57053 39266 57119 39269
rect 59200 39266 60000 39296
rect 57053 39264 60000 39266
rect 57053 39208 57058 39264
rect 57114 39208 60000 39264
rect 57053 39206 60000 39208
rect 57053 39203 57119 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 59200 39176 60000 39206
rect 50290 39135 50606 39136
rect 0 38722 800 38752
rect 1669 38722 1735 38725
rect 0 38720 1735 38722
rect 0 38664 1674 38720
rect 1730 38664 1735 38720
rect 0 38662 1735 38664
rect 0 38632 800 38662
rect 1669 38659 1735 38662
rect 57973 38722 58039 38725
rect 59200 38722 60000 38752
rect 57973 38720 60000 38722
rect 57973 38664 57978 38720
rect 58034 38664 60000 38720
rect 57973 38662 60000 38664
rect 57973 38659 58039 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 59200 38632 60000 38662
rect 34930 38591 35246 38592
rect 22093 38586 22159 38589
rect 23197 38586 23263 38589
rect 23790 38586 23796 38588
rect 22093 38584 23796 38586
rect 22093 38528 22098 38584
rect 22154 38528 23202 38584
rect 23258 38528 23796 38584
rect 22093 38526 23796 38528
rect 22093 38523 22159 38526
rect 23197 38523 23263 38526
rect 23790 38524 23796 38526
rect 23860 38524 23866 38588
rect 58157 38178 58223 38181
rect 59200 38178 60000 38208
rect 58157 38176 60000 38178
rect 58157 38120 58162 38176
rect 58218 38120 60000 38176
rect 58157 38118 60000 38120
rect 58157 38115 58223 38118
rect 19570 38112 19886 38113
rect 0 38042 800 38072
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 59200 38088 60000 38118
rect 50290 38047 50606 38048
rect 1669 38042 1735 38045
rect 0 38040 1735 38042
rect 0 37984 1674 38040
rect 1730 37984 1735 38040
rect 0 37982 1735 37984
rect 0 37952 800 37982
rect 1669 37979 1735 37982
rect 19517 37906 19583 37909
rect 25589 37906 25655 37909
rect 26049 37906 26115 37909
rect 19517 37904 26115 37906
rect 19517 37848 19522 37904
rect 19578 37848 25594 37904
rect 25650 37848 26054 37904
rect 26110 37848 26115 37904
rect 19517 37846 26115 37848
rect 19517 37843 19583 37846
rect 25589 37843 25655 37846
rect 26049 37843 26115 37846
rect 58065 37634 58131 37637
rect 59200 37634 60000 37664
rect 58065 37632 60000 37634
rect 58065 37576 58070 37632
rect 58126 37576 60000 37632
rect 58065 37574 60000 37576
rect 58065 37571 58131 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 59200 37544 60000 37574
rect 34930 37503 35246 37504
rect 0 37362 800 37392
rect 1669 37362 1735 37365
rect 0 37360 1735 37362
rect 0 37304 1674 37360
rect 1730 37304 1735 37360
rect 0 37302 1735 37304
rect 0 37272 800 37302
rect 1669 37299 1735 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 59200 37000 60000 37120
rect 50290 36959 50606 36960
rect 0 36682 800 36712
rect 3049 36682 3115 36685
rect 0 36680 3115 36682
rect 0 36624 3054 36680
rect 3110 36624 3115 36680
rect 0 36622 3115 36624
rect 0 36592 800 36622
rect 3049 36619 3115 36622
rect 17953 36682 18019 36685
rect 19149 36682 19215 36685
rect 17953 36680 19215 36682
rect 17953 36624 17958 36680
rect 18014 36624 19154 36680
rect 19210 36624 19215 36680
rect 17953 36622 19215 36624
rect 17953 36619 18019 36622
rect 19149 36619 19215 36622
rect 58157 36546 58223 36549
rect 59200 36546 60000 36576
rect 58157 36544 60000 36546
rect 58157 36488 58162 36544
rect 58218 36488 60000 36544
rect 58157 36486 60000 36488
rect 58157 36483 58223 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 59200 36456 60000 36486
rect 34930 36415 35246 36416
rect 0 36002 800 36032
rect 1669 36002 1735 36005
rect 0 36000 1735 36002
rect 0 35944 1674 36000
rect 1730 35944 1735 36000
rect 0 35942 1735 35944
rect 0 35912 800 35942
rect 1669 35939 1735 35942
rect 22645 36002 22711 36005
rect 23238 36002 23244 36004
rect 22645 36000 23244 36002
rect 22645 35944 22650 36000
rect 22706 35944 23244 36000
rect 22645 35942 23244 35944
rect 22645 35939 22711 35942
rect 23238 35940 23244 35942
rect 23308 35940 23314 36004
rect 57973 36002 58039 36005
rect 59200 36002 60000 36032
rect 57973 36000 60000 36002
rect 57973 35944 57978 36000
rect 58034 35944 60000 36000
rect 57973 35942 60000 35944
rect 57973 35939 58039 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 59200 35912 60000 35942
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35488
rect 34930 35327 35246 35328
rect 1669 35322 1735 35325
rect 0 35320 1735 35322
rect 0 35264 1674 35320
rect 1730 35264 1735 35320
rect 0 35262 1735 35264
rect 0 35232 800 35262
rect 1669 35259 1735 35262
rect 19701 35050 19767 35053
rect 20161 35050 20227 35053
rect 23013 35050 23079 35053
rect 23473 35050 23539 35053
rect 19701 35048 23539 35050
rect 19701 34992 19706 35048
rect 19762 34992 20166 35048
rect 20222 34992 23018 35048
rect 23074 34992 23478 35048
rect 23534 34992 23539 35048
rect 19701 34990 23539 34992
rect 19701 34987 19767 34990
rect 20161 34987 20227 34990
rect 23013 34987 23079 34990
rect 23473 34987 23539 34990
rect 58157 34914 58223 34917
rect 59200 34914 60000 34944
rect 58157 34912 60000 34914
rect 58157 34856 58162 34912
rect 58218 34856 60000 34912
rect 58157 34854 60000 34856
rect 58157 34851 58223 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 59200 34824 60000 34854
rect 50290 34783 50606 34784
rect 0 34642 800 34672
rect 1669 34642 1735 34645
rect 0 34640 1735 34642
rect 0 34584 1674 34640
rect 1730 34584 1735 34640
rect 0 34582 1735 34584
rect 0 34552 800 34582
rect 1669 34579 1735 34582
rect 22093 34642 22159 34645
rect 23841 34642 23907 34645
rect 22093 34640 23907 34642
rect 22093 34584 22098 34640
rect 22154 34584 23846 34640
rect 23902 34584 23907 34640
rect 22093 34582 23907 34584
rect 22093 34579 22159 34582
rect 23841 34579 23907 34582
rect 22185 34506 22251 34509
rect 22686 34506 22692 34508
rect 22185 34504 22692 34506
rect 22185 34448 22190 34504
rect 22246 34448 22692 34504
rect 22185 34446 22692 34448
rect 22185 34443 22251 34446
rect 22686 34444 22692 34446
rect 22756 34444 22762 34508
rect 57881 34370 57947 34373
rect 59200 34370 60000 34400
rect 57881 34368 60000 34370
rect 57881 34312 57886 34368
rect 57942 34312 60000 34368
rect 57881 34310 60000 34312
rect 57881 34307 57947 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 59200 34280 60000 34310
rect 34930 34239 35246 34240
rect 0 33962 800 33992
rect 1669 33962 1735 33965
rect 0 33960 1735 33962
rect 0 33904 1674 33960
rect 1730 33904 1735 33960
rect 0 33902 1735 33904
rect 0 33872 800 33902
rect 1669 33899 1735 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 59200 33736 60000 33856
rect 50290 33695 50606 33696
rect 0 33282 800 33312
rect 1669 33282 1735 33285
rect 0 33280 1735 33282
rect 0 33224 1674 33280
rect 1730 33224 1735 33280
rect 0 33222 1735 33224
rect 0 33192 800 33222
rect 1669 33219 1735 33222
rect 58157 33282 58223 33285
rect 59200 33282 60000 33312
rect 58157 33280 60000 33282
rect 58157 33224 58162 33280
rect 58218 33224 60000 33280
rect 58157 33222 60000 33224
rect 58157 33219 58223 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 59200 33192 60000 33222
rect 34930 33151 35246 33152
rect 57053 32738 57119 32741
rect 59200 32738 60000 32768
rect 57053 32736 60000 32738
rect 57053 32680 57058 32736
rect 57114 32680 60000 32736
rect 57053 32678 60000 32680
rect 57053 32675 57119 32678
rect 19570 32672 19886 32673
rect 0 32602 800 32632
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 59200 32648 60000 32678
rect 50290 32607 50606 32608
rect 1669 32602 1735 32605
rect 0 32600 1735 32602
rect 0 32544 1674 32600
rect 1730 32544 1735 32600
rect 0 32542 1735 32544
rect 0 32512 800 32542
rect 1669 32539 1735 32542
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 59200 32104 60000 32224
rect 34930 32063 35246 32064
rect 0 31922 800 31952
rect 1669 31922 1735 31925
rect 0 31920 1735 31922
rect 0 31864 1674 31920
rect 1730 31864 1735 31920
rect 0 31862 1735 31864
rect 0 31832 800 31862
rect 1669 31859 1735 31862
rect 57789 31650 57855 31653
rect 59200 31650 60000 31680
rect 57789 31648 60000 31650
rect 57789 31592 57794 31648
rect 57850 31592 60000 31648
rect 57789 31590 60000 31592
rect 57789 31587 57855 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 59200 31560 60000 31590
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 1669 31242 1735 31245
rect 0 31240 1735 31242
rect 0 31184 1674 31240
rect 1730 31184 1735 31240
rect 0 31182 1735 31184
rect 0 31152 800 31182
rect 1669 31179 1735 31182
rect 58065 31106 58131 31109
rect 59200 31106 60000 31136
rect 58065 31104 60000 31106
rect 58065 31048 58070 31104
rect 58126 31048 60000 31104
rect 58065 31046 60000 31048
rect 58065 31043 58131 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 59200 31016 60000 31046
rect 34930 30975 35246 30976
rect 17534 30636 17540 30700
rect 17604 30698 17610 30700
rect 20069 30698 20135 30701
rect 17604 30696 20135 30698
rect 17604 30640 20074 30696
rect 20130 30640 20135 30696
rect 17604 30638 20135 30640
rect 17604 30636 17610 30638
rect 20069 30635 20135 30638
rect 0 30562 800 30592
rect 1669 30562 1735 30565
rect 0 30560 1735 30562
rect 0 30504 1674 30560
rect 1730 30504 1735 30560
rect 0 30502 1735 30504
rect 0 30472 800 30502
rect 1669 30499 1735 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 59200 30472 60000 30592
rect 50290 30431 50606 30432
rect 25129 30290 25195 30293
rect 25681 30290 25747 30293
rect 25129 30288 25747 30290
rect 25129 30232 25134 30288
rect 25190 30232 25686 30288
rect 25742 30232 25747 30288
rect 25129 30230 25747 30232
rect 25129 30227 25195 30230
rect 25681 30227 25747 30230
rect 23933 30154 23999 30157
rect 26325 30154 26391 30157
rect 23933 30152 26391 30154
rect 23933 30096 23938 30152
rect 23994 30096 26330 30152
rect 26386 30096 26391 30152
rect 23933 30094 26391 30096
rect 23933 30091 23999 30094
rect 26325 30091 26391 30094
rect 58157 30018 58223 30021
rect 59200 30018 60000 30048
rect 58157 30016 60000 30018
rect 58157 29960 58162 30016
rect 58218 29960 60000 30016
rect 58157 29958 60000 29960
rect 58157 29955 58223 29958
rect 4210 29952 4526 29953
rect 0 29882 800 29912
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 1761 29882 1827 29885
rect 0 29880 1827 29882
rect 0 29824 1766 29880
rect 1822 29824 1827 29880
rect 0 29822 1827 29824
rect 0 29792 800 29822
rect 1761 29819 1827 29822
rect 57053 29474 57119 29477
rect 59200 29474 60000 29504
rect 57053 29472 60000 29474
rect 57053 29416 57058 29472
rect 57114 29416 60000 29472
rect 57053 29414 60000 29416
rect 57053 29411 57119 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 59200 29384 60000 29414
rect 50290 29343 50606 29344
rect 0 29202 800 29232
rect 1853 29202 1919 29205
rect 0 29200 1919 29202
rect 0 29144 1858 29200
rect 1914 29144 1919 29200
rect 0 29142 1919 29144
rect 0 29112 800 29142
rect 1853 29139 1919 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 59200 28840 60000 28960
rect 34930 28799 35246 28800
rect 0 28522 800 28552
rect 1853 28522 1919 28525
rect 0 28520 1919 28522
rect 0 28464 1858 28520
rect 1914 28464 1919 28520
rect 0 28462 1919 28464
rect 0 28432 800 28462
rect 1853 28459 1919 28462
rect 16062 28460 16068 28524
rect 16132 28522 16138 28524
rect 22553 28522 22619 28525
rect 16132 28520 22619 28522
rect 16132 28464 22558 28520
rect 22614 28464 22619 28520
rect 16132 28462 22619 28464
rect 16132 28460 16138 28462
rect 22553 28459 22619 28462
rect 58157 28386 58223 28389
rect 59200 28386 60000 28416
rect 58157 28384 60000 28386
rect 58157 28328 58162 28384
rect 58218 28328 60000 28384
rect 58157 28326 60000 28328
rect 58157 28323 58223 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 59200 28296 60000 28326
rect 50290 28255 50606 28256
rect 0 27842 800 27872
rect 1761 27842 1827 27845
rect 0 27840 1827 27842
rect 0 27784 1766 27840
rect 1822 27784 1827 27840
rect 0 27782 1827 27784
rect 0 27752 800 27782
rect 1761 27779 1827 27782
rect 58065 27842 58131 27845
rect 59200 27842 60000 27872
rect 58065 27840 60000 27842
rect 58065 27784 58070 27840
rect 58126 27784 60000 27840
rect 58065 27782 60000 27784
rect 58065 27779 58131 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 59200 27752 60000 27782
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 59200 27208 60000 27328
rect 50290 27167 50606 27168
rect 1853 27162 1919 27165
rect 0 27160 1919 27162
rect 0 27104 1858 27160
rect 1914 27104 1919 27160
rect 0 27102 1919 27104
rect 0 27072 800 27102
rect 1853 27099 1919 27102
rect 16430 26964 16436 27028
rect 16500 27026 16506 27028
rect 27153 27026 27219 27029
rect 16500 27024 27219 27026
rect 16500 26968 27158 27024
rect 27214 26968 27219 27024
rect 16500 26966 27219 26968
rect 16500 26964 16506 26966
rect 27153 26963 27219 26966
rect 10501 26890 10567 26893
rect 34094 26890 34100 26892
rect 10501 26888 34100 26890
rect 10501 26832 10506 26888
rect 10562 26832 34100 26888
rect 10501 26830 34100 26832
rect 10501 26827 10567 26830
rect 34094 26828 34100 26830
rect 34164 26828 34170 26892
rect 36670 26828 36676 26892
rect 36740 26890 36746 26892
rect 58525 26890 58591 26893
rect 36740 26888 58591 26890
rect 36740 26832 58530 26888
rect 58586 26832 58591 26888
rect 36740 26830 58591 26832
rect 36740 26828 36746 26830
rect 58525 26827 58591 26830
rect 58157 26754 58223 26757
rect 59200 26754 60000 26784
rect 58157 26752 60000 26754
rect 58157 26696 58162 26752
rect 58218 26696 60000 26752
rect 58157 26694 60000 26696
rect 58157 26691 58223 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 59200 26664 60000 26694
rect 34930 26623 35246 26624
rect 0 26482 800 26512
rect 1761 26482 1827 26485
rect 0 26480 1827 26482
rect 0 26424 1766 26480
rect 1822 26424 1827 26480
rect 0 26422 1827 26424
rect 0 26392 800 26422
rect 1761 26419 1827 26422
rect 31017 26346 31083 26349
rect 36302 26346 36308 26348
rect 31017 26344 36308 26346
rect 31017 26288 31022 26344
rect 31078 26288 36308 26344
rect 31017 26286 36308 26288
rect 31017 26283 31083 26286
rect 36302 26284 36308 26286
rect 36372 26284 36378 26348
rect 57053 26210 57119 26213
rect 59200 26210 60000 26240
rect 57053 26208 60000 26210
rect 57053 26152 57058 26208
rect 57114 26152 60000 26208
rect 57053 26150 60000 26152
rect 57053 26147 57119 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 59200 26120 60000 26150
rect 50290 26079 50606 26080
rect 0 25802 800 25832
rect 1761 25802 1827 25805
rect 0 25800 1827 25802
rect 0 25744 1766 25800
rect 1822 25744 1827 25800
rect 0 25742 1827 25744
rect 0 25712 800 25742
rect 1761 25739 1827 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 59200 25576 60000 25696
rect 34930 25535 35246 25536
rect 0 25122 800 25152
rect 1853 25122 1919 25125
rect 0 25120 1919 25122
rect 0 25064 1858 25120
rect 1914 25064 1919 25120
rect 0 25062 1919 25064
rect 0 25032 800 25062
rect 1853 25059 1919 25062
rect 58157 25122 58223 25125
rect 59200 25122 60000 25152
rect 58157 25120 60000 25122
rect 58157 25064 58162 25120
rect 58218 25064 60000 25120
rect 58157 25062 60000 25064
rect 58157 25059 58223 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 59200 25032 60000 25062
rect 50290 24991 50606 24992
rect 22134 24788 22140 24852
rect 22204 24850 22210 24852
rect 26877 24850 26943 24853
rect 22204 24848 26943 24850
rect 22204 24792 26882 24848
rect 26938 24792 26943 24848
rect 22204 24790 26943 24792
rect 22204 24788 22210 24790
rect 26877 24787 26943 24790
rect 58065 24578 58131 24581
rect 59200 24578 60000 24608
rect 58065 24576 60000 24578
rect 58065 24520 58070 24576
rect 58126 24520 60000 24576
rect 58065 24518 60000 24520
rect 58065 24515 58131 24518
rect 4210 24512 4526 24513
rect 0 24442 800 24472
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 60000 24518
rect 34930 24447 35246 24448
rect 1761 24442 1827 24445
rect 0 24440 1827 24442
rect 0 24384 1766 24440
rect 1822 24384 1827 24440
rect 0 24382 1827 24384
rect 0 24352 800 24382
rect 1761 24379 1827 24382
rect 17217 24306 17283 24309
rect 20110 24306 20116 24308
rect 17217 24304 20116 24306
rect 17217 24248 17222 24304
rect 17278 24248 20116 24304
rect 17217 24246 20116 24248
rect 17217 24243 17283 24246
rect 20110 24244 20116 24246
rect 20180 24244 20186 24308
rect 19425 24170 19491 24173
rect 39430 24170 39436 24172
rect 19425 24168 39436 24170
rect 19425 24112 19430 24168
rect 19486 24112 39436 24168
rect 19425 24110 39436 24112
rect 19425 24107 19491 24110
rect 39430 24108 39436 24110
rect 39500 24108 39506 24172
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 59200 23944 60000 24064
rect 50290 23903 50606 23904
rect 0 23762 800 23792
rect 1853 23762 1919 23765
rect 0 23760 1919 23762
rect 0 23704 1858 23760
rect 1914 23704 1919 23760
rect 0 23702 1919 23704
rect 0 23672 800 23702
rect 1853 23699 1919 23702
rect 23841 23490 23907 23493
rect 23974 23490 23980 23492
rect 23841 23488 23980 23490
rect 23841 23432 23846 23488
rect 23902 23432 23980 23488
rect 23841 23430 23980 23432
rect 23841 23427 23907 23430
rect 23974 23428 23980 23430
rect 24044 23428 24050 23492
rect 58157 23490 58223 23493
rect 59200 23490 60000 23520
rect 58157 23488 60000 23490
rect 58157 23432 58162 23488
rect 58218 23432 60000 23488
rect 58157 23430 60000 23432
rect 58157 23427 58223 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 59200 23400 60000 23430
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 1853 23082 1919 23085
rect 0 23080 1919 23082
rect 0 23024 1858 23080
rect 1914 23024 1919 23080
rect 0 23022 1919 23024
rect 0 22992 800 23022
rect 1853 23019 1919 23022
rect 58065 22946 58131 22949
rect 59200 22946 60000 22976
rect 58065 22944 60000 22946
rect 58065 22888 58070 22944
rect 58126 22888 60000 22944
rect 58065 22886 60000 22888
rect 58065 22883 58131 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 59200 22856 60000 22886
rect 50290 22815 50606 22816
rect 28441 22810 28507 22813
rect 40718 22810 40724 22812
rect 28441 22808 40724 22810
rect 28441 22752 28446 22808
rect 28502 22752 40724 22808
rect 28441 22750 40724 22752
rect 28441 22747 28507 22750
rect 40718 22748 40724 22750
rect 40788 22748 40794 22812
rect 22737 22674 22803 22677
rect 41270 22674 41276 22676
rect 22737 22672 41276 22674
rect 22737 22616 22742 22672
rect 22798 22616 41276 22672
rect 22737 22614 41276 22616
rect 22737 22611 22803 22614
rect 41270 22612 41276 22614
rect 41340 22612 41346 22676
rect 0 22402 800 22432
rect 1761 22402 1827 22405
rect 0 22400 1827 22402
rect 0 22344 1766 22400
rect 1822 22344 1827 22400
rect 0 22342 1827 22344
rect 0 22312 800 22342
rect 1761 22339 1827 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 59200 22312 60000 22432
rect 34930 22271 35246 22272
rect 20294 22068 20300 22132
rect 20364 22130 20370 22132
rect 21449 22130 21515 22133
rect 20364 22128 21515 22130
rect 20364 22072 21454 22128
rect 21510 22072 21515 22128
rect 20364 22070 21515 22072
rect 20364 22068 20370 22070
rect 21449 22067 21515 22070
rect 14406 21932 14412 21996
rect 14476 21994 14482 21996
rect 27429 21994 27495 21997
rect 14476 21992 27495 21994
rect 14476 21936 27434 21992
rect 27490 21936 27495 21992
rect 14476 21934 27495 21936
rect 14476 21932 14482 21934
rect 27429 21931 27495 21934
rect 58157 21858 58223 21861
rect 59200 21858 60000 21888
rect 58157 21856 60000 21858
rect 58157 21800 58162 21856
rect 58218 21800 60000 21856
rect 58157 21798 60000 21800
rect 58157 21795 58223 21798
rect 19570 21792 19886 21793
rect 0 21722 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 59200 21768 60000 21798
rect 50290 21727 50606 21728
rect 1853 21722 1919 21725
rect 0 21720 1919 21722
rect 0 21664 1858 21720
rect 1914 21664 1919 21720
rect 0 21662 1919 21664
rect 0 21632 800 21662
rect 1853 21659 1919 21662
rect 58065 21314 58131 21317
rect 59200 21314 60000 21344
rect 58065 21312 60000 21314
rect 58065 21256 58070 21312
rect 58126 21256 60000 21312
rect 58065 21254 60000 21256
rect 58065 21251 58131 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 59200 21224 60000 21254
rect 34930 21183 35246 21184
rect 0 21042 800 21072
rect 1761 21042 1827 21045
rect 0 21040 1827 21042
rect 0 20984 1766 21040
rect 1822 20984 1827 21040
rect 0 20982 1827 20984
rect 0 20952 800 20982
rect 1761 20979 1827 20982
rect 38009 20770 38075 20773
rect 40534 20770 40540 20772
rect 38009 20768 40540 20770
rect 38009 20712 38014 20768
rect 38070 20712 40540 20768
rect 38009 20710 40540 20712
rect 38009 20707 38075 20710
rect 40534 20708 40540 20710
rect 40604 20708 40610 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 59200 20680 60000 20800
rect 50290 20639 50606 20640
rect 0 20362 800 20392
rect 1761 20362 1827 20365
rect 0 20360 1827 20362
rect 0 20304 1766 20360
rect 1822 20304 1827 20360
rect 0 20302 1827 20304
rect 0 20272 800 20302
rect 1761 20299 1827 20302
rect 58157 20226 58223 20229
rect 59200 20226 60000 20256
rect 58157 20224 60000 20226
rect 58157 20168 58162 20224
rect 58218 20168 60000 20224
rect 58157 20166 60000 20168
rect 58157 20163 58223 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 59200 20136 60000 20166
rect 34930 20095 35246 20096
rect 24761 19954 24827 19957
rect 25221 19954 25287 19957
rect 24761 19952 25287 19954
rect 24761 19896 24766 19952
rect 24822 19896 25226 19952
rect 25282 19896 25287 19952
rect 24761 19894 25287 19896
rect 24761 19891 24827 19894
rect 25221 19891 25287 19894
rect 18045 19818 18111 19821
rect 22093 19818 22159 19821
rect 18045 19816 22159 19818
rect 18045 19760 18050 19816
rect 18106 19760 22098 19816
rect 22154 19760 22159 19816
rect 18045 19758 22159 19760
rect 18045 19755 18111 19758
rect 22093 19755 22159 19758
rect 24577 19818 24643 19821
rect 25681 19818 25747 19821
rect 24577 19816 25747 19818
rect 24577 19760 24582 19816
rect 24638 19760 25686 19816
rect 25742 19760 25747 19816
rect 24577 19758 25747 19760
rect 24577 19755 24643 19758
rect 25681 19755 25747 19758
rect 0 19682 800 19712
rect 1853 19682 1919 19685
rect 0 19680 1919 19682
rect 0 19624 1858 19680
rect 1914 19624 1919 19680
rect 0 19622 1919 19624
rect 0 19592 800 19622
rect 1853 19619 1919 19622
rect 58065 19682 58131 19685
rect 59200 19682 60000 19712
rect 58065 19680 60000 19682
rect 58065 19624 58070 19680
rect 58126 19624 60000 19680
rect 58065 19622 60000 19624
rect 58065 19619 58131 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 59200 19592 60000 19622
rect 50290 19551 50606 19552
rect 21633 19546 21699 19549
rect 22185 19546 22251 19549
rect 22737 19546 22803 19549
rect 21633 19544 22803 19546
rect 21633 19488 21638 19544
rect 21694 19488 22190 19544
rect 22246 19488 22742 19544
rect 22798 19488 22803 19544
rect 21633 19486 22803 19488
rect 21633 19483 21699 19486
rect 22185 19483 22251 19486
rect 22737 19483 22803 19486
rect 35065 19546 35131 19549
rect 35801 19546 35867 19549
rect 35065 19544 35867 19546
rect 35065 19488 35070 19544
rect 35126 19488 35806 19544
rect 35862 19488 35867 19544
rect 35065 19486 35867 19488
rect 35065 19483 35131 19486
rect 35801 19483 35867 19486
rect 48221 19546 48287 19549
rect 48681 19546 48747 19549
rect 48221 19544 48747 19546
rect 48221 19488 48226 19544
rect 48282 19488 48686 19544
rect 48742 19488 48747 19544
rect 48221 19486 48747 19488
rect 48221 19483 48287 19486
rect 48681 19483 48747 19486
rect 22645 19410 22711 19413
rect 24761 19410 24827 19413
rect 21958 19408 24827 19410
rect 21958 19352 22650 19408
rect 22706 19352 24766 19408
rect 24822 19352 24827 19408
rect 21958 19350 24827 19352
rect 21958 19348 22067 19350
rect 21958 19292 22006 19348
rect 22062 19292 22067 19348
rect 22645 19347 22711 19350
rect 24761 19347 24827 19350
rect 47761 19410 47827 19413
rect 48957 19410 49023 19413
rect 47761 19408 49023 19410
rect 47761 19352 47766 19408
rect 47822 19352 48962 19408
rect 49018 19352 49023 19408
rect 47761 19350 49023 19352
rect 47761 19347 47827 19350
rect 48957 19347 49023 19350
rect 21958 19290 22067 19292
rect 22001 19287 22067 19290
rect 23749 19274 23815 19277
rect 34421 19274 34487 19277
rect 23749 19272 34487 19274
rect 23749 19216 23754 19272
rect 23810 19216 34426 19272
rect 34482 19216 34487 19272
rect 23749 19214 34487 19216
rect 23749 19211 23815 19214
rect 34421 19211 34487 19214
rect 40677 19274 40743 19277
rect 41229 19274 41295 19277
rect 40677 19272 41295 19274
rect 40677 19216 40682 19272
rect 40738 19216 41234 19272
rect 41290 19216 41295 19272
rect 40677 19214 41295 19216
rect 40677 19211 40743 19214
rect 41229 19211 41295 19214
rect 17585 19138 17651 19141
rect 18965 19138 19031 19141
rect 17585 19136 19031 19138
rect 17585 19080 17590 19136
rect 17646 19080 18970 19136
rect 19026 19080 19031 19136
rect 17585 19078 19031 19080
rect 17585 19075 17651 19078
rect 18965 19075 19031 19078
rect 22369 19138 22435 19141
rect 29269 19138 29335 19141
rect 22369 19136 29335 19138
rect 22369 19080 22374 19136
rect 22430 19080 29274 19136
rect 29330 19080 29335 19136
rect 22369 19078 29335 19080
rect 22369 19075 22435 19078
rect 29269 19075 29335 19078
rect 40585 19138 40651 19141
rect 48129 19138 48195 19141
rect 40585 19136 48195 19138
rect 40585 19080 40590 19136
rect 40646 19080 48134 19136
rect 48190 19080 48195 19136
rect 40585 19078 48195 19080
rect 40585 19075 40651 19078
rect 48129 19075 48195 19078
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19168
rect 34930 19007 35246 19008
rect 1853 19002 1919 19005
rect 39849 19004 39915 19005
rect 0 19000 1919 19002
rect 0 18944 1858 19000
rect 1914 18944 1919 19000
rect 0 18942 1919 18944
rect 0 18912 800 18942
rect 1853 18939 1919 18942
rect 39798 18940 39804 19004
rect 39868 19002 39915 19004
rect 39868 19000 39960 19002
rect 39910 18944 39960 19000
rect 39868 18942 39960 18944
rect 39868 18940 39915 18942
rect 39849 18939 39915 18940
rect 34881 18866 34947 18869
rect 36261 18866 36327 18869
rect 34881 18864 36327 18866
rect 34881 18808 34886 18864
rect 34942 18808 36266 18864
rect 36322 18808 36327 18864
rect 34881 18806 36327 18808
rect 34881 18803 34947 18806
rect 36261 18803 36327 18806
rect 48589 18866 48655 18869
rect 57881 18866 57947 18869
rect 48589 18864 57947 18866
rect 48589 18808 48594 18864
rect 48650 18808 57886 18864
rect 57942 18808 57947 18864
rect 48589 18806 57947 18808
rect 48589 18803 48655 18806
rect 57881 18803 57947 18806
rect 13302 18668 13308 18732
rect 13372 18730 13378 18732
rect 30281 18730 30347 18733
rect 13372 18728 30347 18730
rect 13372 18672 30286 18728
rect 30342 18672 30347 18728
rect 13372 18670 30347 18672
rect 13372 18668 13378 18670
rect 30281 18667 30347 18670
rect 48221 18730 48287 18733
rect 49141 18730 49207 18733
rect 48221 18728 49207 18730
rect 48221 18672 48226 18728
rect 48282 18672 49146 18728
rect 49202 18672 49207 18728
rect 48221 18670 49207 18672
rect 48221 18667 48287 18670
rect 49141 18667 49207 18670
rect 58157 18594 58223 18597
rect 59200 18594 60000 18624
rect 58157 18592 60000 18594
rect 58157 18536 58162 18592
rect 58218 18536 60000 18592
rect 58157 18534 60000 18536
rect 58157 18531 58223 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 59200 18504 60000 18534
rect 50290 18463 50606 18464
rect 0 18322 800 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 800 18262
rect 1853 18259 1919 18262
rect 24301 18322 24367 18325
rect 27521 18322 27587 18325
rect 24301 18320 27587 18322
rect 24301 18264 24306 18320
rect 24362 18264 27526 18320
rect 27582 18264 27587 18320
rect 24301 18262 27587 18264
rect 24301 18259 24367 18262
rect 27521 18259 27587 18262
rect 26049 18186 26115 18189
rect 27429 18186 27495 18189
rect 26049 18184 27495 18186
rect 26049 18128 26054 18184
rect 26110 18128 27434 18184
rect 27490 18128 27495 18184
rect 26049 18126 27495 18128
rect 26049 18123 26115 18126
rect 27429 18123 27495 18126
rect 14457 18050 14523 18053
rect 22737 18052 22803 18053
rect 17350 18050 17356 18052
rect 14457 18048 17356 18050
rect 14457 17992 14462 18048
rect 14518 17992 17356 18048
rect 14457 17990 17356 17992
rect 14457 17987 14523 17990
rect 17350 17988 17356 17990
rect 17420 17988 17426 18052
rect 22686 18050 22692 18052
rect 22646 17990 22692 18050
rect 22756 18048 22803 18052
rect 22798 17992 22803 18048
rect 22686 17988 22692 17990
rect 22756 17988 22803 17992
rect 22737 17987 22803 17988
rect 58065 18050 58131 18053
rect 59200 18050 60000 18080
rect 58065 18048 60000 18050
rect 58065 17992 58070 18048
rect 58126 17992 60000 18048
rect 58065 17990 60000 17992
rect 58065 17987 58131 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 59200 17960 60000 17990
rect 34930 17919 35246 17920
rect 17125 17914 17191 17917
rect 20662 17914 20668 17916
rect 17125 17912 20668 17914
rect 17125 17856 17130 17912
rect 17186 17856 20668 17912
rect 17125 17854 20668 17856
rect 17125 17851 17191 17854
rect 20662 17852 20668 17854
rect 20732 17852 20738 17916
rect 16757 17778 16823 17781
rect 21766 17778 21772 17780
rect 16757 17776 21772 17778
rect 16757 17720 16762 17776
rect 16818 17720 21772 17776
rect 16757 17718 21772 17720
rect 16757 17715 16823 17718
rect 21766 17716 21772 17718
rect 21836 17716 21842 17780
rect 24577 17778 24643 17781
rect 26417 17778 26483 17781
rect 24577 17776 26483 17778
rect 24577 17720 24582 17776
rect 24638 17720 26422 17776
rect 26478 17720 26483 17776
rect 24577 17718 26483 17720
rect 24577 17715 24643 17718
rect 26417 17715 26483 17718
rect 27889 17778 27955 17781
rect 28993 17778 29059 17781
rect 27889 17776 29059 17778
rect 27889 17720 27894 17776
rect 27950 17720 28998 17776
rect 29054 17720 29059 17776
rect 27889 17718 29059 17720
rect 27889 17715 27955 17718
rect 28993 17715 29059 17718
rect 34881 17778 34947 17781
rect 38101 17778 38167 17781
rect 34881 17776 38167 17778
rect 34881 17720 34886 17776
rect 34942 17720 38106 17776
rect 38162 17720 38167 17776
rect 34881 17718 38167 17720
rect 34881 17715 34947 17718
rect 38101 17715 38167 17718
rect 0 17642 800 17672
rect 1853 17642 1919 17645
rect 0 17640 1919 17642
rect 0 17584 1858 17640
rect 1914 17584 1919 17640
rect 0 17582 1919 17584
rect 0 17552 800 17582
rect 1853 17579 1919 17582
rect 21725 17642 21791 17645
rect 39205 17642 39271 17645
rect 21725 17640 39271 17642
rect 21725 17584 21730 17640
rect 21786 17584 39210 17640
rect 39266 17584 39271 17640
rect 21725 17582 39271 17584
rect 21725 17579 21791 17582
rect 39205 17579 39271 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 59200 17416 60000 17536
rect 50290 17375 50606 17376
rect 17401 17234 17467 17237
rect 17902 17234 17908 17236
rect 17401 17232 17908 17234
rect 17401 17176 17406 17232
rect 17462 17176 17908 17232
rect 17401 17174 17908 17176
rect 17401 17171 17467 17174
rect 17902 17172 17908 17174
rect 17972 17172 17978 17236
rect 31201 17098 31267 17101
rect 33685 17098 33751 17101
rect 31201 17096 33751 17098
rect 31201 17040 31206 17096
rect 31262 17040 33690 17096
rect 33746 17040 33751 17096
rect 31201 17038 33751 17040
rect 31201 17035 31267 17038
rect 33685 17035 33751 17038
rect 0 16962 800 16992
rect 1761 16962 1827 16965
rect 0 16960 1827 16962
rect 0 16904 1766 16960
rect 1822 16904 1827 16960
rect 0 16902 1827 16904
rect 0 16872 800 16902
rect 1761 16899 1827 16902
rect 18454 16900 18460 16964
rect 18524 16962 18530 16964
rect 18873 16962 18939 16965
rect 18524 16960 18939 16962
rect 18524 16904 18878 16960
rect 18934 16904 18939 16960
rect 18524 16902 18939 16904
rect 18524 16900 18530 16902
rect 18873 16899 18939 16902
rect 58157 16962 58223 16965
rect 59200 16962 60000 16992
rect 58157 16960 60000 16962
rect 58157 16904 58162 16960
rect 58218 16904 60000 16960
rect 58157 16902 60000 16904
rect 58157 16899 58223 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 59200 16872 60000 16902
rect 34930 16831 35246 16832
rect 35709 16690 35775 16693
rect 37181 16690 37247 16693
rect 37549 16690 37615 16693
rect 35709 16688 37615 16690
rect 35709 16632 35714 16688
rect 35770 16632 37186 16688
rect 37242 16632 37554 16688
rect 37610 16632 37615 16688
rect 35709 16630 37615 16632
rect 35709 16627 35775 16630
rect 37181 16627 37247 16630
rect 37549 16627 37615 16630
rect 27613 16418 27679 16421
rect 31109 16418 31175 16421
rect 27613 16416 31175 16418
rect 27613 16360 27618 16416
rect 27674 16360 31114 16416
rect 31170 16360 31175 16416
rect 27613 16358 31175 16360
rect 27613 16355 27679 16358
rect 31109 16355 31175 16358
rect 57053 16418 57119 16421
rect 59200 16418 60000 16448
rect 57053 16416 60000 16418
rect 57053 16360 57058 16416
rect 57114 16360 60000 16416
rect 57053 16358 60000 16360
rect 57053 16355 57119 16358
rect 19570 16352 19886 16353
rect 0 16282 800 16312
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 59200 16328 60000 16358
rect 50290 16287 50606 16288
rect 1853 16282 1919 16285
rect 0 16280 1919 16282
rect 0 16224 1858 16280
rect 1914 16224 1919 16280
rect 0 16222 1919 16224
rect 0 16192 800 16222
rect 1853 16219 1919 16222
rect 32121 16282 32187 16285
rect 33726 16282 33732 16284
rect 32121 16280 33732 16282
rect 32121 16224 32126 16280
rect 32182 16224 33732 16280
rect 32121 16222 33732 16224
rect 32121 16219 32187 16222
rect 33726 16220 33732 16222
rect 33796 16220 33802 16284
rect 30005 16010 30071 16013
rect 36905 16010 36971 16013
rect 30005 16008 36971 16010
rect 30005 15952 30010 16008
rect 30066 15952 36910 16008
rect 36966 15952 36971 16008
rect 30005 15950 36971 15952
rect 30005 15947 30071 15950
rect 36905 15947 36971 15950
rect 37222 15948 37228 16012
rect 37292 16010 37298 16012
rect 37733 16010 37799 16013
rect 37292 16008 37799 16010
rect 37292 15952 37738 16008
rect 37794 15952 37799 16008
rect 37292 15950 37799 15952
rect 37292 15948 37298 15950
rect 37733 15947 37799 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 59200 15784 60000 15904
rect 34930 15743 35246 15744
rect 30373 15738 30439 15741
rect 34053 15738 34119 15741
rect 30373 15736 34119 15738
rect 30373 15680 30378 15736
rect 30434 15680 34058 15736
rect 34114 15680 34119 15736
rect 30373 15678 34119 15680
rect 30373 15675 30439 15678
rect 34053 15675 34119 15678
rect 0 15602 800 15632
rect 1761 15602 1827 15605
rect 0 15600 1827 15602
rect 0 15544 1766 15600
rect 1822 15544 1827 15600
rect 0 15542 1827 15544
rect 0 15512 800 15542
rect 1761 15539 1827 15542
rect 17166 15540 17172 15604
rect 17236 15602 17242 15604
rect 19977 15602 20043 15605
rect 17236 15600 20043 15602
rect 17236 15544 19982 15600
rect 20038 15544 20043 15600
rect 17236 15542 20043 15544
rect 17236 15540 17242 15542
rect 19977 15539 20043 15542
rect 28993 15602 29059 15605
rect 35801 15602 35867 15605
rect 28993 15600 35867 15602
rect 28993 15544 28998 15600
rect 29054 15544 35806 15600
rect 35862 15544 35867 15600
rect 28993 15542 35867 15544
rect 28993 15539 29059 15542
rect 35801 15539 35867 15542
rect 14917 15466 14983 15469
rect 20478 15466 20484 15468
rect 14917 15464 20484 15466
rect 14917 15408 14922 15464
rect 14978 15408 20484 15464
rect 14917 15406 20484 15408
rect 14917 15403 14983 15406
rect 20478 15404 20484 15406
rect 20548 15404 20554 15468
rect 22001 15466 22067 15469
rect 37733 15466 37799 15469
rect 22001 15464 37799 15466
rect 22001 15408 22006 15464
rect 22062 15408 37738 15464
rect 37794 15408 37799 15464
rect 22001 15406 37799 15408
rect 22001 15403 22067 15406
rect 37733 15403 37799 15406
rect 38837 15466 38903 15469
rect 40585 15466 40651 15469
rect 38837 15464 40651 15466
rect 38837 15408 38842 15464
rect 38898 15408 40590 15464
rect 40646 15408 40651 15464
rect 38837 15406 40651 15408
rect 38837 15403 38903 15406
rect 40585 15403 40651 15406
rect 20529 15330 20595 15333
rect 42701 15330 42767 15333
rect 20529 15328 42767 15330
rect 20529 15272 20534 15328
rect 20590 15272 42706 15328
rect 42762 15272 42767 15328
rect 20529 15270 42767 15272
rect 20529 15267 20595 15270
rect 42701 15267 42767 15270
rect 58157 15330 58223 15333
rect 59200 15330 60000 15360
rect 58157 15328 60000 15330
rect 58157 15272 58162 15328
rect 58218 15272 60000 15328
rect 58157 15270 60000 15272
rect 58157 15267 58223 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 59200 15240 60000 15270
rect 50290 15199 50606 15200
rect 32213 15194 32279 15197
rect 35065 15194 35131 15197
rect 32213 15192 35131 15194
rect 32213 15136 32218 15192
rect 32274 15136 35070 15192
rect 35126 15136 35131 15192
rect 32213 15134 35131 15136
rect 32213 15131 32279 15134
rect 35065 15131 35131 15134
rect 38837 15194 38903 15197
rect 40309 15194 40375 15197
rect 38837 15192 40375 15194
rect 38837 15136 38842 15192
rect 38898 15136 40314 15192
rect 40370 15136 40375 15192
rect 38837 15134 40375 15136
rect 38837 15131 38903 15134
rect 40309 15131 40375 15134
rect 11237 15058 11303 15061
rect 15009 15058 15075 15061
rect 11237 15056 15075 15058
rect 11237 15000 11242 15056
rect 11298 15000 15014 15056
rect 15070 15000 15075 15056
rect 11237 14998 15075 15000
rect 11237 14995 11303 14998
rect 15009 14995 15075 14998
rect 30189 15058 30255 15061
rect 36629 15058 36695 15061
rect 30189 15056 36695 15058
rect 30189 15000 30194 15056
rect 30250 15000 36634 15056
rect 36690 15000 36695 15056
rect 30189 14998 36695 15000
rect 30189 14995 30255 14998
rect 36629 14995 36695 14998
rect 38745 15058 38811 15061
rect 46473 15058 46539 15061
rect 38745 15056 46539 15058
rect 38745 15000 38750 15056
rect 38806 15000 46478 15056
rect 46534 15000 46539 15056
rect 38745 14998 46539 15000
rect 38745 14995 38811 14998
rect 46473 14995 46539 14998
rect 0 14922 800 14952
rect 1761 14922 1827 14925
rect 0 14920 1827 14922
rect 0 14864 1766 14920
rect 1822 14864 1827 14920
rect 0 14862 1827 14864
rect 0 14832 800 14862
rect 1761 14859 1827 14862
rect 2405 14922 2471 14925
rect 21030 14922 21036 14924
rect 2405 14920 21036 14922
rect 2405 14864 2410 14920
rect 2466 14864 21036 14920
rect 2405 14862 21036 14864
rect 2405 14859 2471 14862
rect 21030 14860 21036 14862
rect 21100 14860 21106 14924
rect 22093 14922 22159 14925
rect 23565 14922 23631 14925
rect 22093 14920 23631 14922
rect 22093 14864 22098 14920
rect 22154 14864 23570 14920
rect 23626 14864 23631 14920
rect 22093 14862 23631 14864
rect 22093 14859 22159 14862
rect 23565 14859 23631 14862
rect 34053 14922 34119 14925
rect 35525 14922 35591 14925
rect 34053 14920 35591 14922
rect 34053 14864 34058 14920
rect 34114 14864 35530 14920
rect 35586 14864 35591 14920
rect 34053 14862 35591 14864
rect 34053 14859 34119 14862
rect 35525 14859 35591 14862
rect 39113 14922 39179 14925
rect 41413 14922 41479 14925
rect 39113 14920 41479 14922
rect 39113 14864 39118 14920
rect 39174 14864 41418 14920
rect 41474 14864 41479 14920
rect 39113 14862 41479 14864
rect 39113 14859 39179 14862
rect 41413 14859 41479 14862
rect 11789 14786 11855 14789
rect 30741 14786 30807 14789
rect 11789 14784 30807 14786
rect 11789 14728 11794 14784
rect 11850 14728 30746 14784
rect 30802 14728 30807 14784
rect 11789 14726 30807 14728
rect 11789 14723 11855 14726
rect 30741 14723 30807 14726
rect 57973 14786 58039 14789
rect 59200 14786 60000 14816
rect 57973 14784 60000 14786
rect 57973 14728 57978 14784
rect 58034 14728 60000 14784
rect 57973 14726 60000 14728
rect 57973 14723 58039 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 59200 14696 60000 14726
rect 34930 14655 35246 14656
rect 18638 14588 18644 14652
rect 18708 14650 18714 14652
rect 33777 14650 33843 14653
rect 33961 14650 34027 14653
rect 18708 14648 34027 14650
rect 18708 14592 33782 14648
rect 33838 14592 33966 14648
rect 34022 14592 34027 14648
rect 18708 14590 34027 14592
rect 18708 14588 18714 14590
rect 33777 14587 33843 14590
rect 33961 14587 34027 14590
rect 36629 14650 36695 14653
rect 37549 14650 37615 14653
rect 36629 14648 37615 14650
rect 36629 14592 36634 14648
rect 36690 14592 37554 14648
rect 37610 14592 37615 14648
rect 36629 14590 37615 14592
rect 36629 14587 36695 14590
rect 37549 14587 37615 14590
rect 40125 14650 40191 14653
rect 41045 14650 41111 14653
rect 40125 14648 41111 14650
rect 40125 14592 40130 14648
rect 40186 14592 41050 14648
rect 41106 14592 41111 14648
rect 40125 14590 41111 14592
rect 40125 14587 40191 14590
rect 41045 14587 41111 14590
rect 20345 14514 20411 14517
rect 25773 14514 25839 14517
rect 42701 14514 42767 14517
rect 20345 14512 42767 14514
rect 20345 14456 20350 14512
rect 20406 14456 25778 14512
rect 25834 14456 42706 14512
rect 42762 14456 42767 14512
rect 20345 14454 42767 14456
rect 20345 14451 20411 14454
rect 25773 14451 25839 14454
rect 42701 14451 42767 14454
rect 2405 14378 2471 14381
rect 22870 14378 22876 14380
rect 2405 14376 22876 14378
rect 2405 14320 2410 14376
rect 2466 14320 22876 14376
rect 2405 14318 22876 14320
rect 2405 14315 2471 14318
rect 22870 14316 22876 14318
rect 22940 14316 22946 14380
rect 24025 14378 24091 14381
rect 25497 14378 25563 14381
rect 24025 14376 25563 14378
rect 24025 14320 24030 14376
rect 24086 14320 25502 14376
rect 25558 14320 25563 14376
rect 24025 14318 25563 14320
rect 24025 14315 24091 14318
rect 25497 14315 25563 14318
rect 28533 14378 28599 14381
rect 58065 14378 58131 14381
rect 28533 14376 58131 14378
rect 28533 14320 28538 14376
rect 28594 14320 58070 14376
rect 58126 14320 58131 14376
rect 28533 14318 58131 14320
rect 28533 14315 28599 14318
rect 58065 14315 58131 14318
rect 0 14242 800 14272
rect 1853 14242 1919 14245
rect 0 14240 1919 14242
rect 0 14184 1858 14240
rect 1914 14184 1919 14240
rect 0 14182 1919 14184
rect 0 14152 800 14182
rect 1853 14179 1919 14182
rect 13261 14242 13327 14245
rect 15837 14242 15903 14245
rect 19241 14242 19307 14245
rect 13261 14240 19307 14242
rect 13261 14184 13266 14240
rect 13322 14184 15842 14240
rect 15898 14184 19246 14240
rect 19302 14184 19307 14240
rect 13261 14182 19307 14184
rect 13261 14179 13327 14182
rect 15837 14179 15903 14182
rect 19241 14179 19307 14182
rect 24710 14180 24716 14244
rect 24780 14242 24786 14244
rect 39389 14242 39455 14245
rect 24780 14240 39455 14242
rect 24780 14184 39394 14240
rect 39450 14184 39455 14240
rect 24780 14182 39455 14184
rect 24780 14180 24786 14182
rect 39389 14179 39455 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 59200 14152 60000 14272
rect 50290 14111 50606 14112
rect 24117 14106 24183 14109
rect 34237 14106 34303 14109
rect 24117 14104 34303 14106
rect 24117 14048 24122 14104
rect 24178 14048 34242 14104
rect 34298 14048 34303 14104
rect 24117 14046 34303 14048
rect 24117 14043 24183 14046
rect 34237 14043 34303 14046
rect 34513 14106 34579 14109
rect 36905 14106 36971 14109
rect 34513 14104 36971 14106
rect 34513 14048 34518 14104
rect 34574 14048 36910 14104
rect 36966 14048 36971 14104
rect 34513 14046 36971 14048
rect 34513 14043 34579 14046
rect 36905 14043 36971 14046
rect 38745 14106 38811 14109
rect 40585 14106 40651 14109
rect 42333 14106 42399 14109
rect 43345 14106 43411 14109
rect 43805 14106 43871 14109
rect 38745 14104 43871 14106
rect 38745 14048 38750 14104
rect 38806 14048 40590 14104
rect 40646 14048 42338 14104
rect 42394 14048 43350 14104
rect 43406 14048 43810 14104
rect 43866 14048 43871 14104
rect 38745 14046 43871 14048
rect 38745 14043 38811 14046
rect 40585 14043 40651 14046
rect 42333 14043 42399 14046
rect 43345 14043 43411 14046
rect 43805 14043 43871 14046
rect 17861 13970 17927 13973
rect 34697 13970 34763 13973
rect 17861 13968 34763 13970
rect 17861 13912 17866 13968
rect 17922 13912 34702 13968
rect 34758 13912 34763 13968
rect 17861 13910 34763 13912
rect 17861 13907 17927 13910
rect 34697 13907 34763 13910
rect 34881 13970 34947 13973
rect 37181 13970 37247 13973
rect 34881 13968 37247 13970
rect 34881 13912 34886 13968
rect 34942 13912 37186 13968
rect 37242 13912 37247 13968
rect 34881 13910 37247 13912
rect 34881 13907 34947 13910
rect 37181 13907 37247 13910
rect 10225 13834 10291 13837
rect 18045 13834 18111 13837
rect 10225 13832 18111 13834
rect 10225 13776 10230 13832
rect 10286 13776 18050 13832
rect 18106 13776 18111 13832
rect 10225 13774 18111 13776
rect 10225 13771 10291 13774
rect 18045 13771 18111 13774
rect 27245 13834 27311 13837
rect 35566 13834 35572 13836
rect 27245 13832 35572 13834
rect 27245 13776 27250 13832
rect 27306 13776 35572 13832
rect 27245 13774 35572 13776
rect 27245 13771 27311 13774
rect 35566 13772 35572 13774
rect 35636 13834 35642 13836
rect 37641 13834 37707 13837
rect 38193 13834 38259 13837
rect 35636 13832 38259 13834
rect 35636 13776 37646 13832
rect 37702 13776 38198 13832
rect 38254 13776 38259 13832
rect 35636 13774 38259 13776
rect 35636 13772 35642 13774
rect 37641 13771 37707 13774
rect 38193 13771 38259 13774
rect 43846 13772 43852 13836
rect 43916 13834 43922 13836
rect 44081 13834 44147 13837
rect 43916 13832 44147 13834
rect 43916 13776 44086 13832
rect 44142 13776 44147 13832
rect 43916 13774 44147 13776
rect 43916 13772 43922 13774
rect 44081 13771 44147 13774
rect 13537 13698 13603 13701
rect 14365 13698 14431 13701
rect 16205 13698 16271 13701
rect 13537 13696 16271 13698
rect 13537 13640 13542 13696
rect 13598 13640 14370 13696
rect 14426 13640 16210 13696
rect 16266 13640 16271 13696
rect 13537 13638 16271 13640
rect 13537 13635 13603 13638
rect 14365 13635 14431 13638
rect 16205 13635 16271 13638
rect 16982 13636 16988 13700
rect 17052 13698 17058 13700
rect 27102 13698 27108 13700
rect 17052 13638 27108 13698
rect 17052 13636 17058 13638
rect 27102 13636 27108 13638
rect 27172 13636 27178 13700
rect 35433 13698 35499 13701
rect 37733 13698 37799 13701
rect 35433 13696 37799 13698
rect 35433 13640 35438 13696
rect 35494 13640 37738 13696
rect 37794 13640 37799 13696
rect 35433 13638 37799 13640
rect 35433 13635 35499 13638
rect 37733 13635 37799 13638
rect 40309 13698 40375 13701
rect 41597 13698 41663 13701
rect 42149 13698 42215 13701
rect 40309 13696 42215 13698
rect 40309 13640 40314 13696
rect 40370 13640 41602 13696
rect 41658 13640 42154 13696
rect 42210 13640 42215 13696
rect 40309 13638 42215 13640
rect 40309 13635 40375 13638
rect 41597 13635 41663 13638
rect 42149 13635 42215 13638
rect 58157 13698 58223 13701
rect 59200 13698 60000 13728
rect 58157 13696 60000 13698
rect 58157 13640 58162 13696
rect 58218 13640 60000 13696
rect 58157 13638 60000 13640
rect 58157 13635 58223 13638
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 1761 13562 1827 13565
rect 0 13560 1827 13562
rect 0 13504 1766 13560
rect 1822 13504 1827 13560
rect 0 13502 1827 13504
rect 0 13472 800 13502
rect 1761 13499 1827 13502
rect 11421 13562 11487 13565
rect 17401 13562 17467 13565
rect 11421 13560 17467 13562
rect 11421 13504 11426 13560
rect 11482 13504 17406 13560
rect 17462 13504 17467 13560
rect 11421 13502 17467 13504
rect 11421 13499 11487 13502
rect 17401 13499 17467 13502
rect 19374 13500 19380 13564
rect 19444 13562 19450 13564
rect 23749 13562 23815 13565
rect 19444 13560 23815 13562
rect 19444 13504 23754 13560
rect 23810 13504 23815 13560
rect 19444 13502 23815 13504
rect 19444 13500 19450 13502
rect 23749 13499 23815 13502
rect 30097 13562 30163 13565
rect 34278 13562 34284 13564
rect 30097 13560 34284 13562
rect 30097 13504 30102 13560
rect 30158 13504 34284 13560
rect 30097 13502 34284 13504
rect 30097 13499 30163 13502
rect 34278 13500 34284 13502
rect 34348 13500 34354 13564
rect 37089 13562 37155 13565
rect 37222 13562 37228 13564
rect 37089 13560 37228 13562
rect 37089 13504 37094 13560
rect 37150 13504 37228 13560
rect 37089 13502 37228 13504
rect 37089 13499 37155 13502
rect 37222 13500 37228 13502
rect 37292 13500 37298 13564
rect 41137 13562 41203 13565
rect 41094 13560 41203 13562
rect 41094 13504 41142 13560
rect 41198 13504 41203 13560
rect 41094 13499 41203 13504
rect 16021 13426 16087 13429
rect 36813 13426 36879 13429
rect 16021 13424 36879 13426
rect 16021 13368 16026 13424
rect 16082 13368 36818 13424
rect 36874 13368 36879 13424
rect 16021 13366 36879 13368
rect 16021 13363 16087 13366
rect 36813 13363 36879 13366
rect 12341 13290 12407 13293
rect 22829 13290 22895 13293
rect 12341 13288 22895 13290
rect 12341 13232 12346 13288
rect 12402 13232 22834 13288
rect 22890 13232 22895 13288
rect 12341 13230 22895 13232
rect 12341 13227 12407 13230
rect 22829 13227 22895 13230
rect 32397 13290 32463 13293
rect 37733 13290 37799 13293
rect 32397 13288 37799 13290
rect 32397 13232 32402 13288
rect 32458 13232 37738 13288
rect 37794 13232 37799 13288
rect 32397 13230 37799 13232
rect 32397 13227 32463 13230
rect 37733 13227 37799 13230
rect 12985 13154 13051 13157
rect 13537 13154 13603 13157
rect 12985 13152 13603 13154
rect 12985 13096 12990 13152
rect 13046 13096 13542 13152
rect 13598 13096 13603 13152
rect 12985 13094 13603 13096
rect 12985 13091 13051 13094
rect 13537 13091 13603 13094
rect 20805 13154 20871 13157
rect 26509 13154 26575 13157
rect 20805 13152 26575 13154
rect 20805 13096 20810 13152
rect 20866 13096 26514 13152
rect 26570 13096 26575 13152
rect 20805 13094 26575 13096
rect 20805 13091 20871 13094
rect 26509 13091 26575 13094
rect 27521 13154 27587 13157
rect 29729 13154 29795 13157
rect 27521 13152 29795 13154
rect 27521 13096 27526 13152
rect 27582 13096 29734 13152
rect 29790 13096 29795 13152
rect 27521 13094 29795 13096
rect 27521 13091 27587 13094
rect 29729 13091 29795 13094
rect 30005 13154 30071 13157
rect 32581 13154 32647 13157
rect 30005 13152 32647 13154
rect 30005 13096 30010 13152
rect 30066 13096 32586 13152
rect 32642 13096 32647 13152
rect 30005 13094 32647 13096
rect 30005 13091 30071 13094
rect 32581 13091 32647 13094
rect 34973 13154 35039 13157
rect 35801 13154 35867 13157
rect 34973 13152 35867 13154
rect 34973 13096 34978 13152
rect 35034 13096 35806 13152
rect 35862 13096 35867 13152
rect 34973 13094 35867 13096
rect 34973 13091 35039 13094
rect 35801 13091 35867 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 12617 13018 12683 13021
rect 14733 13018 14799 13021
rect 12617 13016 14799 13018
rect 12617 12960 12622 13016
rect 12678 12960 14738 13016
rect 14794 12960 14799 13016
rect 12617 12958 14799 12960
rect 12617 12955 12683 12958
rect 14733 12955 14799 12958
rect 15653 13018 15719 13021
rect 21541 13018 21607 13021
rect 33133 13018 33199 13021
rect 36445 13018 36511 13021
rect 15653 13016 18292 13018
rect 15653 12960 15658 13016
rect 15714 12960 18292 13016
rect 15653 12958 18292 12960
rect 15653 12955 15719 12958
rect 0 12882 800 12912
rect 18232 12885 18292 12958
rect 20118 13016 33199 13018
rect 20118 12960 21546 13016
rect 21602 12960 33138 13016
rect 33194 12960 33199 13016
rect 20118 12958 33199 12960
rect 1853 12882 1919 12885
rect 0 12880 1919 12882
rect 0 12824 1858 12880
rect 1914 12824 1919 12880
rect 0 12822 1919 12824
rect 0 12792 800 12822
rect 1853 12819 1919 12822
rect 10593 12882 10659 12885
rect 17493 12882 17559 12885
rect 10593 12880 17559 12882
rect 10593 12824 10598 12880
rect 10654 12824 17498 12880
rect 17554 12824 17559 12880
rect 10593 12822 17559 12824
rect 10593 12819 10659 12822
rect 17493 12819 17559 12822
rect 18229 12880 18295 12885
rect 18229 12824 18234 12880
rect 18290 12824 18295 12880
rect 18229 12819 18295 12824
rect 18454 12820 18460 12884
rect 18524 12882 18530 12884
rect 20118 12882 20178 12958
rect 21541 12955 21607 12958
rect 33133 12955 33199 12958
rect 34700 13016 36511 13018
rect 34700 12960 36450 13016
rect 36506 12960 36511 13016
rect 34700 12958 36511 12960
rect 18524 12822 20178 12882
rect 21633 12882 21699 12885
rect 24025 12882 24091 12885
rect 32489 12882 32555 12885
rect 21633 12880 24091 12882
rect 21633 12824 21638 12880
rect 21694 12824 24030 12880
rect 24086 12824 24091 12880
rect 21633 12822 24091 12824
rect 18524 12820 18530 12822
rect 21633 12819 21699 12822
rect 24025 12819 24091 12822
rect 26926 12880 32555 12882
rect 26926 12824 32494 12880
rect 32550 12824 32555 12880
rect 26926 12822 32555 12824
rect 11881 12746 11947 12749
rect 12433 12746 12499 12749
rect 14825 12746 14891 12749
rect 18597 12746 18663 12749
rect 11881 12744 18663 12746
rect 11881 12688 11886 12744
rect 11942 12688 12438 12744
rect 12494 12688 14830 12744
rect 14886 12688 18602 12744
rect 18658 12688 18663 12744
rect 11881 12686 18663 12688
rect 11881 12683 11947 12686
rect 12433 12683 12499 12686
rect 14825 12683 14891 12686
rect 18597 12683 18663 12686
rect 19190 12684 19196 12748
rect 19260 12746 19266 12748
rect 26926 12746 26986 12822
rect 32489 12819 32555 12822
rect 33041 12882 33107 12885
rect 34700 12882 34760 12958
rect 36445 12955 36511 12958
rect 33041 12880 34760 12882
rect 33041 12824 33046 12880
rect 33102 12824 34760 12880
rect 33041 12822 34760 12824
rect 35525 12882 35591 12885
rect 38561 12882 38627 12885
rect 41094 12882 41154 13499
rect 57053 13154 57119 13157
rect 59200 13154 60000 13184
rect 57053 13152 60000 13154
rect 57053 13096 57058 13152
rect 57114 13096 60000 13152
rect 57053 13094 60000 13096
rect 57053 13091 57119 13094
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 59200 13064 60000 13094
rect 50290 13023 50606 13024
rect 35525 12880 38627 12882
rect 35525 12824 35530 12880
rect 35586 12824 38566 12880
rect 38622 12824 38627 12880
rect 35525 12822 38627 12824
rect 33041 12819 33107 12822
rect 35525 12819 35591 12822
rect 38561 12819 38627 12822
rect 40358 12822 41154 12882
rect 19260 12686 26986 12746
rect 19260 12684 19266 12686
rect 27102 12684 27108 12748
rect 27172 12746 27178 12748
rect 39941 12746 40007 12749
rect 40358 12746 40418 12822
rect 27172 12744 40418 12746
rect 27172 12688 39946 12744
rect 40002 12688 40418 12744
rect 27172 12686 40418 12688
rect 40493 12746 40559 12749
rect 40493 12744 41154 12746
rect 40493 12688 40498 12744
rect 40554 12688 41154 12744
rect 40493 12686 41154 12688
rect 27172 12684 27178 12686
rect 39941 12683 40007 12686
rect 40493 12683 40559 12686
rect 15653 12610 15719 12613
rect 26969 12610 27035 12613
rect 15653 12608 27035 12610
rect 15653 12552 15658 12608
rect 15714 12552 26974 12608
rect 27030 12552 27035 12608
rect 15653 12550 27035 12552
rect 15653 12547 15719 12550
rect 26969 12547 27035 12550
rect 27153 12610 27219 12613
rect 27797 12610 27863 12613
rect 32673 12610 32739 12613
rect 33593 12612 33659 12613
rect 33542 12610 33548 12612
rect 27153 12608 32739 12610
rect 27153 12552 27158 12608
rect 27214 12552 27802 12608
rect 27858 12552 32678 12608
rect 32734 12552 32739 12608
rect 27153 12550 32739 12552
rect 33502 12550 33548 12610
rect 33612 12608 33659 12612
rect 33654 12552 33659 12608
rect 27153 12547 27219 12550
rect 27797 12547 27863 12550
rect 32673 12547 32739 12550
rect 33542 12548 33548 12550
rect 33612 12548 33659 12552
rect 41094 12610 41154 12686
rect 41229 12610 41295 12613
rect 41094 12608 41295 12610
rect 41094 12552 41234 12608
rect 41290 12552 41295 12608
rect 41094 12550 41295 12552
rect 33593 12547 33659 12548
rect 41229 12547 41295 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 59200 12520 60000 12640
rect 34930 12479 35246 12480
rect 15469 12474 15535 12477
rect 23565 12474 23631 12477
rect 15469 12472 23631 12474
rect 15469 12416 15474 12472
rect 15530 12416 23570 12472
rect 23626 12416 23631 12472
rect 15469 12414 23631 12416
rect 15469 12411 15535 12414
rect 23565 12411 23631 12414
rect 32765 12474 32831 12477
rect 34513 12474 34579 12477
rect 32765 12472 34579 12474
rect 32765 12416 32770 12472
rect 32826 12416 34518 12472
rect 34574 12416 34579 12472
rect 32765 12414 34579 12416
rect 32765 12411 32831 12414
rect 34513 12411 34579 12414
rect 40033 12474 40099 12477
rect 41505 12474 41571 12477
rect 40033 12472 41571 12474
rect 40033 12416 40038 12472
rect 40094 12416 41510 12472
rect 41566 12416 41571 12472
rect 40033 12414 41571 12416
rect 40033 12411 40099 12414
rect 41505 12411 41571 12414
rect 42057 12474 42123 12477
rect 43253 12474 43319 12477
rect 42057 12472 43319 12474
rect 42057 12416 42062 12472
rect 42118 12416 43258 12472
rect 43314 12416 43319 12472
rect 42057 12414 43319 12416
rect 42057 12411 42123 12414
rect 43253 12411 43319 12414
rect 10777 12338 10843 12341
rect 15101 12338 15167 12341
rect 10777 12336 15167 12338
rect 10777 12280 10782 12336
rect 10838 12280 15106 12336
rect 15162 12280 15167 12336
rect 10777 12278 15167 12280
rect 10777 12275 10843 12278
rect 15101 12275 15167 12278
rect 15745 12338 15811 12341
rect 16113 12338 16179 12341
rect 15745 12336 16179 12338
rect 15745 12280 15750 12336
rect 15806 12280 16118 12336
rect 16174 12280 16179 12336
rect 15745 12278 16179 12280
rect 15745 12275 15811 12278
rect 16113 12275 16179 12278
rect 18045 12338 18111 12341
rect 35617 12338 35683 12341
rect 18045 12336 35683 12338
rect 18045 12280 18050 12336
rect 18106 12280 35622 12336
rect 35678 12280 35683 12336
rect 18045 12278 35683 12280
rect 18045 12275 18111 12278
rect 35617 12275 35683 12278
rect 0 12202 800 12232
rect 1853 12202 1919 12205
rect 0 12200 1919 12202
rect 0 12144 1858 12200
rect 1914 12144 1919 12200
rect 0 12142 1919 12144
rect 0 12112 800 12142
rect 1853 12139 1919 12142
rect 11697 12202 11763 12205
rect 30097 12202 30163 12205
rect 33501 12202 33567 12205
rect 11697 12200 33567 12202
rect 11697 12144 11702 12200
rect 11758 12144 30102 12200
rect 30158 12144 33506 12200
rect 33562 12144 33567 12200
rect 11697 12142 33567 12144
rect 11697 12139 11763 12142
rect 30097 12139 30163 12142
rect 33501 12139 33567 12142
rect 34881 12202 34947 12205
rect 37549 12202 37615 12205
rect 34881 12200 37615 12202
rect 34881 12144 34886 12200
rect 34942 12144 37554 12200
rect 37610 12144 37615 12200
rect 34881 12142 37615 12144
rect 34881 12139 34947 12142
rect 37549 12139 37615 12142
rect 12801 12066 12867 12069
rect 16849 12066 16915 12069
rect 12801 12064 16915 12066
rect 12801 12008 12806 12064
rect 12862 12008 16854 12064
rect 16910 12008 16915 12064
rect 12801 12006 16915 12008
rect 12801 12003 12867 12006
rect 16849 12003 16915 12006
rect 24577 12066 24643 12069
rect 25773 12066 25839 12069
rect 40125 12066 40191 12069
rect 24577 12064 24962 12066
rect 24577 12008 24582 12064
rect 24638 12008 24962 12064
rect 24577 12006 24962 12008
rect 24577 12003 24643 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 10685 11930 10751 11933
rect 15009 11930 15075 11933
rect 10685 11928 15075 11930
rect 10685 11872 10690 11928
rect 10746 11872 15014 11928
rect 15070 11872 15075 11928
rect 10685 11870 15075 11872
rect 24902 11930 24962 12006
rect 25773 12064 40191 12066
rect 25773 12008 25778 12064
rect 25834 12008 40130 12064
rect 40186 12008 40191 12064
rect 25773 12006 40191 12008
rect 25773 12003 25839 12006
rect 40125 12003 40191 12006
rect 58157 12066 58223 12069
rect 59200 12066 60000 12096
rect 58157 12064 60000 12066
rect 58157 12008 58162 12064
rect 58218 12008 60000 12064
rect 58157 12006 60000 12008
rect 58157 12003 58223 12006
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 59200 11976 60000 12006
rect 50290 11935 50606 11936
rect 34329 11930 34395 11933
rect 35157 11930 35223 11933
rect 24902 11928 35223 11930
rect 24902 11872 34334 11928
rect 34390 11872 35162 11928
rect 35218 11872 35223 11928
rect 24902 11870 35223 11872
rect 10685 11867 10751 11870
rect 15009 11867 15075 11870
rect 34329 11867 34395 11870
rect 35157 11867 35223 11870
rect 14181 11794 14247 11797
rect 20345 11794 20411 11797
rect 14181 11792 20411 11794
rect 14181 11736 14186 11792
rect 14242 11736 20350 11792
rect 20406 11736 20411 11792
rect 14181 11734 20411 11736
rect 14181 11731 14247 11734
rect 20345 11731 20411 11734
rect 20805 11794 20871 11797
rect 36261 11794 36327 11797
rect 20805 11792 36327 11794
rect 20805 11736 20810 11792
rect 20866 11736 36266 11792
rect 36322 11736 36327 11792
rect 20805 11734 36327 11736
rect 20805 11731 20871 11734
rect 36261 11731 36327 11734
rect 15193 11658 15259 11661
rect 43069 11658 43135 11661
rect 15193 11656 43135 11658
rect 15193 11600 15198 11656
rect 15254 11600 43074 11656
rect 43130 11600 43135 11656
rect 15193 11598 43135 11600
rect 15193 11595 15259 11598
rect 43069 11595 43135 11598
rect 0 11522 800 11552
rect 1761 11522 1827 11525
rect 0 11520 1827 11522
rect 0 11464 1766 11520
rect 1822 11464 1827 11520
rect 0 11462 1827 11464
rect 0 11432 800 11462
rect 1761 11459 1827 11462
rect 15929 11522 15995 11525
rect 16062 11522 16068 11524
rect 15929 11520 16068 11522
rect 15929 11464 15934 11520
rect 15990 11464 16068 11520
rect 15929 11462 16068 11464
rect 15929 11459 15995 11462
rect 16062 11460 16068 11462
rect 16132 11460 16138 11524
rect 17585 11522 17651 11525
rect 20805 11522 20871 11525
rect 17585 11520 20871 11522
rect 17585 11464 17590 11520
rect 17646 11464 20810 11520
rect 20866 11464 20871 11520
rect 17585 11462 20871 11464
rect 17585 11459 17651 11462
rect 20805 11459 20871 11462
rect 21909 11522 21975 11525
rect 25589 11522 25655 11525
rect 21909 11520 25655 11522
rect 21909 11464 21914 11520
rect 21970 11464 25594 11520
rect 25650 11464 25655 11520
rect 21909 11462 25655 11464
rect 21909 11459 21975 11462
rect 25589 11459 25655 11462
rect 29913 11522 29979 11525
rect 32857 11522 32923 11525
rect 34697 11522 34763 11525
rect 29913 11520 32690 11522
rect 29913 11464 29918 11520
rect 29974 11464 32690 11520
rect 29913 11462 32690 11464
rect 29913 11459 29979 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 11605 11386 11671 11389
rect 16941 11386 17007 11389
rect 11605 11384 17007 11386
rect 11605 11328 11610 11384
rect 11666 11328 16946 11384
rect 17002 11328 17007 11384
rect 11605 11326 17007 11328
rect 11605 11323 11671 11326
rect 16941 11323 17007 11326
rect 18873 11386 18939 11389
rect 32630 11386 32690 11462
rect 32857 11520 34763 11522
rect 32857 11464 32862 11520
rect 32918 11464 34702 11520
rect 34758 11464 34763 11520
rect 32857 11462 34763 11464
rect 32857 11459 32923 11462
rect 34697 11459 34763 11462
rect 36077 11522 36143 11525
rect 38561 11522 38627 11525
rect 36077 11520 38627 11522
rect 36077 11464 36082 11520
rect 36138 11464 38566 11520
rect 38622 11464 38627 11520
rect 36077 11462 38627 11464
rect 36077 11459 36143 11462
rect 38561 11459 38627 11462
rect 40677 11522 40743 11525
rect 46749 11522 46815 11525
rect 40677 11520 46815 11522
rect 40677 11464 40682 11520
rect 40738 11464 46754 11520
rect 46810 11464 46815 11520
rect 40677 11462 46815 11464
rect 40677 11459 40743 11462
rect 46749 11459 46815 11462
rect 58065 11522 58131 11525
rect 59200 11522 60000 11552
rect 58065 11520 60000 11522
rect 58065 11464 58070 11520
rect 58126 11464 60000 11520
rect 58065 11462 60000 11464
rect 58065 11459 58131 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 59200 11432 60000 11462
rect 34930 11391 35246 11392
rect 34053 11386 34119 11389
rect 18873 11384 31770 11386
rect 18873 11328 18878 11384
rect 18934 11328 31770 11384
rect 18873 11326 31770 11328
rect 32630 11384 34119 11386
rect 32630 11328 34058 11384
rect 34114 11328 34119 11384
rect 32630 11326 34119 11328
rect 18873 11323 18939 11326
rect 13353 11250 13419 11253
rect 17033 11250 17099 11253
rect 13353 11248 17099 11250
rect 13353 11192 13358 11248
rect 13414 11192 17038 11248
rect 17094 11192 17099 11248
rect 13353 11190 17099 11192
rect 13353 11187 13419 11190
rect 17033 11187 17099 11190
rect 17309 11250 17375 11253
rect 23841 11250 23907 11253
rect 17309 11248 23907 11250
rect 17309 11192 17314 11248
rect 17370 11192 23846 11248
rect 23902 11192 23907 11248
rect 17309 11190 23907 11192
rect 31710 11250 31770 11326
rect 34053 11323 34119 11326
rect 34462 11324 34468 11388
rect 34532 11386 34538 11388
rect 34605 11386 34671 11389
rect 34532 11384 34671 11386
rect 34532 11328 34610 11384
rect 34666 11328 34671 11384
rect 34532 11326 34671 11328
rect 34532 11324 34538 11326
rect 34605 11323 34671 11326
rect 36261 11386 36327 11389
rect 37365 11386 37431 11389
rect 36261 11384 37431 11386
rect 36261 11328 36266 11384
rect 36322 11328 37370 11384
rect 37426 11328 37431 11384
rect 36261 11326 37431 11328
rect 36261 11323 36327 11326
rect 37365 11323 37431 11326
rect 40350 11324 40356 11388
rect 40420 11386 40426 11388
rect 40861 11386 40927 11389
rect 40420 11384 40927 11386
rect 40420 11328 40866 11384
rect 40922 11328 40927 11384
rect 40420 11326 40927 11328
rect 40420 11324 40426 11326
rect 40861 11323 40927 11326
rect 36629 11250 36695 11253
rect 31710 11248 36695 11250
rect 31710 11192 36634 11248
rect 36690 11192 36695 11248
rect 31710 11190 36695 11192
rect 17309 11187 17375 11190
rect 23841 11187 23907 11190
rect 36629 11187 36695 11190
rect 43621 11250 43687 11253
rect 44081 11250 44147 11253
rect 43621 11248 44147 11250
rect 43621 11192 43626 11248
rect 43682 11192 44086 11248
rect 44142 11192 44147 11248
rect 43621 11190 44147 11192
rect 43621 11187 43687 11190
rect 44081 11187 44147 11190
rect 13261 11114 13327 11117
rect 16665 11114 16731 11117
rect 13261 11112 16731 11114
rect 13261 11056 13266 11112
rect 13322 11056 16670 11112
rect 16726 11056 16731 11112
rect 13261 11054 16731 11056
rect 13261 11051 13327 11054
rect 16665 11051 16731 11054
rect 17401 11114 17467 11117
rect 21265 11114 21331 11117
rect 17401 11112 21331 11114
rect 17401 11056 17406 11112
rect 17462 11056 21270 11112
rect 21326 11056 21331 11112
rect 17401 11054 21331 11056
rect 17401 11051 17467 11054
rect 21265 11051 21331 11054
rect 21909 11114 21975 11117
rect 22185 11114 22251 11117
rect 21909 11112 22251 11114
rect 21909 11056 21914 11112
rect 21970 11056 22190 11112
rect 22246 11056 22251 11112
rect 21909 11054 22251 11056
rect 21909 11051 21975 11054
rect 22185 11051 22251 11054
rect 29913 11114 29979 11117
rect 33317 11114 33383 11117
rect 29913 11112 33383 11114
rect 29913 11056 29918 11112
rect 29974 11056 33322 11112
rect 33378 11056 33383 11112
rect 29913 11054 33383 11056
rect 29913 11051 29979 11054
rect 33317 11051 33383 11054
rect 34237 11114 34303 11117
rect 35525 11114 35591 11117
rect 34237 11112 35591 11114
rect 34237 11056 34242 11112
rect 34298 11056 35530 11112
rect 35586 11056 35591 11112
rect 34237 11054 35591 11056
rect 34237 11051 34303 11054
rect 35525 11051 35591 11054
rect 35801 11114 35867 11117
rect 36169 11114 36235 11117
rect 35801 11112 36235 11114
rect 35801 11056 35806 11112
rect 35862 11056 36174 11112
rect 36230 11056 36235 11112
rect 35801 11054 36235 11056
rect 35801 11051 35867 11054
rect 36169 11051 36235 11054
rect 39246 11052 39252 11116
rect 39316 11114 39322 11116
rect 40166 11114 40172 11116
rect 39316 11054 40172 11114
rect 39316 11052 39322 11054
rect 40166 11052 40172 11054
rect 40236 11052 40242 11116
rect 50613 11114 50679 11117
rect 53005 11114 53071 11117
rect 50613 11112 53071 11114
rect 50613 11056 50618 11112
rect 50674 11056 53010 11112
rect 53066 11056 53071 11112
rect 50613 11054 53071 11056
rect 50613 11051 50679 11054
rect 53005 11051 53071 11054
rect 14549 10978 14615 10981
rect 17217 10978 17283 10981
rect 14549 10976 17283 10978
rect 14549 10920 14554 10976
rect 14610 10920 17222 10976
rect 17278 10920 17283 10976
rect 14549 10918 17283 10920
rect 14549 10915 14615 10918
rect 17217 10915 17283 10918
rect 17902 10916 17908 10980
rect 17972 10978 17978 10980
rect 18321 10978 18387 10981
rect 17972 10976 18387 10978
rect 17972 10920 18326 10976
rect 18382 10920 18387 10976
rect 17972 10918 18387 10920
rect 17972 10916 17978 10918
rect 18321 10915 18387 10918
rect 20345 10978 20411 10981
rect 20805 10978 20871 10981
rect 20345 10976 20871 10978
rect 20345 10920 20350 10976
rect 20406 10920 20810 10976
rect 20866 10920 20871 10976
rect 20345 10918 20871 10920
rect 20345 10915 20411 10918
rect 20805 10915 20871 10918
rect 21541 10978 21607 10981
rect 23657 10978 23723 10981
rect 21541 10976 23723 10978
rect 21541 10920 21546 10976
rect 21602 10920 23662 10976
rect 23718 10920 23723 10976
rect 21541 10918 23723 10920
rect 21541 10915 21607 10918
rect 23657 10915 23723 10918
rect 25957 10978 26023 10981
rect 33685 10978 33751 10981
rect 36077 10978 36143 10981
rect 25957 10976 36143 10978
rect 25957 10920 25962 10976
rect 26018 10920 33690 10976
rect 33746 10920 36082 10976
rect 36138 10920 36143 10976
rect 25957 10918 36143 10920
rect 25957 10915 26023 10918
rect 33685 10915 33751 10918
rect 36077 10915 36143 10918
rect 36302 10916 36308 10980
rect 36372 10978 36378 10980
rect 36629 10978 36695 10981
rect 36372 10976 36695 10978
rect 36372 10920 36634 10976
rect 36690 10920 36695 10976
rect 36372 10918 36695 10920
rect 36372 10916 36378 10918
rect 36629 10915 36695 10918
rect 38101 10978 38167 10981
rect 38653 10978 38719 10981
rect 38101 10976 38719 10978
rect 38101 10920 38106 10976
rect 38162 10920 38658 10976
rect 38714 10920 38719 10976
rect 38101 10918 38719 10920
rect 38101 10915 38167 10918
rect 38653 10915 38719 10918
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 60000 11008
rect 50290 10847 50606 10848
rect 1853 10842 1919 10845
rect 0 10840 1919 10842
rect 0 10784 1858 10840
rect 1914 10784 1919 10840
rect 0 10782 1919 10784
rect 0 10752 800 10782
rect 1853 10779 1919 10782
rect 12617 10842 12683 10845
rect 18597 10842 18663 10845
rect 12617 10840 18663 10842
rect 12617 10784 12622 10840
rect 12678 10784 18602 10840
rect 18658 10784 18663 10840
rect 12617 10782 18663 10784
rect 12617 10779 12683 10782
rect 18597 10779 18663 10782
rect 20437 10842 20503 10845
rect 26693 10842 26759 10845
rect 20437 10840 26759 10842
rect 20437 10784 20442 10840
rect 20498 10784 26698 10840
rect 26754 10784 26759 10840
rect 20437 10782 26759 10784
rect 20437 10779 20503 10782
rect 26693 10779 26759 10782
rect 30005 10842 30071 10845
rect 31293 10842 31359 10845
rect 48957 10842 49023 10845
rect 30005 10840 49023 10842
rect 30005 10784 30010 10840
rect 30066 10784 31298 10840
rect 31354 10784 48962 10840
rect 49018 10784 49023 10840
rect 30005 10782 49023 10784
rect 30005 10779 30071 10782
rect 31293 10779 31359 10782
rect 48957 10779 49023 10782
rect 1577 10706 1643 10709
rect 19241 10706 19307 10709
rect 21909 10706 21975 10709
rect 22185 10708 22251 10709
rect 22134 10706 22140 10708
rect 1577 10704 12450 10706
rect 1577 10648 1582 10704
rect 1638 10648 12450 10704
rect 1577 10646 12450 10648
rect 1577 10643 1643 10646
rect 12390 10434 12450 10646
rect 19241 10704 21975 10706
rect 19241 10648 19246 10704
rect 19302 10648 21914 10704
rect 21970 10648 21975 10704
rect 19241 10646 21975 10648
rect 22094 10646 22140 10706
rect 22204 10704 22251 10708
rect 22246 10648 22251 10704
rect 19241 10643 19307 10646
rect 21909 10643 21975 10646
rect 22134 10644 22140 10646
rect 22204 10644 22251 10648
rect 22185 10643 22251 10644
rect 22369 10706 22435 10709
rect 24025 10706 24091 10709
rect 22369 10704 24091 10706
rect 22369 10648 22374 10704
rect 22430 10648 24030 10704
rect 24086 10648 24091 10704
rect 22369 10646 24091 10648
rect 22369 10643 22435 10646
rect 24025 10643 24091 10646
rect 32581 10706 32647 10709
rect 42609 10706 42675 10709
rect 32581 10704 42675 10706
rect 32581 10648 32586 10704
rect 32642 10648 42614 10704
rect 42670 10648 42675 10704
rect 32581 10646 42675 10648
rect 32581 10643 32647 10646
rect 42609 10643 42675 10646
rect 15745 10570 15811 10573
rect 41505 10570 41571 10573
rect 15745 10568 41571 10570
rect 15745 10512 15750 10568
rect 15806 10512 41510 10568
rect 41566 10512 41571 10568
rect 15745 10510 41571 10512
rect 15745 10507 15811 10510
rect 41505 10507 41571 10510
rect 28809 10434 28875 10437
rect 12390 10432 28875 10434
rect 12390 10376 28814 10432
rect 28870 10376 28875 10432
rect 12390 10374 28875 10376
rect 28809 10371 28875 10374
rect 32857 10434 32923 10437
rect 34053 10434 34119 10437
rect 34697 10436 34763 10437
rect 34646 10434 34652 10436
rect 32857 10432 34119 10434
rect 32857 10376 32862 10432
rect 32918 10376 34058 10432
rect 34114 10376 34119 10432
rect 32857 10374 34119 10376
rect 34606 10374 34652 10434
rect 34716 10432 34763 10436
rect 34758 10376 34763 10432
rect 32857 10371 32923 10374
rect 34053 10371 34119 10374
rect 34646 10372 34652 10374
rect 34716 10372 34763 10376
rect 34697 10371 34763 10372
rect 35525 10434 35591 10437
rect 38101 10434 38167 10437
rect 35525 10432 38167 10434
rect 35525 10376 35530 10432
rect 35586 10376 38106 10432
rect 38162 10376 38167 10432
rect 35525 10374 38167 10376
rect 35525 10371 35591 10374
rect 38101 10371 38167 10374
rect 40677 10436 40743 10437
rect 40677 10432 40724 10436
rect 40788 10434 40794 10436
rect 57881 10434 57947 10437
rect 59200 10434 60000 10464
rect 40677 10376 40682 10432
rect 40677 10372 40724 10376
rect 40788 10374 40834 10434
rect 57881 10432 60000 10434
rect 57881 10376 57886 10432
rect 57942 10376 60000 10432
rect 57881 10374 60000 10376
rect 40788 10372 40794 10374
rect 40677 10371 40743 10372
rect 57881 10371 57947 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 59200 10344 60000 10374
rect 34930 10303 35246 10304
rect 16849 10298 16915 10301
rect 24117 10298 24183 10301
rect 16849 10296 24183 10298
rect 16849 10240 16854 10296
rect 16910 10240 24122 10296
rect 24178 10240 24183 10296
rect 16849 10238 24183 10240
rect 16849 10235 16915 10238
rect 24117 10235 24183 10238
rect 27613 10298 27679 10301
rect 33961 10298 34027 10301
rect 34329 10298 34395 10301
rect 27613 10296 34395 10298
rect 27613 10240 27618 10296
rect 27674 10240 33966 10296
rect 34022 10240 34334 10296
rect 34390 10240 34395 10296
rect 27613 10238 34395 10240
rect 27613 10235 27679 10238
rect 33961 10235 34027 10238
rect 34329 10235 34395 10238
rect 34462 10236 34468 10300
rect 34532 10298 34538 10300
rect 34789 10298 34855 10301
rect 34532 10296 34855 10298
rect 34532 10240 34794 10296
rect 34850 10240 34855 10296
rect 34532 10238 34855 10240
rect 34532 10236 34538 10238
rect 34789 10235 34855 10238
rect 35709 10298 35775 10301
rect 38745 10298 38811 10301
rect 35709 10296 38811 10298
rect 35709 10240 35714 10296
rect 35770 10240 38750 10296
rect 38806 10240 38811 10296
rect 35709 10238 38811 10240
rect 35709 10235 35775 10238
rect 38745 10235 38811 10238
rect 39982 10236 39988 10300
rect 40052 10298 40058 10300
rect 51809 10298 51875 10301
rect 40052 10296 51875 10298
rect 40052 10240 51814 10296
rect 51870 10240 51875 10296
rect 40052 10238 51875 10240
rect 40052 10236 40058 10238
rect 51809 10235 51875 10238
rect 0 10162 800 10192
rect 1761 10162 1827 10165
rect 0 10160 1827 10162
rect 0 10104 1766 10160
rect 1822 10104 1827 10160
rect 0 10102 1827 10104
rect 0 10072 800 10102
rect 1761 10099 1827 10102
rect 15101 10162 15167 10165
rect 16941 10162 17007 10165
rect 15101 10160 17007 10162
rect 15101 10104 15106 10160
rect 15162 10104 16946 10160
rect 17002 10104 17007 10160
rect 15101 10102 17007 10104
rect 15101 10099 15167 10102
rect 16941 10099 17007 10102
rect 17493 10162 17559 10165
rect 31845 10162 31911 10165
rect 37549 10162 37615 10165
rect 17493 10160 31770 10162
rect 17493 10104 17498 10160
rect 17554 10104 31770 10160
rect 17493 10102 31770 10104
rect 17493 10099 17559 10102
rect 19425 10028 19491 10029
rect 19374 9964 19380 10028
rect 19444 10026 19491 10028
rect 19793 10026 19859 10029
rect 20110 10026 20116 10028
rect 19444 10024 19536 10026
rect 19486 9968 19536 10024
rect 19444 9966 19536 9968
rect 19793 10024 20116 10026
rect 19793 9968 19798 10024
rect 19854 9968 20116 10024
rect 19793 9966 20116 9968
rect 19444 9964 19491 9966
rect 19425 9963 19491 9964
rect 19793 9963 19859 9966
rect 20110 9964 20116 9966
rect 20180 9964 20186 10028
rect 22318 9964 22324 10028
rect 22388 10026 22394 10028
rect 23657 10026 23723 10029
rect 22388 10024 23723 10026
rect 22388 9968 23662 10024
rect 23718 9968 23723 10024
rect 22388 9966 23723 9968
rect 22388 9964 22394 9966
rect 23657 9963 23723 9966
rect 24669 10026 24735 10029
rect 26693 10026 26759 10029
rect 24669 10024 26759 10026
rect 24669 9968 24674 10024
rect 24730 9968 26698 10024
rect 26754 9968 26759 10024
rect 24669 9966 26759 9968
rect 31710 10026 31770 10102
rect 31845 10160 37615 10162
rect 31845 10104 31850 10160
rect 31906 10104 37554 10160
rect 37610 10104 37615 10160
rect 31845 10102 37615 10104
rect 31845 10099 31911 10102
rect 37549 10099 37615 10102
rect 40309 10026 40375 10029
rect 31710 10024 40375 10026
rect 31710 9968 40314 10024
rect 40370 9968 40375 10024
rect 31710 9966 40375 9968
rect 24669 9963 24735 9966
rect 26693 9963 26759 9966
rect 40309 9963 40375 9966
rect 16113 9890 16179 9893
rect 18689 9890 18755 9893
rect 16113 9888 18755 9890
rect 16113 9832 16118 9888
rect 16174 9832 18694 9888
rect 18750 9832 18755 9888
rect 16113 9830 18755 9832
rect 16113 9827 16179 9830
rect 18689 9827 18755 9830
rect 20437 9890 20503 9893
rect 23974 9890 23980 9892
rect 20437 9888 23980 9890
rect 20437 9832 20442 9888
rect 20498 9832 23980 9888
rect 20437 9830 23980 9832
rect 20437 9827 20503 9830
rect 23974 9828 23980 9830
rect 24044 9890 24050 9892
rect 24669 9890 24735 9893
rect 24044 9888 24735 9890
rect 24044 9832 24674 9888
rect 24730 9832 24735 9888
rect 24044 9830 24735 9832
rect 24044 9828 24050 9830
rect 24669 9827 24735 9830
rect 34053 9890 34119 9893
rect 35249 9890 35315 9893
rect 34053 9888 35315 9890
rect 34053 9832 34058 9888
rect 34114 9832 35254 9888
rect 35310 9832 35315 9888
rect 34053 9830 35315 9832
rect 34053 9827 34119 9830
rect 35249 9827 35315 9830
rect 35433 9890 35499 9893
rect 35985 9890 36051 9893
rect 35433 9888 36051 9890
rect 35433 9832 35438 9888
rect 35494 9832 35990 9888
rect 36046 9832 36051 9888
rect 35433 9830 36051 9832
rect 35433 9827 35499 9830
rect 35985 9827 36051 9830
rect 36169 9890 36235 9893
rect 36905 9890 36971 9893
rect 36169 9888 36971 9890
rect 36169 9832 36174 9888
rect 36230 9832 36910 9888
rect 36966 9832 36971 9888
rect 36169 9830 36971 9832
rect 36169 9827 36235 9830
rect 36905 9827 36971 9830
rect 58065 9890 58131 9893
rect 59200 9890 60000 9920
rect 58065 9888 60000 9890
rect 58065 9832 58070 9888
rect 58126 9832 60000 9888
rect 58065 9830 60000 9832
rect 58065 9827 58131 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 59200 9800 60000 9830
rect 50290 9759 50606 9760
rect 15837 9754 15903 9757
rect 18413 9754 18479 9757
rect 18873 9754 18939 9757
rect 15837 9752 18939 9754
rect 15837 9696 15842 9752
rect 15898 9696 18418 9752
rect 18474 9696 18878 9752
rect 18934 9696 18939 9752
rect 15837 9694 18939 9696
rect 15837 9691 15903 9694
rect 18413 9691 18479 9694
rect 18873 9691 18939 9694
rect 20713 9754 20779 9757
rect 26417 9754 26483 9757
rect 27889 9754 27955 9757
rect 20713 9752 27955 9754
rect 20713 9696 20718 9752
rect 20774 9696 26422 9752
rect 26478 9696 27894 9752
rect 27950 9696 27955 9752
rect 20713 9694 27955 9696
rect 20713 9691 20779 9694
rect 26417 9691 26483 9694
rect 27889 9691 27955 9694
rect 30097 9754 30163 9757
rect 32673 9754 32739 9757
rect 30097 9752 32739 9754
rect 30097 9696 30102 9752
rect 30158 9696 32678 9752
rect 32734 9696 32739 9752
rect 30097 9694 32739 9696
rect 30097 9691 30163 9694
rect 32673 9691 32739 9694
rect 33501 9754 33567 9757
rect 38009 9754 38075 9757
rect 33501 9752 38075 9754
rect 33501 9696 33506 9752
rect 33562 9696 38014 9752
rect 38070 9696 38075 9752
rect 33501 9694 38075 9696
rect 33501 9691 33567 9694
rect 38009 9691 38075 9694
rect 38929 9754 38995 9757
rect 39573 9754 39639 9757
rect 38929 9752 39639 9754
rect 38929 9696 38934 9752
rect 38990 9696 39578 9752
rect 39634 9696 39639 9752
rect 38929 9694 39639 9696
rect 38929 9691 38995 9694
rect 39573 9691 39639 9694
rect 39798 9692 39804 9756
rect 39868 9754 39874 9756
rect 40217 9754 40283 9757
rect 39868 9752 40283 9754
rect 39868 9696 40222 9752
rect 40278 9696 40283 9752
rect 39868 9694 40283 9696
rect 39868 9692 39874 9694
rect 40217 9691 40283 9694
rect 1577 9618 1643 9621
rect 31201 9618 31267 9621
rect 1577 9616 31267 9618
rect 1577 9560 1582 9616
rect 1638 9560 31206 9616
rect 31262 9560 31267 9616
rect 1577 9558 31267 9560
rect 1577 9555 1643 9558
rect 31201 9555 31267 9558
rect 31569 9618 31635 9621
rect 32949 9618 33015 9621
rect 31569 9616 33015 9618
rect 31569 9560 31574 9616
rect 31630 9560 32954 9616
rect 33010 9560 33015 9616
rect 31569 9558 33015 9560
rect 31569 9555 31635 9558
rect 32949 9555 33015 9558
rect 33542 9556 33548 9620
rect 33612 9618 33618 9620
rect 34053 9618 34119 9621
rect 33612 9616 34119 9618
rect 33612 9560 34058 9616
rect 34114 9560 34119 9616
rect 33612 9558 34119 9560
rect 33612 9556 33618 9558
rect 34053 9555 34119 9558
rect 34237 9620 34303 9621
rect 34237 9616 34284 9620
rect 34348 9618 34354 9620
rect 34237 9560 34242 9616
rect 34237 9556 34284 9560
rect 34348 9558 34394 9618
rect 34348 9556 34354 9558
rect 34462 9556 34468 9620
rect 34532 9618 34538 9620
rect 34973 9618 35039 9621
rect 35382 9618 35388 9620
rect 34532 9616 35388 9618
rect 34532 9560 34978 9616
rect 35034 9560 35388 9616
rect 34532 9558 35388 9560
rect 34532 9556 34538 9558
rect 34237 9555 34303 9556
rect 34973 9555 35039 9558
rect 35382 9556 35388 9558
rect 35452 9556 35458 9620
rect 35801 9618 35867 9621
rect 36118 9618 36124 9620
rect 35801 9616 36124 9618
rect 35801 9560 35806 9616
rect 35862 9560 36124 9616
rect 35801 9558 36124 9560
rect 35801 9555 35867 9558
rect 36118 9556 36124 9558
rect 36188 9556 36194 9620
rect 38377 9618 38443 9621
rect 38510 9618 38516 9620
rect 38377 9616 38516 9618
rect 38377 9560 38382 9616
rect 38438 9560 38516 9616
rect 38377 9558 38516 9560
rect 38377 9555 38443 9558
rect 38510 9556 38516 9558
rect 38580 9556 38586 9620
rect 39757 9618 39823 9621
rect 45921 9618 45987 9621
rect 39757 9616 45987 9618
rect 39757 9560 39762 9616
rect 39818 9560 45926 9616
rect 45982 9560 45987 9616
rect 39757 9558 45987 9560
rect 39757 9555 39823 9558
rect 45921 9555 45987 9558
rect 0 9482 800 9512
rect 1761 9482 1827 9485
rect 0 9480 1827 9482
rect 0 9424 1766 9480
rect 1822 9424 1827 9480
rect 0 9422 1827 9424
rect 0 9392 800 9422
rect 1761 9419 1827 9422
rect 16062 9420 16068 9484
rect 16132 9482 16138 9484
rect 16941 9482 17007 9485
rect 16132 9480 17007 9482
rect 16132 9424 16946 9480
rect 17002 9424 17007 9480
rect 16132 9422 17007 9424
rect 16132 9420 16138 9422
rect 16941 9419 17007 9422
rect 19793 9482 19859 9485
rect 20294 9482 20300 9484
rect 19793 9480 20300 9482
rect 19793 9424 19798 9480
rect 19854 9424 20300 9480
rect 19793 9422 20300 9424
rect 19793 9419 19859 9422
rect 20294 9420 20300 9422
rect 20364 9420 20370 9484
rect 20621 9482 20687 9485
rect 20846 9482 20852 9484
rect 20621 9480 20852 9482
rect 20621 9424 20626 9480
rect 20682 9424 20852 9480
rect 20621 9422 20852 9424
rect 20621 9419 20687 9422
rect 20846 9420 20852 9422
rect 20916 9420 20922 9484
rect 25773 9482 25839 9485
rect 22050 9480 25839 9482
rect 22050 9424 25778 9480
rect 25834 9424 25839 9480
rect 22050 9422 25839 9424
rect 14457 9346 14523 9349
rect 17401 9346 17467 9349
rect 14457 9344 17467 9346
rect 14457 9288 14462 9344
rect 14518 9288 17406 9344
rect 17462 9288 17467 9344
rect 14457 9286 17467 9288
rect 14457 9283 14523 9286
rect 17401 9283 17467 9286
rect 18505 9346 18571 9349
rect 22050 9346 22110 9422
rect 25773 9419 25839 9422
rect 28901 9482 28967 9485
rect 36077 9482 36143 9485
rect 28901 9480 36143 9482
rect 28901 9424 28906 9480
rect 28962 9424 36082 9480
rect 36138 9424 36143 9480
rect 28901 9422 36143 9424
rect 28901 9419 28967 9422
rect 36077 9419 36143 9422
rect 38653 9484 38719 9485
rect 38653 9480 38700 9484
rect 38764 9482 38770 9484
rect 38653 9424 38658 9480
rect 38653 9420 38700 9424
rect 38764 9422 38810 9482
rect 38764 9420 38770 9422
rect 38653 9419 38719 9420
rect 18505 9344 22110 9346
rect 18505 9288 18510 9344
rect 18566 9288 22110 9344
rect 18505 9286 22110 9288
rect 22921 9346 22987 9349
rect 23054 9346 23060 9348
rect 22921 9344 23060 9346
rect 22921 9288 22926 9344
rect 22982 9288 23060 9344
rect 22921 9286 23060 9288
rect 18505 9283 18571 9286
rect 22921 9283 22987 9286
rect 23054 9284 23060 9286
rect 23124 9284 23130 9348
rect 23657 9346 23723 9349
rect 29913 9346 29979 9349
rect 23657 9344 29979 9346
rect 23657 9288 23662 9344
rect 23718 9288 29918 9344
rect 29974 9288 29979 9344
rect 23657 9286 29979 9288
rect 23657 9283 23723 9286
rect 29913 9283 29979 9286
rect 30097 9346 30163 9349
rect 33409 9346 33475 9349
rect 33961 9346 34027 9349
rect 30097 9344 31954 9346
rect 30097 9288 30102 9344
rect 30158 9288 31954 9344
rect 30097 9286 31954 9288
rect 30097 9283 30163 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 17401 9212 17467 9213
rect 17350 9148 17356 9212
rect 17420 9210 17467 9212
rect 18781 9210 18847 9213
rect 20621 9210 20687 9213
rect 26049 9210 26115 9213
rect 17420 9208 17512 9210
rect 17462 9152 17512 9208
rect 17420 9150 17512 9152
rect 18781 9208 26115 9210
rect 18781 9152 18786 9208
rect 18842 9152 20626 9208
rect 20682 9152 26054 9208
rect 26110 9152 26115 9208
rect 18781 9150 26115 9152
rect 17420 9148 17467 9150
rect 17401 9147 17467 9148
rect 18781 9147 18847 9150
rect 20621 9147 20687 9150
rect 26049 9147 26115 9150
rect 29453 9210 29519 9213
rect 30741 9210 30807 9213
rect 31753 9210 31819 9213
rect 29453 9208 29930 9210
rect 29453 9152 29458 9208
rect 29514 9152 29930 9208
rect 29453 9150 29930 9152
rect 29453 9147 29519 9150
rect 13629 9074 13695 9077
rect 27429 9074 27495 9077
rect 13629 9072 27495 9074
rect 13629 9016 13634 9072
rect 13690 9016 27434 9072
rect 27490 9016 27495 9072
rect 13629 9014 27495 9016
rect 13629 9011 13695 9014
rect 27429 9011 27495 9014
rect 29453 9074 29519 9077
rect 29637 9074 29703 9077
rect 29453 9072 29703 9074
rect 29453 9016 29458 9072
rect 29514 9016 29642 9072
rect 29698 9016 29703 9072
rect 29453 9014 29703 9016
rect 29870 9074 29930 9150
rect 30741 9208 31819 9210
rect 30741 9152 30746 9208
rect 30802 9152 31758 9208
rect 31814 9152 31819 9208
rect 30741 9150 31819 9152
rect 31894 9210 31954 9286
rect 33409 9344 34027 9346
rect 33409 9288 33414 9344
rect 33470 9288 33966 9344
rect 34022 9288 34027 9344
rect 33409 9286 34027 9288
rect 33409 9283 33475 9286
rect 33961 9283 34027 9286
rect 34462 9284 34468 9348
rect 34532 9346 34538 9348
rect 34605 9346 34671 9349
rect 34532 9344 34671 9346
rect 34532 9288 34610 9344
rect 34666 9288 34671 9344
rect 34532 9286 34671 9288
rect 34532 9284 34538 9286
rect 34605 9283 34671 9286
rect 34789 9344 34855 9349
rect 34789 9288 34794 9344
rect 34850 9288 34855 9344
rect 34789 9283 34855 9288
rect 35617 9346 35683 9349
rect 35985 9346 36051 9349
rect 37181 9346 37247 9349
rect 35617 9344 35910 9346
rect 35617 9288 35622 9344
rect 35678 9288 35910 9344
rect 35617 9286 35910 9288
rect 35617 9283 35683 9286
rect 34792 9210 34852 9283
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 31894 9150 34852 9210
rect 35850 9210 35910 9286
rect 35985 9344 37247 9346
rect 35985 9288 35990 9344
rect 36046 9288 37186 9344
rect 37242 9288 37247 9344
rect 35985 9286 37247 9288
rect 35985 9283 36051 9286
rect 37181 9283 37247 9286
rect 39665 9346 39731 9349
rect 40125 9346 40191 9349
rect 39665 9344 40191 9346
rect 39665 9288 39670 9344
rect 39726 9288 40130 9344
rect 40186 9288 40191 9344
rect 39665 9286 40191 9288
rect 39665 9283 39731 9286
rect 40125 9283 40191 9286
rect 59200 9256 60000 9376
rect 36537 9210 36603 9213
rect 35850 9208 36603 9210
rect 35850 9152 36542 9208
rect 36598 9152 36603 9208
rect 35850 9150 36603 9152
rect 30741 9147 30807 9150
rect 31753 9147 31819 9150
rect 36537 9147 36603 9150
rect 39573 9210 39639 9213
rect 44265 9210 44331 9213
rect 39573 9208 44331 9210
rect 39573 9152 39578 9208
rect 39634 9152 44270 9208
rect 44326 9152 44331 9208
rect 39573 9150 44331 9152
rect 39573 9147 39639 9150
rect 44265 9147 44331 9150
rect 33317 9074 33383 9077
rect 42609 9074 42675 9077
rect 29870 9072 42675 9074
rect 29870 9016 33322 9072
rect 33378 9016 42614 9072
rect 42670 9016 42675 9072
rect 29870 9014 42675 9016
rect 29453 9011 29519 9014
rect 29637 9011 29703 9014
rect 33317 9011 33383 9014
rect 42609 9011 42675 9014
rect 16205 8938 16271 8941
rect 16430 8938 16436 8940
rect 16205 8936 16436 8938
rect 16205 8880 16210 8936
rect 16266 8880 16436 8936
rect 16205 8878 16436 8880
rect 16205 8875 16271 8878
rect 16430 8876 16436 8878
rect 16500 8876 16506 8940
rect 17953 8938 18019 8941
rect 19057 8938 19123 8941
rect 17953 8936 19123 8938
rect 17953 8880 17958 8936
rect 18014 8880 19062 8936
rect 19118 8880 19123 8936
rect 17953 8878 19123 8880
rect 17953 8875 18019 8878
rect 19057 8875 19123 8878
rect 19701 8938 19767 8941
rect 32949 8938 33015 8941
rect 55397 8938 55463 8941
rect 19701 8936 20500 8938
rect 19701 8880 19706 8936
rect 19762 8880 20500 8936
rect 19701 8878 20500 8880
rect 19701 8875 19767 8878
rect 0 8802 800 8832
rect 20440 8805 20500 8878
rect 20670 8878 31770 8938
rect 1853 8802 1919 8805
rect 0 8800 1919 8802
rect 0 8744 1858 8800
rect 1914 8744 1919 8800
rect 0 8742 1919 8744
rect 0 8712 800 8742
rect 1853 8739 1919 8742
rect 16297 8802 16363 8805
rect 18965 8802 19031 8805
rect 16297 8800 19031 8802
rect 16297 8744 16302 8800
rect 16358 8744 18970 8800
rect 19026 8744 19031 8800
rect 16297 8742 19031 8744
rect 16297 8739 16363 8742
rect 18965 8739 19031 8742
rect 20437 8800 20503 8805
rect 20437 8744 20442 8800
rect 20498 8744 20503 8800
rect 20437 8739 20503 8744
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 19977 8666 20043 8669
rect 20110 8666 20116 8668
rect 19977 8664 20116 8666
rect 19977 8608 19982 8664
rect 20038 8608 20116 8664
rect 19977 8606 20116 8608
rect 19977 8603 20043 8606
rect 20110 8604 20116 8606
rect 20180 8604 20186 8668
rect 17677 8530 17743 8533
rect 20670 8530 20730 8878
rect 22093 8802 22159 8805
rect 22369 8802 22435 8805
rect 23289 8802 23355 8805
rect 24209 8802 24275 8805
rect 31569 8802 31635 8805
rect 22093 8800 23355 8802
rect 22093 8744 22098 8800
rect 22154 8744 22374 8800
rect 22430 8744 23294 8800
rect 23350 8744 23355 8800
rect 22093 8742 23355 8744
rect 22093 8739 22159 8742
rect 22369 8739 22435 8742
rect 23289 8739 23355 8742
rect 23430 8800 31635 8802
rect 23430 8744 24214 8800
rect 24270 8744 31574 8800
rect 31630 8744 31635 8800
rect 23430 8742 31635 8744
rect 31710 8802 31770 8878
rect 32949 8936 55463 8938
rect 32949 8880 32954 8936
rect 33010 8880 55402 8936
rect 55458 8880 55463 8936
rect 32949 8878 55463 8880
rect 32949 8875 33015 8878
rect 55397 8875 55463 8878
rect 40861 8802 40927 8805
rect 41229 8802 41295 8805
rect 31710 8800 41295 8802
rect 31710 8744 40866 8800
rect 40922 8744 41234 8800
rect 41290 8744 41295 8800
rect 31710 8742 41295 8744
rect 21081 8666 21147 8669
rect 23430 8666 23490 8742
rect 24209 8739 24275 8742
rect 31569 8739 31635 8742
rect 40861 8739 40927 8742
rect 41229 8739 41295 8742
rect 58157 8802 58223 8805
rect 59200 8802 60000 8832
rect 58157 8800 60000 8802
rect 58157 8744 58162 8800
rect 58218 8744 60000 8800
rect 58157 8742 60000 8744
rect 58157 8739 58223 8742
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 59200 8712 60000 8742
rect 50290 8671 50606 8672
rect 21081 8664 23490 8666
rect 21081 8608 21086 8664
rect 21142 8608 23490 8664
rect 21081 8606 23490 8608
rect 23749 8666 23815 8669
rect 26969 8666 27035 8669
rect 34237 8666 34303 8669
rect 23749 8664 24042 8666
rect 23749 8608 23754 8664
rect 23810 8608 24042 8664
rect 23749 8606 24042 8608
rect 21081 8603 21147 8606
rect 23749 8603 23815 8606
rect 23749 8532 23815 8533
rect 23749 8530 23796 8532
rect 17677 8528 20730 8530
rect 17677 8472 17682 8528
rect 17738 8472 20730 8528
rect 17677 8470 20730 8472
rect 23704 8528 23796 8530
rect 23704 8472 23754 8528
rect 23704 8470 23796 8472
rect 17677 8467 17743 8470
rect 23749 8468 23796 8470
rect 23860 8468 23866 8532
rect 23982 8530 24042 8606
rect 26969 8664 34303 8666
rect 26969 8608 26974 8664
rect 27030 8608 34242 8664
rect 34298 8608 34303 8664
rect 26969 8606 34303 8608
rect 26969 8603 27035 8606
rect 34237 8603 34303 8606
rect 34513 8666 34579 8669
rect 35249 8666 35315 8669
rect 34513 8664 35315 8666
rect 34513 8608 34518 8664
rect 34574 8608 35254 8664
rect 35310 8608 35315 8664
rect 34513 8606 35315 8608
rect 34513 8603 34579 8606
rect 35249 8603 35315 8606
rect 35382 8604 35388 8668
rect 35452 8666 35458 8668
rect 38929 8666 38995 8669
rect 35452 8664 38995 8666
rect 35452 8608 38934 8664
rect 38990 8608 38995 8664
rect 35452 8606 38995 8608
rect 35452 8604 35458 8606
rect 38929 8603 38995 8606
rect 24393 8530 24459 8533
rect 32121 8530 32187 8533
rect 23982 8528 32187 8530
rect 23982 8472 24398 8528
rect 24454 8472 32126 8528
rect 32182 8472 32187 8528
rect 23982 8470 32187 8472
rect 23749 8467 23815 8468
rect 24393 8467 24459 8470
rect 32121 8467 32187 8470
rect 34881 8530 34947 8533
rect 35341 8530 35407 8533
rect 35566 8530 35572 8532
rect 34881 8528 35572 8530
rect 34881 8472 34886 8528
rect 34942 8472 35346 8528
rect 35402 8472 35572 8528
rect 34881 8470 35572 8472
rect 34881 8467 34947 8470
rect 35341 8467 35407 8470
rect 35566 8468 35572 8470
rect 35636 8468 35642 8532
rect 36670 8468 36676 8532
rect 36740 8530 36746 8532
rect 36905 8530 36971 8533
rect 36740 8528 36971 8530
rect 36740 8472 36910 8528
rect 36966 8472 36971 8528
rect 36740 8470 36971 8472
rect 36740 8468 36746 8470
rect 36905 8467 36971 8470
rect 39665 8530 39731 8533
rect 40493 8530 40559 8533
rect 39665 8528 40559 8530
rect 39665 8472 39670 8528
rect 39726 8472 40498 8528
rect 40554 8472 40559 8528
rect 39665 8470 40559 8472
rect 39665 8467 39731 8470
rect 40493 8467 40559 8470
rect 18229 8394 18295 8397
rect 19057 8394 19123 8397
rect 18229 8392 19123 8394
rect 18229 8336 18234 8392
rect 18290 8336 19062 8392
rect 19118 8336 19123 8392
rect 18229 8334 19123 8336
rect 18229 8331 18295 8334
rect 19057 8331 19123 8334
rect 19333 8394 19399 8397
rect 19977 8394 20043 8397
rect 19333 8392 20043 8394
rect 19333 8336 19338 8392
rect 19394 8336 19982 8392
rect 20038 8336 20043 8392
rect 19333 8334 20043 8336
rect 19333 8331 19399 8334
rect 19977 8331 20043 8334
rect 20253 8394 20319 8397
rect 22318 8394 22324 8396
rect 20253 8392 22324 8394
rect 20253 8336 20258 8392
rect 20314 8336 22324 8392
rect 20253 8334 22324 8336
rect 20253 8331 20319 8334
rect 22318 8332 22324 8334
rect 22388 8332 22394 8396
rect 22553 8394 22619 8397
rect 23289 8394 23355 8397
rect 28901 8394 28967 8397
rect 22553 8392 28967 8394
rect 22553 8336 22558 8392
rect 22614 8336 23294 8392
rect 23350 8336 28906 8392
rect 28962 8336 28967 8392
rect 22553 8334 28967 8336
rect 22553 8331 22619 8334
rect 23289 8331 23355 8334
rect 28901 8331 28967 8334
rect 31937 8394 32003 8397
rect 33542 8394 33548 8396
rect 31937 8392 33548 8394
rect 31937 8336 31942 8392
rect 31998 8336 33548 8392
rect 31937 8334 33548 8336
rect 31937 8331 32003 8334
rect 33542 8332 33548 8334
rect 33612 8332 33618 8396
rect 33726 8332 33732 8396
rect 33796 8394 33802 8396
rect 40677 8394 40743 8397
rect 33796 8334 35450 8394
rect 33796 8332 33802 8334
rect 11881 8258 11947 8261
rect 30097 8258 30163 8261
rect 33869 8260 33935 8261
rect 34605 8260 34671 8261
rect 30230 8258 30236 8260
rect 11881 8256 26986 8258
rect 11881 8200 11886 8256
rect 11942 8200 26986 8256
rect 11881 8198 26986 8200
rect 11881 8195 11947 8198
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 1761 8122 1827 8125
rect 0 8120 1827 8122
rect 0 8064 1766 8120
rect 1822 8064 1827 8120
rect 0 8062 1827 8064
rect 0 8032 800 8062
rect 1761 8059 1827 8062
rect 18597 8122 18663 8125
rect 19149 8122 19215 8125
rect 20529 8122 20595 8125
rect 22553 8122 22619 8125
rect 23238 8122 23244 8124
rect 18597 8120 22110 8122
rect 18597 8064 18602 8120
rect 18658 8064 19154 8120
rect 19210 8064 20534 8120
rect 20590 8064 22110 8120
rect 18597 8062 22110 8064
rect 18597 8059 18663 8062
rect 19149 8059 19215 8062
rect 20529 8059 20595 8062
rect 12934 7924 12940 7988
rect 13004 7986 13010 7988
rect 18413 7986 18479 7989
rect 13004 7984 18479 7986
rect 13004 7928 18418 7984
rect 18474 7928 18479 7984
rect 13004 7926 18479 7928
rect 13004 7924 13010 7926
rect 18413 7923 18479 7926
rect 19793 7986 19859 7989
rect 20253 7986 20319 7989
rect 21909 7986 21975 7989
rect 19793 7984 20178 7986
rect 19793 7928 19798 7984
rect 19854 7928 20178 7984
rect 19793 7926 20178 7928
rect 19793 7923 19859 7926
rect 10317 7850 10383 7853
rect 13077 7850 13143 7853
rect 20118 7850 20178 7926
rect 20253 7984 21975 7986
rect 20253 7928 20258 7984
rect 20314 7928 21914 7984
rect 21970 7928 21975 7984
rect 20253 7926 21975 7928
rect 22050 7986 22110 8062
rect 22553 8120 23244 8122
rect 22553 8064 22558 8120
rect 22614 8064 23244 8120
rect 22553 8062 23244 8064
rect 22553 8059 22619 8062
rect 23238 8060 23244 8062
rect 23308 8060 23314 8124
rect 26926 8122 26986 8198
rect 30097 8256 30236 8258
rect 30097 8200 30102 8256
rect 30158 8200 30236 8256
rect 30097 8198 30236 8200
rect 30097 8195 30163 8198
rect 30230 8196 30236 8198
rect 30300 8196 30306 8260
rect 33869 8258 33916 8260
rect 33824 8256 33916 8258
rect 33824 8200 33874 8256
rect 33824 8198 33916 8200
rect 33869 8196 33916 8198
rect 33980 8196 33986 8260
rect 34605 8258 34652 8260
rect 34560 8256 34652 8258
rect 34560 8200 34610 8256
rect 34560 8198 34652 8200
rect 34605 8196 34652 8198
rect 34716 8196 34722 8260
rect 35390 8258 35450 8334
rect 35942 8392 40743 8394
rect 35942 8336 40682 8392
rect 40738 8336 40743 8392
rect 35942 8334 40743 8336
rect 35942 8258 36002 8334
rect 40677 8331 40743 8334
rect 35390 8198 36002 8258
rect 36353 8258 36419 8261
rect 37273 8258 37339 8261
rect 36353 8256 37339 8258
rect 36353 8200 36358 8256
rect 36414 8200 37278 8256
rect 37334 8200 37339 8256
rect 36353 8198 37339 8200
rect 33869 8195 33935 8196
rect 34605 8195 34671 8196
rect 36353 8195 36419 8198
rect 37273 8195 37339 8198
rect 38193 8258 38259 8261
rect 38561 8258 38627 8261
rect 38193 8256 38627 8258
rect 38193 8200 38198 8256
rect 38254 8200 38566 8256
rect 38622 8200 38627 8256
rect 38193 8198 38627 8200
rect 38193 8195 38259 8198
rect 38561 8195 38627 8198
rect 39757 8258 39823 8261
rect 39982 8258 39988 8260
rect 39757 8256 39988 8258
rect 39757 8200 39762 8256
rect 39818 8200 39988 8256
rect 39757 8198 39988 8200
rect 39757 8195 39823 8198
rect 39982 8196 39988 8198
rect 40052 8196 40058 8260
rect 40166 8196 40172 8260
rect 40236 8258 40242 8260
rect 40861 8258 40927 8261
rect 40236 8256 40927 8258
rect 40236 8200 40866 8256
rect 40922 8200 40927 8256
rect 40236 8198 40927 8200
rect 40236 8196 40242 8198
rect 40861 8195 40927 8198
rect 57145 8258 57211 8261
rect 59200 8258 60000 8288
rect 57145 8256 60000 8258
rect 57145 8200 57150 8256
rect 57206 8200 60000 8256
rect 57145 8198 60000 8200
rect 57145 8195 57211 8198
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 31661 8122 31727 8125
rect 26926 8120 31727 8122
rect 26926 8064 31666 8120
rect 31722 8064 31727 8120
rect 26926 8062 31727 8064
rect 31661 8059 31727 8062
rect 35801 8122 35867 8125
rect 49693 8122 49759 8125
rect 35801 8120 49759 8122
rect 35801 8064 35806 8120
rect 35862 8064 49698 8120
rect 49754 8064 49759 8120
rect 35801 8062 49759 8064
rect 35801 8059 35867 8062
rect 49693 8059 49759 8062
rect 25129 7986 25195 7989
rect 38469 7986 38535 7989
rect 38745 7988 38811 7989
rect 22050 7984 38535 7986
rect 22050 7928 25134 7984
rect 25190 7928 38474 7984
rect 38530 7928 38535 7984
rect 22050 7926 38535 7928
rect 20253 7923 20319 7926
rect 21909 7923 21975 7926
rect 25129 7923 25195 7926
rect 38469 7923 38535 7926
rect 38694 7924 38700 7988
rect 38764 7986 38811 7988
rect 40033 7986 40099 7989
rect 44541 7986 44607 7989
rect 38764 7984 38856 7986
rect 38806 7928 38856 7984
rect 38764 7926 38856 7928
rect 40033 7984 44607 7986
rect 40033 7928 40038 7984
rect 40094 7928 44546 7984
rect 44602 7928 44607 7984
rect 40033 7926 44607 7928
rect 38764 7924 38811 7926
rect 38745 7923 38811 7924
rect 40033 7923 40099 7926
rect 44541 7923 44607 7926
rect 20805 7850 20871 7853
rect 10317 7848 18844 7850
rect 10317 7792 10322 7848
rect 10378 7792 13082 7848
rect 13138 7792 18844 7848
rect 10317 7790 18844 7792
rect 20118 7848 20871 7850
rect 20118 7792 20810 7848
rect 20866 7792 20871 7848
rect 20118 7790 20871 7792
rect 10317 7787 10383 7790
rect 13077 7787 13143 7790
rect 18784 7717 18844 7790
rect 20805 7787 20871 7790
rect 23105 7850 23171 7853
rect 39113 7850 39179 7853
rect 23105 7848 39179 7850
rect 23105 7792 23110 7848
rect 23166 7792 39118 7848
rect 39174 7792 39179 7848
rect 23105 7790 39179 7792
rect 23105 7787 23171 7790
rect 39113 7787 39179 7790
rect 13721 7714 13787 7717
rect 14406 7714 14412 7716
rect 13721 7712 14412 7714
rect 13721 7656 13726 7712
rect 13782 7656 14412 7712
rect 13721 7654 14412 7656
rect 13721 7651 13787 7654
rect 14406 7652 14412 7654
rect 14476 7652 14482 7716
rect 14733 7714 14799 7717
rect 16982 7714 16988 7716
rect 14733 7712 16988 7714
rect 14733 7656 14738 7712
rect 14794 7656 16988 7712
rect 14733 7654 16988 7656
rect 14733 7651 14799 7654
rect 16982 7652 16988 7654
rect 17052 7652 17058 7716
rect 18781 7714 18847 7717
rect 19149 7714 19215 7717
rect 22277 7714 22343 7717
rect 18781 7712 19215 7714
rect 18781 7656 18786 7712
rect 18842 7656 19154 7712
rect 19210 7656 19215 7712
rect 18781 7654 19215 7656
rect 18781 7651 18847 7654
rect 19149 7651 19215 7654
rect 19980 7712 22343 7714
rect 19980 7656 22282 7712
rect 22338 7656 22343 7712
rect 19980 7654 22343 7656
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 19980 7581 20040 7654
rect 22277 7651 22343 7654
rect 27981 7714 28047 7717
rect 30281 7714 30347 7717
rect 27981 7712 30347 7714
rect 27981 7656 27986 7712
rect 28042 7656 30286 7712
rect 30342 7656 30347 7712
rect 27981 7654 30347 7656
rect 27981 7651 28047 7654
rect 30281 7651 30347 7654
rect 31109 7714 31175 7717
rect 42241 7714 42307 7717
rect 31109 7712 42307 7714
rect 31109 7656 31114 7712
rect 31170 7656 42246 7712
rect 42302 7656 42307 7712
rect 31109 7654 42307 7656
rect 31109 7651 31175 7654
rect 42241 7651 42307 7654
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 59200 7624 60000 7744
rect 50290 7583 50606 7584
rect 19425 7580 19491 7581
rect 19374 7578 19380 7580
rect 19334 7518 19380 7578
rect 19444 7576 19491 7580
rect 19486 7520 19491 7576
rect 19374 7516 19380 7518
rect 19444 7516 19491 7520
rect 19425 7515 19491 7516
rect 19977 7576 20043 7581
rect 19977 7520 19982 7576
rect 20038 7520 20043 7576
rect 19977 7515 20043 7520
rect 20897 7578 20963 7581
rect 21449 7578 21515 7581
rect 22001 7580 22067 7581
rect 21950 7578 21956 7580
rect 20897 7576 21515 7578
rect 20897 7520 20902 7576
rect 20958 7520 21454 7576
rect 21510 7520 21515 7576
rect 20897 7518 21515 7520
rect 21910 7518 21956 7578
rect 22020 7576 22067 7580
rect 22062 7520 22067 7576
rect 20897 7515 20963 7518
rect 21449 7515 21515 7518
rect 21950 7516 21956 7518
rect 22020 7516 22067 7520
rect 22001 7515 22067 7516
rect 33961 7578 34027 7581
rect 41229 7578 41295 7581
rect 33961 7576 41295 7578
rect 33961 7520 33966 7576
rect 34022 7520 41234 7576
rect 41290 7520 41295 7576
rect 33961 7518 41295 7520
rect 33961 7515 34027 7518
rect 41229 7515 41295 7518
rect 0 7442 800 7472
rect 1853 7442 1919 7445
rect 0 7440 1919 7442
rect 0 7384 1858 7440
rect 1914 7384 1919 7440
rect 0 7382 1919 7384
rect 0 7352 800 7382
rect 1853 7379 1919 7382
rect 15653 7442 15719 7445
rect 35249 7442 35315 7445
rect 39205 7442 39271 7445
rect 15653 7440 39271 7442
rect 15653 7384 15658 7440
rect 15714 7384 35254 7440
rect 35310 7384 39210 7440
rect 39266 7384 39271 7440
rect 15653 7382 39271 7384
rect 15653 7379 15719 7382
rect 35249 7379 35315 7382
rect 39205 7379 39271 7382
rect 9397 7306 9463 7309
rect 25773 7306 25839 7309
rect 9397 7304 25839 7306
rect 9397 7248 9402 7304
rect 9458 7248 25778 7304
rect 25834 7248 25839 7304
rect 9397 7246 25839 7248
rect 9397 7243 9463 7246
rect 25773 7243 25839 7246
rect 32397 7306 32463 7309
rect 36353 7306 36419 7309
rect 32397 7304 36419 7306
rect 32397 7248 32402 7304
rect 32458 7248 36358 7304
rect 36414 7248 36419 7304
rect 32397 7246 36419 7248
rect 32397 7243 32463 7246
rect 36353 7243 36419 7246
rect 38837 7306 38903 7309
rect 39113 7306 39179 7309
rect 38837 7304 39179 7306
rect 38837 7248 38842 7304
rect 38898 7248 39118 7304
rect 39174 7248 39179 7304
rect 38837 7246 39179 7248
rect 38837 7243 38903 7246
rect 39113 7243 39179 7246
rect 13905 7170 13971 7173
rect 21541 7170 21607 7173
rect 13905 7168 21607 7170
rect 13905 7112 13910 7168
rect 13966 7112 21546 7168
rect 21602 7112 21607 7168
rect 13905 7110 21607 7112
rect 13905 7107 13971 7110
rect 21541 7107 21607 7110
rect 27521 7170 27587 7173
rect 34145 7170 34211 7173
rect 27521 7168 34211 7170
rect 27521 7112 27526 7168
rect 27582 7112 34150 7168
rect 34206 7112 34211 7168
rect 27521 7110 34211 7112
rect 27521 7107 27587 7110
rect 34145 7107 34211 7110
rect 35341 7170 35407 7173
rect 35801 7170 35867 7173
rect 35341 7168 35867 7170
rect 35341 7112 35346 7168
rect 35402 7112 35806 7168
rect 35862 7112 35867 7168
rect 35341 7110 35867 7112
rect 35341 7107 35407 7110
rect 35801 7107 35867 7110
rect 36537 7170 36603 7173
rect 38469 7170 38535 7173
rect 36537 7168 38535 7170
rect 36537 7112 36542 7168
rect 36598 7112 38474 7168
rect 38530 7112 38535 7168
rect 36537 7110 38535 7112
rect 36537 7107 36603 7110
rect 38469 7107 38535 7110
rect 57329 7170 57395 7173
rect 59200 7170 60000 7200
rect 57329 7168 60000 7170
rect 57329 7112 57334 7168
rect 57390 7112 60000 7168
rect 57329 7110 60000 7112
rect 57329 7107 57395 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 59200 7080 60000 7110
rect 34930 7039 35246 7040
rect 13997 7034 14063 7037
rect 34605 7034 34671 7037
rect 37641 7034 37707 7037
rect 13997 7032 34671 7034
rect 13997 6976 14002 7032
rect 14058 6976 34610 7032
rect 34666 6976 34671 7032
rect 13997 6974 34671 6976
rect 13997 6971 14063 6974
rect 34605 6971 34671 6974
rect 35390 7032 37707 7034
rect 35390 6976 37646 7032
rect 37702 6976 37707 7032
rect 35390 6974 37707 6976
rect 18413 6900 18479 6901
rect 18413 6896 18460 6900
rect 18524 6898 18530 6900
rect 20253 6898 20319 6901
rect 20713 6898 20779 6901
rect 20846 6898 20852 6900
rect 18413 6840 18418 6896
rect 18413 6836 18460 6840
rect 18524 6838 18570 6898
rect 20253 6896 20852 6898
rect 20253 6840 20258 6896
rect 20314 6840 20718 6896
rect 20774 6840 20852 6896
rect 20253 6838 20852 6840
rect 18524 6836 18530 6838
rect 18413 6835 18479 6836
rect 20253 6835 20319 6838
rect 20713 6835 20779 6838
rect 20846 6836 20852 6838
rect 20916 6836 20922 6900
rect 22318 6836 22324 6900
rect 22388 6898 22394 6900
rect 22461 6898 22527 6901
rect 22388 6896 22527 6898
rect 22388 6840 22466 6896
rect 22522 6840 22527 6896
rect 22388 6838 22527 6840
rect 22388 6836 22394 6838
rect 22461 6835 22527 6838
rect 23473 6898 23539 6901
rect 27521 6898 27587 6901
rect 23473 6896 27587 6898
rect 23473 6840 23478 6896
rect 23534 6840 27526 6896
rect 27582 6840 27587 6896
rect 23473 6838 27587 6840
rect 23473 6835 23539 6838
rect 27521 6835 27587 6838
rect 29729 6898 29795 6901
rect 31109 6900 31175 6901
rect 29862 6898 29868 6900
rect 29729 6896 29868 6898
rect 29729 6840 29734 6896
rect 29790 6840 29868 6896
rect 29729 6838 29868 6840
rect 29729 6835 29795 6838
rect 29862 6836 29868 6838
rect 29932 6836 29938 6900
rect 31109 6898 31156 6900
rect 31064 6896 31156 6898
rect 31064 6840 31114 6896
rect 31064 6838 31156 6840
rect 31109 6836 31156 6838
rect 31220 6836 31226 6900
rect 32673 6898 32739 6901
rect 32806 6898 32812 6900
rect 32673 6896 32812 6898
rect 32673 6840 32678 6896
rect 32734 6840 32812 6896
rect 32673 6838 32812 6840
rect 31109 6835 31175 6836
rect 32673 6835 32739 6838
rect 32806 6836 32812 6838
rect 32876 6836 32882 6900
rect 33225 6898 33291 6901
rect 34697 6898 34763 6901
rect 33225 6896 34763 6898
rect 33225 6840 33230 6896
rect 33286 6840 34702 6896
rect 34758 6840 34763 6896
rect 33225 6838 34763 6840
rect 33225 6835 33291 6838
rect 34697 6835 34763 6838
rect 34881 6898 34947 6901
rect 35390 6898 35450 6974
rect 37641 6971 37707 6974
rect 34881 6896 35450 6898
rect 34881 6840 34886 6896
rect 34942 6840 35450 6896
rect 34881 6838 35450 6840
rect 35525 6898 35591 6901
rect 37549 6898 37615 6901
rect 35525 6896 37615 6898
rect 35525 6840 35530 6896
rect 35586 6840 37554 6896
rect 37610 6840 37615 6896
rect 35525 6838 37615 6840
rect 34881 6835 34947 6838
rect 35525 6835 35591 6838
rect 37549 6835 37615 6838
rect 43805 6900 43871 6901
rect 43805 6896 43852 6900
rect 43916 6898 43922 6900
rect 43805 6840 43810 6896
rect 43805 6836 43852 6840
rect 43916 6838 43962 6898
rect 43916 6836 43922 6838
rect 43805 6835 43871 6836
rect 0 6762 800 6792
rect 1853 6762 1919 6765
rect 0 6760 1919 6762
rect 0 6704 1858 6760
rect 1914 6704 1919 6760
rect 0 6702 1919 6704
rect 0 6672 800 6702
rect 1853 6699 1919 6702
rect 17217 6762 17283 6765
rect 22093 6762 22159 6765
rect 17217 6760 22159 6762
rect 17217 6704 17222 6760
rect 17278 6704 22098 6760
rect 22154 6704 22159 6760
rect 17217 6702 22159 6704
rect 17217 6699 17283 6702
rect 22093 6699 22159 6702
rect 23013 6762 23079 6765
rect 51257 6762 51323 6765
rect 23013 6760 51323 6762
rect 23013 6704 23018 6760
rect 23074 6704 51262 6760
rect 51318 6704 51323 6760
rect 23013 6702 51323 6704
rect 23013 6699 23079 6702
rect 51257 6699 51323 6702
rect 18321 6626 18387 6629
rect 19057 6626 19123 6629
rect 18321 6624 19123 6626
rect 18321 6568 18326 6624
rect 18382 6568 19062 6624
rect 19118 6568 19123 6624
rect 18321 6566 19123 6568
rect 18321 6563 18387 6566
rect 19057 6563 19123 6566
rect 24945 6626 25011 6629
rect 31201 6626 31267 6629
rect 36169 6626 36235 6629
rect 24945 6624 36235 6626
rect 24945 6568 24950 6624
rect 25006 6568 31206 6624
rect 31262 6568 36174 6624
rect 36230 6568 36235 6624
rect 24945 6566 36235 6568
rect 24945 6563 25011 6566
rect 31201 6563 31267 6566
rect 36169 6563 36235 6566
rect 36997 6626 37063 6629
rect 38193 6626 38259 6629
rect 36997 6624 38259 6626
rect 36997 6568 37002 6624
rect 37058 6568 38198 6624
rect 38254 6568 38259 6624
rect 36997 6566 38259 6568
rect 36997 6563 37063 6566
rect 38193 6563 38259 6566
rect 58065 6626 58131 6629
rect 59200 6626 60000 6656
rect 58065 6624 60000 6626
rect 58065 6568 58070 6624
rect 58126 6568 60000 6624
rect 58065 6566 60000 6568
rect 58065 6563 58131 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 59200 6536 60000 6566
rect 50290 6495 50606 6496
rect 14917 6490 14983 6493
rect 19333 6492 19399 6493
rect 19190 6490 19196 6492
rect 14917 6488 19196 6490
rect 14917 6432 14922 6488
rect 14978 6432 19196 6488
rect 14917 6430 19196 6432
rect 14917 6427 14983 6430
rect 19190 6428 19196 6430
rect 19260 6428 19266 6492
rect 19333 6488 19380 6492
rect 19444 6490 19450 6492
rect 22461 6490 22527 6493
rect 32581 6490 32647 6493
rect 19333 6432 19338 6488
rect 19333 6428 19380 6432
rect 19444 6430 19490 6490
rect 19980 6488 31770 6490
rect 19980 6432 22466 6488
rect 22522 6432 31770 6488
rect 19980 6430 31770 6432
rect 19444 6428 19450 6430
rect 19333 6427 19399 6428
rect 18229 6354 18295 6357
rect 19241 6354 19307 6357
rect 18229 6352 19307 6354
rect 18229 6296 18234 6352
rect 18290 6296 19246 6352
rect 19302 6296 19307 6352
rect 18229 6294 19307 6296
rect 18229 6291 18295 6294
rect 19241 6291 19307 6294
rect 19374 6292 19380 6356
rect 19444 6354 19450 6356
rect 19980 6354 20040 6430
rect 22461 6427 22527 6430
rect 19444 6294 20040 6354
rect 20437 6354 20503 6357
rect 23289 6354 23355 6357
rect 29177 6354 29243 6357
rect 20437 6352 23355 6354
rect 20437 6296 20442 6352
rect 20498 6296 23294 6352
rect 23350 6296 23355 6352
rect 20437 6294 23355 6296
rect 19444 6292 19450 6294
rect 20437 6291 20503 6294
rect 23289 6291 23355 6294
rect 26926 6352 29243 6354
rect 26926 6296 29182 6352
rect 29238 6296 29243 6352
rect 26926 6294 29243 6296
rect 31710 6354 31770 6430
rect 32581 6488 41430 6490
rect 32581 6432 32586 6488
rect 32642 6432 41430 6488
rect 32581 6430 41430 6432
rect 32581 6427 32647 6430
rect 39665 6354 39731 6357
rect 31710 6352 39731 6354
rect 31710 6296 39670 6352
rect 39726 6296 39731 6352
rect 31710 6294 39731 6296
rect 17493 6218 17559 6221
rect 26926 6218 26986 6294
rect 29177 6291 29243 6294
rect 39665 6291 39731 6294
rect 17493 6216 26986 6218
rect 17493 6160 17498 6216
rect 17554 6160 26986 6216
rect 17493 6158 26986 6160
rect 30097 6218 30163 6221
rect 37365 6218 37431 6221
rect 30097 6216 37431 6218
rect 30097 6160 30102 6216
rect 30158 6160 37370 6216
rect 37426 6160 37431 6216
rect 30097 6158 37431 6160
rect 41370 6218 41430 6430
rect 55213 6218 55279 6221
rect 41370 6216 55279 6218
rect 41370 6160 55218 6216
rect 55274 6160 55279 6216
rect 41370 6158 55279 6160
rect 17493 6155 17559 6158
rect 30097 6155 30163 6158
rect 37365 6155 37431 6158
rect 55213 6155 55279 6158
rect 0 6082 800 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 800 6022
rect 1761 6019 1827 6022
rect 21909 6082 21975 6085
rect 22093 6082 22159 6085
rect 21909 6080 22159 6082
rect 21909 6024 21914 6080
rect 21970 6024 22098 6080
rect 22154 6024 22159 6080
rect 21909 6022 22159 6024
rect 21909 6019 21975 6022
rect 22093 6019 22159 6022
rect 23381 6082 23447 6085
rect 31017 6082 31083 6085
rect 23381 6080 31083 6082
rect 23381 6024 23386 6080
rect 23442 6024 31022 6080
rect 31078 6024 31083 6080
rect 23381 6022 31083 6024
rect 23381 6019 23447 6022
rect 31017 6019 31083 6022
rect 33317 6082 33383 6085
rect 34605 6082 34671 6085
rect 33317 6080 34671 6082
rect 33317 6024 33322 6080
rect 33378 6024 34610 6080
rect 34666 6024 34671 6080
rect 33317 6022 34671 6024
rect 33317 6019 33383 6022
rect 34605 6019 34671 6022
rect 35525 6082 35591 6085
rect 36905 6082 36971 6085
rect 35525 6080 36971 6082
rect 35525 6024 35530 6080
rect 35586 6024 36910 6080
rect 36966 6024 36971 6080
rect 35525 6022 36971 6024
rect 35525 6019 35591 6022
rect 36905 6019 36971 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 59200 5992 60000 6112
rect 34930 5951 35246 5952
rect 17585 5946 17651 5949
rect 22829 5946 22895 5949
rect 17585 5944 22895 5946
rect 17585 5888 17590 5944
rect 17646 5888 22834 5944
rect 22890 5888 22895 5944
rect 17585 5886 22895 5888
rect 17585 5883 17651 5886
rect 22829 5883 22895 5886
rect 24485 5946 24551 5949
rect 27337 5946 27403 5949
rect 24485 5944 27403 5946
rect 24485 5888 24490 5944
rect 24546 5888 27342 5944
rect 27398 5888 27403 5944
rect 24485 5886 27403 5888
rect 24485 5883 24551 5886
rect 27337 5883 27403 5886
rect 30005 5946 30071 5949
rect 30649 5946 30715 5949
rect 30005 5944 30715 5946
rect 30005 5888 30010 5944
rect 30066 5888 30654 5944
rect 30710 5888 30715 5944
rect 30005 5886 30715 5888
rect 30005 5883 30071 5886
rect 30649 5883 30715 5886
rect 32397 5946 32463 5949
rect 33593 5946 33659 5949
rect 32397 5944 33659 5946
rect 32397 5888 32402 5944
rect 32458 5888 33598 5944
rect 33654 5888 33659 5944
rect 32397 5886 33659 5888
rect 32397 5883 32463 5886
rect 33593 5883 33659 5886
rect 34513 5946 34579 5949
rect 34646 5946 34652 5948
rect 34513 5944 34652 5946
rect 34513 5888 34518 5944
rect 34574 5888 34652 5944
rect 34513 5886 34652 5888
rect 34513 5883 34579 5886
rect 34646 5884 34652 5886
rect 34716 5884 34722 5948
rect 17585 5812 17651 5813
rect 17534 5748 17540 5812
rect 17604 5810 17651 5812
rect 30281 5810 30347 5813
rect 17604 5808 30347 5810
rect 17646 5752 30286 5808
rect 30342 5752 30347 5808
rect 17604 5750 30347 5752
rect 17604 5748 17651 5750
rect 17585 5747 17651 5748
rect 30281 5747 30347 5750
rect 31017 5810 31083 5813
rect 33593 5810 33659 5813
rect 31017 5808 33659 5810
rect 31017 5752 31022 5808
rect 31078 5752 33598 5808
rect 33654 5752 33659 5808
rect 31017 5750 33659 5752
rect 31017 5747 31083 5750
rect 33593 5747 33659 5750
rect 33961 5810 34027 5813
rect 35750 5810 35756 5812
rect 33961 5808 35756 5810
rect 33961 5752 33966 5808
rect 34022 5752 35756 5808
rect 33961 5750 35756 5752
rect 33961 5747 34027 5750
rect 35750 5748 35756 5750
rect 35820 5748 35826 5812
rect 15469 5674 15535 5677
rect 32397 5674 32463 5677
rect 15469 5672 32463 5674
rect 15469 5616 15474 5672
rect 15530 5616 32402 5672
rect 32458 5616 32463 5672
rect 15469 5614 32463 5616
rect 15469 5611 15535 5614
rect 32397 5611 32463 5614
rect 33225 5674 33291 5677
rect 36169 5674 36235 5677
rect 33225 5672 36235 5674
rect 33225 5616 33230 5672
rect 33286 5616 36174 5672
rect 36230 5616 36235 5672
rect 33225 5614 36235 5616
rect 33225 5611 33291 5614
rect 36169 5611 36235 5614
rect 20161 5538 20227 5541
rect 23657 5538 23723 5541
rect 20161 5536 23723 5538
rect 20161 5480 20166 5536
rect 20222 5480 23662 5536
rect 23718 5480 23723 5536
rect 20161 5478 23723 5480
rect 20161 5475 20227 5478
rect 23657 5475 23723 5478
rect 24301 5538 24367 5541
rect 25589 5538 25655 5541
rect 24301 5536 25655 5538
rect 24301 5480 24306 5536
rect 24362 5480 25594 5536
rect 25650 5480 25655 5536
rect 24301 5478 25655 5480
rect 24301 5475 24367 5478
rect 25589 5475 25655 5478
rect 27797 5538 27863 5541
rect 30649 5538 30715 5541
rect 27797 5536 30715 5538
rect 27797 5480 27802 5536
rect 27858 5480 30654 5536
rect 30710 5480 30715 5536
rect 27797 5478 30715 5480
rect 27797 5475 27863 5478
rect 30649 5475 30715 5478
rect 31661 5538 31727 5541
rect 31845 5538 31911 5541
rect 31661 5536 31911 5538
rect 31661 5480 31666 5536
rect 31722 5480 31850 5536
rect 31906 5480 31911 5536
rect 31661 5478 31911 5480
rect 31661 5475 31727 5478
rect 31845 5475 31911 5478
rect 42333 5540 42399 5541
rect 42333 5536 42380 5540
rect 42444 5538 42450 5540
rect 58157 5538 58223 5541
rect 59200 5538 60000 5568
rect 42333 5480 42338 5536
rect 42333 5476 42380 5480
rect 42444 5478 42490 5538
rect 58157 5536 60000 5538
rect 58157 5480 58162 5536
rect 58218 5480 60000 5536
rect 58157 5478 60000 5480
rect 42444 5476 42450 5478
rect 42333 5475 42399 5476
rect 58157 5475 58223 5478
rect 19570 5472 19886 5473
rect 0 5402 800 5432
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 59200 5448 60000 5478
rect 50290 5407 50606 5408
rect 1853 5402 1919 5405
rect 0 5400 1919 5402
rect 0 5344 1858 5400
rect 1914 5344 1919 5400
rect 0 5342 1919 5344
rect 0 5312 800 5342
rect 1853 5339 1919 5342
rect 20253 5404 20319 5405
rect 20253 5400 20300 5404
rect 20364 5402 20370 5404
rect 28901 5402 28967 5405
rect 31845 5402 31911 5405
rect 20253 5344 20258 5400
rect 20253 5340 20300 5344
rect 20364 5342 20410 5402
rect 28901 5400 31911 5402
rect 28901 5344 28906 5400
rect 28962 5344 31850 5400
rect 31906 5344 31911 5400
rect 28901 5342 31911 5344
rect 20364 5340 20370 5342
rect 20253 5339 20319 5340
rect 28901 5339 28967 5342
rect 31845 5339 31911 5342
rect 35433 5402 35499 5405
rect 43989 5402 44055 5405
rect 35433 5400 44055 5402
rect 35433 5344 35438 5400
rect 35494 5344 43994 5400
rect 44050 5344 44055 5400
rect 35433 5342 44055 5344
rect 35433 5339 35499 5342
rect 43989 5339 44055 5342
rect 12157 5266 12223 5269
rect 14089 5266 14155 5269
rect 12157 5264 14155 5266
rect 12157 5208 12162 5264
rect 12218 5208 14094 5264
rect 14150 5208 14155 5264
rect 12157 5206 14155 5208
rect 12157 5203 12223 5206
rect 14089 5203 14155 5206
rect 18137 5266 18203 5269
rect 22829 5266 22895 5269
rect 32397 5266 32463 5269
rect 36813 5266 36879 5269
rect 18137 5264 36879 5266
rect 18137 5208 18142 5264
rect 18198 5208 22834 5264
rect 22890 5208 32402 5264
rect 32458 5208 36818 5264
rect 36874 5208 36879 5264
rect 18137 5206 36879 5208
rect 18137 5203 18203 5206
rect 22829 5203 22895 5206
rect 32397 5203 32463 5206
rect 36813 5203 36879 5206
rect 3141 5130 3207 5133
rect 18781 5130 18847 5133
rect 3141 5128 18847 5130
rect 3141 5072 3146 5128
rect 3202 5072 18786 5128
rect 18842 5072 18847 5128
rect 3141 5070 18847 5072
rect 3141 5067 3207 5070
rect 18781 5067 18847 5070
rect 19333 5130 19399 5133
rect 20345 5130 20411 5133
rect 19333 5128 20411 5130
rect 19333 5072 19338 5128
rect 19394 5072 20350 5128
rect 20406 5072 20411 5128
rect 19333 5070 20411 5072
rect 19333 5067 19399 5070
rect 20345 5067 20411 5070
rect 23473 5130 23539 5133
rect 24710 5130 24716 5132
rect 23473 5128 24716 5130
rect 23473 5072 23478 5128
rect 23534 5072 24716 5128
rect 23473 5070 24716 5072
rect 23473 5067 23539 5070
rect 24710 5068 24716 5070
rect 24780 5068 24786 5132
rect 31385 5130 31451 5133
rect 35893 5130 35959 5133
rect 31385 5128 35959 5130
rect 31385 5072 31390 5128
rect 31446 5072 35898 5128
rect 35954 5072 35959 5128
rect 31385 5070 35959 5072
rect 31385 5067 31451 5070
rect 35893 5067 35959 5070
rect 9305 4994 9371 4997
rect 18413 4994 18479 4997
rect 32765 4994 32831 4997
rect 9305 4992 17970 4994
rect 9305 4936 9310 4992
rect 9366 4936 17970 4992
rect 9305 4934 17970 4936
rect 9305 4931 9371 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 8661 4858 8727 4861
rect 9581 4858 9647 4861
rect 8661 4856 9647 4858
rect 8661 4800 8666 4856
rect 8722 4800 9586 4856
rect 9642 4800 9647 4856
rect 8661 4798 9647 4800
rect 17910 4858 17970 4934
rect 18413 4992 32831 4994
rect 18413 4936 18418 4992
rect 18474 4936 32770 4992
rect 32826 4936 32831 4992
rect 18413 4934 32831 4936
rect 18413 4931 18479 4934
rect 32765 4931 32831 4934
rect 58065 4994 58131 4997
rect 59200 4994 60000 5024
rect 58065 4992 60000 4994
rect 58065 4936 58070 4992
rect 58126 4936 60000 4992
rect 58065 4934 60000 4936
rect 58065 4931 58131 4934
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 59200 4904 60000 4934
rect 34930 4863 35246 4864
rect 28809 4858 28875 4861
rect 17910 4856 28875 4858
rect 17910 4800 28814 4856
rect 28870 4800 28875 4856
rect 17910 4798 28875 4800
rect 8661 4795 8727 4798
rect 9581 4795 9647 4798
rect 28809 4795 28875 4798
rect 36261 4858 36327 4861
rect 37825 4858 37891 4861
rect 36261 4856 37891 4858
rect 36261 4800 36266 4856
rect 36322 4800 37830 4856
rect 37886 4800 37891 4856
rect 36261 4798 37891 4800
rect 36261 4795 36327 4798
rect 37825 4795 37891 4798
rect 0 4722 800 4752
rect 1761 4722 1827 4725
rect 28349 4722 28415 4725
rect 0 4720 1827 4722
rect 0 4664 1766 4720
rect 1822 4664 1827 4720
rect 0 4662 1827 4664
rect 0 4632 800 4662
rect 1761 4659 1827 4662
rect 9630 4720 28415 4722
rect 9630 4664 28354 4720
rect 28410 4664 28415 4720
rect 9630 4662 28415 4664
rect 9213 4314 9279 4317
rect 9630 4314 9690 4662
rect 28349 4659 28415 4662
rect 28625 4722 28691 4725
rect 32673 4722 32739 4725
rect 28625 4720 32739 4722
rect 28625 4664 28630 4720
rect 28686 4664 32678 4720
rect 32734 4664 32739 4720
rect 28625 4662 32739 4664
rect 28625 4659 28691 4662
rect 32673 4659 32739 4662
rect 34421 4724 34487 4725
rect 34421 4720 34468 4724
rect 34532 4722 34538 4724
rect 35525 4722 35591 4725
rect 38377 4722 38443 4725
rect 34421 4664 34426 4720
rect 34421 4660 34468 4664
rect 34532 4662 34578 4722
rect 35525 4720 38443 4722
rect 35525 4664 35530 4720
rect 35586 4664 38382 4720
rect 38438 4664 38443 4720
rect 35525 4662 38443 4664
rect 34532 4660 34538 4662
rect 34421 4659 34487 4660
rect 35525 4659 35591 4662
rect 38377 4659 38443 4662
rect 43253 4722 43319 4725
rect 45553 4722 45619 4725
rect 43253 4720 45619 4722
rect 43253 4664 43258 4720
rect 43314 4664 45558 4720
rect 45614 4664 45619 4720
rect 43253 4662 45619 4664
rect 43253 4659 43319 4662
rect 45553 4659 45619 4662
rect 10593 4586 10659 4589
rect 28165 4586 28231 4589
rect 10593 4584 28231 4586
rect 10593 4528 10598 4584
rect 10654 4528 28170 4584
rect 28226 4528 28231 4584
rect 10593 4526 28231 4528
rect 10593 4523 10659 4526
rect 28165 4523 28231 4526
rect 29361 4586 29427 4589
rect 32949 4586 33015 4589
rect 43713 4586 43779 4589
rect 52821 4586 52887 4589
rect 29361 4584 33015 4586
rect 29361 4528 29366 4584
rect 29422 4528 32954 4584
rect 33010 4528 33015 4584
rect 29361 4526 33015 4528
rect 29361 4523 29427 4526
rect 32949 4523 33015 4526
rect 41370 4584 52887 4586
rect 41370 4528 43718 4584
rect 43774 4528 52826 4584
rect 52882 4528 52887 4584
rect 41370 4526 52887 4528
rect 19977 4450 20043 4453
rect 22461 4450 22527 4453
rect 41370 4450 41430 4526
rect 43713 4523 43779 4526
rect 52821 4523 52887 4526
rect 19977 4448 21834 4450
rect 19977 4392 19982 4448
rect 20038 4392 21834 4448
rect 19977 4390 21834 4392
rect 19977 4387 20043 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 9213 4312 9690 4314
rect 9213 4256 9218 4312
rect 9274 4256 9690 4312
rect 9213 4254 9690 4256
rect 9213 4251 9279 4254
rect 20110 4252 20116 4316
rect 20180 4314 20186 4316
rect 20437 4314 20503 4317
rect 20180 4312 20503 4314
rect 20180 4256 20442 4312
rect 20498 4256 20503 4312
rect 20180 4254 20503 4256
rect 20180 4252 20186 4254
rect 20437 4251 20503 4254
rect 20713 4314 20779 4317
rect 21541 4314 21607 4317
rect 20713 4312 21607 4314
rect 20713 4256 20718 4312
rect 20774 4256 21546 4312
rect 21602 4256 21607 4312
rect 20713 4254 21607 4256
rect 21774 4314 21834 4390
rect 22461 4448 41430 4450
rect 22461 4392 22466 4448
rect 22522 4392 41430 4448
rect 22461 4390 41430 4392
rect 22461 4387 22527 4390
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 59200 4360 60000 4480
rect 50290 4319 50606 4320
rect 23105 4314 23171 4317
rect 21774 4312 23171 4314
rect 21774 4256 23110 4312
rect 23166 4256 23171 4312
rect 21774 4254 23171 4256
rect 20713 4251 20779 4254
rect 21541 4251 21607 4254
rect 23105 4251 23171 4254
rect 27981 4314 28047 4317
rect 36261 4314 36327 4317
rect 27981 4312 36327 4314
rect 27981 4256 27986 4312
rect 28042 4256 36266 4312
rect 36322 4256 36327 4312
rect 27981 4254 36327 4256
rect 27981 4251 28047 4254
rect 36261 4251 36327 4254
rect 9121 4178 9187 4181
rect 12985 4178 13051 4181
rect 9121 4176 13051 4178
rect 9121 4120 9126 4176
rect 9182 4120 12990 4176
rect 13046 4120 13051 4176
rect 9121 4118 13051 4120
rect 9121 4115 9187 4118
rect 12985 4115 13051 4118
rect 16941 4178 17007 4181
rect 26417 4178 26483 4181
rect 16941 4176 26483 4178
rect 16941 4120 16946 4176
rect 17002 4120 26422 4176
rect 26478 4120 26483 4176
rect 16941 4118 26483 4120
rect 16941 4115 17007 4118
rect 26417 4115 26483 4118
rect 29453 4178 29519 4181
rect 30465 4178 30531 4181
rect 31753 4178 31819 4181
rect 29453 4176 31819 4178
rect 29453 4120 29458 4176
rect 29514 4120 30470 4176
rect 30526 4120 31758 4176
rect 31814 4120 31819 4176
rect 29453 4118 31819 4120
rect 29453 4115 29519 4118
rect 30465 4115 30531 4118
rect 31753 4115 31819 4118
rect 33501 4178 33567 4181
rect 35893 4178 35959 4181
rect 33501 4176 35959 4178
rect 33501 4120 33506 4176
rect 33562 4120 35898 4176
rect 35954 4120 35959 4176
rect 33501 4118 35959 4120
rect 33501 4115 33567 4118
rect 35893 4115 35959 4118
rect 42977 4178 43043 4181
rect 44541 4178 44607 4181
rect 42977 4176 44607 4178
rect 42977 4120 42982 4176
rect 43038 4120 44546 4176
rect 44602 4120 44607 4176
rect 42977 4118 44607 4120
rect 42977 4115 43043 4118
rect 44541 4115 44607 4118
rect 0 4042 800 4072
rect 1761 4042 1827 4045
rect 0 4040 1827 4042
rect 0 3984 1766 4040
rect 1822 3984 1827 4040
rect 0 3982 1827 3984
rect 0 3952 800 3982
rect 1761 3979 1827 3982
rect 17125 4044 17191 4045
rect 17125 4040 17172 4044
rect 17236 4042 17242 4044
rect 18505 4042 18571 4045
rect 18638 4042 18644 4044
rect 17125 3984 17130 4040
rect 17125 3980 17172 3984
rect 17236 3982 17282 4042
rect 18505 4040 18644 4042
rect 18505 3984 18510 4040
rect 18566 3984 18644 4040
rect 18505 3982 18644 3984
rect 17236 3980 17242 3982
rect 17125 3979 17191 3980
rect 18505 3979 18571 3982
rect 18638 3980 18644 3982
rect 18708 3980 18714 4044
rect 19425 4042 19491 4045
rect 20478 4042 20484 4044
rect 19425 4040 20484 4042
rect 19425 3984 19430 4040
rect 19486 3984 20484 4040
rect 19425 3982 20484 3984
rect 19425 3979 19491 3982
rect 20478 3980 20484 3982
rect 20548 3980 20554 4044
rect 22318 3980 22324 4044
rect 22388 4042 22394 4044
rect 22737 4042 22803 4045
rect 22388 4040 22803 4042
rect 22388 3984 22742 4040
rect 22798 3984 22803 4040
rect 22388 3982 22803 3984
rect 22388 3980 22394 3982
rect 22737 3979 22803 3982
rect 29453 4042 29519 4045
rect 30005 4042 30071 4045
rect 29453 4040 30071 4042
rect 29453 3984 29458 4040
rect 29514 3984 30010 4040
rect 30066 3984 30071 4040
rect 29453 3982 30071 3984
rect 29453 3979 29519 3982
rect 30005 3979 30071 3982
rect 36721 4042 36787 4045
rect 36854 4042 36860 4044
rect 36721 4040 36860 4042
rect 36721 3984 36726 4040
rect 36782 3984 36860 4040
rect 36721 3982 36860 3984
rect 36721 3979 36787 3982
rect 36854 3980 36860 3982
rect 36924 3980 36930 4044
rect 39021 4042 39087 4045
rect 40585 4044 40651 4045
rect 40534 4042 40540 4044
rect 37782 4040 39087 4042
rect 37782 3984 39026 4040
rect 39082 3984 39087 4040
rect 37782 3982 39087 3984
rect 40494 3982 40540 4042
rect 40604 4040 40651 4044
rect 40646 3984 40651 4040
rect 12525 3906 12591 3909
rect 21909 3906 21975 3909
rect 12525 3904 21975 3906
rect 12525 3848 12530 3904
rect 12586 3848 21914 3904
rect 21970 3848 21975 3904
rect 12525 3846 21975 3848
rect 12525 3843 12591 3846
rect 21909 3843 21975 3846
rect 24393 3906 24459 3909
rect 28625 3906 28691 3909
rect 24393 3904 28691 3906
rect 24393 3848 24398 3904
rect 24454 3848 28630 3904
rect 28686 3848 28691 3904
rect 24393 3846 28691 3848
rect 24393 3843 24459 3846
rect 28625 3843 28691 3846
rect 35709 3906 35775 3909
rect 37782 3906 37842 3982
rect 39021 3979 39087 3982
rect 40534 3980 40540 3982
rect 40604 3980 40651 3984
rect 41822 3980 41828 4044
rect 41892 4042 41898 4044
rect 41965 4042 42031 4045
rect 41892 4040 42031 4042
rect 41892 3984 41970 4040
rect 42026 3984 42031 4040
rect 41892 3982 42031 3984
rect 41892 3980 41898 3982
rect 40585 3979 40651 3980
rect 41965 3979 42031 3982
rect 43345 4042 43411 4045
rect 43478 4042 43484 4044
rect 43345 4040 43484 4042
rect 43345 3984 43350 4040
rect 43406 3984 43484 4040
rect 43345 3982 43484 3984
rect 43345 3979 43411 3982
rect 43478 3980 43484 3982
rect 43548 3980 43554 4044
rect 53373 4042 53439 4045
rect 51030 4040 53439 4042
rect 51030 3984 53378 4040
rect 53434 3984 53439 4040
rect 51030 3982 53439 3984
rect 35709 3904 37842 3906
rect 35709 3848 35714 3904
rect 35770 3848 37842 3904
rect 35709 3846 37842 3848
rect 38009 3906 38075 3909
rect 49325 3906 49391 3909
rect 38009 3904 49391 3906
rect 38009 3848 38014 3904
rect 38070 3848 49330 3904
rect 49386 3848 49391 3904
rect 38009 3846 49391 3848
rect 35709 3843 35775 3846
rect 38009 3843 38075 3846
rect 49325 3843 49391 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 18505 3770 18571 3773
rect 19374 3770 19380 3772
rect 18505 3768 19380 3770
rect 18505 3712 18510 3768
rect 18566 3712 19380 3768
rect 18505 3710 19380 3712
rect 18505 3707 18571 3710
rect 19374 3708 19380 3710
rect 19444 3770 19450 3772
rect 19609 3770 19675 3773
rect 20621 3772 20687 3773
rect 20621 3770 20668 3772
rect 19444 3768 19675 3770
rect 19444 3712 19614 3768
rect 19670 3712 19675 3768
rect 19444 3710 19675 3712
rect 20576 3768 20668 3770
rect 20576 3712 20626 3768
rect 20576 3710 20668 3712
rect 19444 3708 19450 3710
rect 19609 3707 19675 3710
rect 20621 3708 20668 3710
rect 20732 3708 20738 3772
rect 21817 3770 21883 3773
rect 25497 3770 25563 3773
rect 21817 3768 25563 3770
rect 21817 3712 21822 3768
rect 21878 3712 25502 3768
rect 25558 3712 25563 3768
rect 21817 3710 25563 3712
rect 20621 3707 20687 3708
rect 21817 3707 21883 3710
rect 25497 3707 25563 3710
rect 35893 3770 35959 3773
rect 51030 3770 51090 3982
rect 53373 3979 53439 3982
rect 57881 3906 57947 3909
rect 59200 3906 60000 3936
rect 57881 3904 60000 3906
rect 57881 3848 57886 3904
rect 57942 3848 60000 3904
rect 57881 3846 60000 3848
rect 57881 3843 57947 3846
rect 59200 3816 60000 3846
rect 35893 3768 51090 3770
rect 35893 3712 35898 3768
rect 35954 3712 51090 3768
rect 35893 3710 51090 3712
rect 35893 3707 35959 3710
rect 15285 3634 15351 3637
rect 21265 3634 21331 3637
rect 15285 3632 21331 3634
rect 15285 3576 15290 3632
rect 15346 3576 21270 3632
rect 21326 3576 21331 3632
rect 15285 3574 21331 3576
rect 15285 3571 15351 3574
rect 21265 3571 21331 3574
rect 24393 3634 24459 3637
rect 24945 3634 25011 3637
rect 24393 3632 25011 3634
rect 24393 3576 24398 3632
rect 24454 3576 24950 3632
rect 25006 3576 25011 3632
rect 24393 3574 25011 3576
rect 24393 3571 24459 3574
rect 24945 3571 25011 3574
rect 25129 3634 25195 3637
rect 25773 3634 25839 3637
rect 25129 3632 25839 3634
rect 25129 3576 25134 3632
rect 25190 3576 25778 3632
rect 25834 3576 25839 3632
rect 25129 3574 25839 3576
rect 25129 3571 25195 3574
rect 25773 3571 25839 3574
rect 28993 3634 29059 3637
rect 33225 3634 33291 3637
rect 28993 3632 33291 3634
rect 28993 3576 28998 3632
rect 29054 3576 33230 3632
rect 33286 3576 33291 3632
rect 28993 3574 33291 3576
rect 28993 3571 29059 3574
rect 33225 3571 33291 3574
rect 36905 3634 36971 3637
rect 43529 3634 43595 3637
rect 49693 3634 49759 3637
rect 36905 3632 41430 3634
rect 36905 3576 36910 3632
rect 36966 3576 41430 3632
rect 36905 3574 41430 3576
rect 36905 3571 36971 3574
rect 12433 3498 12499 3501
rect 22185 3498 22251 3501
rect 12433 3496 22251 3498
rect 12433 3440 12438 3496
rect 12494 3440 22190 3496
rect 22246 3440 22251 3496
rect 12433 3438 22251 3440
rect 12433 3435 12499 3438
rect 22185 3435 22251 3438
rect 23105 3498 23171 3501
rect 39297 3498 39363 3501
rect 23105 3496 39363 3498
rect 23105 3440 23110 3496
rect 23166 3440 39302 3496
rect 39358 3440 39363 3496
rect 23105 3438 39363 3440
rect 23105 3435 23171 3438
rect 39297 3435 39363 3438
rect 0 3362 800 3392
rect 1853 3362 1919 3365
rect 0 3360 1919 3362
rect 0 3304 1858 3360
rect 1914 3304 1919 3360
rect 0 3302 1919 3304
rect 0 3272 800 3302
rect 1853 3299 1919 3302
rect 7465 3362 7531 3365
rect 9489 3362 9555 3365
rect 7465 3360 9555 3362
rect 7465 3304 7470 3360
rect 7526 3304 9494 3360
rect 9550 3304 9555 3360
rect 7465 3302 9555 3304
rect 7465 3299 7531 3302
rect 9489 3299 9555 3302
rect 20897 3362 20963 3365
rect 35433 3362 35499 3365
rect 20897 3360 35499 3362
rect 20897 3304 20902 3360
rect 20958 3304 35438 3360
rect 35494 3304 35499 3360
rect 20897 3302 35499 3304
rect 20897 3299 20963 3302
rect 35433 3299 35499 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 5165 3226 5231 3229
rect 11513 3226 11579 3229
rect 5165 3224 11579 3226
rect 5165 3168 5170 3224
rect 5226 3168 11518 3224
rect 11574 3168 11579 3224
rect 5165 3166 11579 3168
rect 5165 3163 5231 3166
rect 11513 3163 11579 3166
rect 12065 3226 12131 3229
rect 18597 3226 18663 3229
rect 19425 3228 19491 3229
rect 19374 3226 19380 3228
rect 12065 3224 18663 3226
rect 12065 3168 12070 3224
rect 12126 3168 18602 3224
rect 18658 3168 18663 3224
rect 12065 3166 18663 3168
rect 19334 3166 19380 3226
rect 19444 3224 19491 3228
rect 19486 3168 19491 3224
rect 12065 3163 12131 3166
rect 18597 3163 18663 3166
rect 19374 3164 19380 3166
rect 19444 3164 19491 3168
rect 19425 3163 19491 3164
rect 20069 3226 20135 3229
rect 23933 3226 23999 3229
rect 20069 3224 23999 3226
rect 20069 3168 20074 3224
rect 20130 3168 23938 3224
rect 23994 3168 23999 3224
rect 20069 3166 23999 3168
rect 20069 3163 20135 3166
rect 23933 3163 23999 3166
rect 24117 3226 24183 3229
rect 32305 3226 32371 3229
rect 24117 3224 32371 3226
rect 24117 3168 24122 3224
rect 24178 3168 32310 3224
rect 32366 3168 32371 3224
rect 24117 3166 32371 3168
rect 24117 3163 24183 3166
rect 32305 3163 32371 3166
rect 34145 3226 34211 3229
rect 37457 3226 37523 3229
rect 34145 3224 37523 3226
rect 34145 3168 34150 3224
rect 34206 3168 37462 3224
rect 37518 3168 37523 3224
rect 34145 3166 37523 3168
rect 41370 3226 41430 3574
rect 43529 3632 49759 3634
rect 43529 3576 43534 3632
rect 43590 3576 49698 3632
rect 49754 3576 49759 3632
rect 43529 3574 49759 3576
rect 43529 3571 43595 3574
rect 49693 3571 49759 3574
rect 42149 3498 42215 3501
rect 46565 3498 46631 3501
rect 42149 3496 46631 3498
rect 42149 3440 42154 3496
rect 42210 3440 46570 3496
rect 46626 3440 46631 3496
rect 42149 3438 46631 3440
rect 42149 3435 42215 3438
rect 46565 3435 46631 3438
rect 42609 3362 42675 3365
rect 48037 3362 48103 3365
rect 42609 3360 48103 3362
rect 42609 3304 42614 3360
rect 42670 3304 48042 3360
rect 48098 3304 48103 3360
rect 42609 3302 48103 3304
rect 42609 3299 42675 3302
rect 48037 3299 48103 3302
rect 58157 3362 58223 3365
rect 59200 3362 60000 3392
rect 58157 3360 60000 3362
rect 58157 3304 58162 3360
rect 58218 3304 60000 3360
rect 58157 3302 60000 3304
rect 58157 3299 58223 3302
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 59200 3272 60000 3302
rect 50290 3231 50606 3232
rect 49693 3226 49759 3229
rect 41370 3224 49759 3226
rect 41370 3168 49698 3224
rect 49754 3168 49759 3224
rect 41370 3166 49759 3168
rect 34145 3163 34211 3166
rect 37457 3163 37523 3166
rect 49693 3163 49759 3166
rect 16573 3090 16639 3093
rect 22093 3090 22159 3093
rect 16573 3088 22159 3090
rect 16573 3032 16578 3088
rect 16634 3032 22098 3088
rect 22154 3032 22159 3088
rect 16573 3030 22159 3032
rect 16573 3027 16639 3030
rect 22093 3027 22159 3030
rect 22921 3090 22987 3093
rect 28533 3090 28599 3093
rect 22921 3088 28599 3090
rect 22921 3032 22926 3088
rect 22982 3032 28538 3088
rect 28594 3032 28599 3088
rect 22921 3030 28599 3032
rect 22921 3027 22987 3030
rect 28533 3027 28599 3030
rect 41965 3090 42031 3093
rect 44357 3090 44423 3093
rect 41965 3088 44423 3090
rect 41965 3032 41970 3088
rect 42026 3032 44362 3088
rect 44418 3032 44423 3088
rect 41965 3030 44423 3032
rect 41965 3027 42031 3030
rect 44357 3027 44423 3030
rect 6729 2954 6795 2957
rect 9857 2954 9923 2957
rect 6729 2952 9923 2954
rect 6729 2896 6734 2952
rect 6790 2896 9862 2952
rect 9918 2896 9923 2952
rect 6729 2894 9923 2896
rect 6729 2891 6795 2894
rect 9857 2891 9923 2894
rect 15837 2954 15903 2957
rect 19793 2954 19859 2957
rect 15837 2952 19859 2954
rect 15837 2896 15842 2952
rect 15898 2896 19798 2952
rect 19854 2896 19859 2952
rect 15837 2894 19859 2896
rect 15837 2891 15903 2894
rect 19793 2891 19859 2894
rect 19977 2954 20043 2957
rect 30097 2954 30163 2957
rect 19977 2952 30163 2954
rect 19977 2896 19982 2952
rect 20038 2896 30102 2952
rect 30158 2896 30163 2952
rect 19977 2894 30163 2896
rect 19977 2891 20043 2894
rect 30097 2891 30163 2894
rect 44357 2954 44423 2957
rect 44817 2954 44883 2957
rect 44357 2952 44883 2954
rect 44357 2896 44362 2952
rect 44418 2896 44822 2952
rect 44878 2896 44883 2952
rect 44357 2894 44883 2896
rect 44357 2891 44423 2894
rect 44817 2891 44883 2894
rect 14273 2818 14339 2821
rect 20069 2818 20135 2821
rect 14273 2816 20135 2818
rect 14273 2760 14278 2816
rect 14334 2760 20074 2816
rect 20130 2760 20135 2816
rect 14273 2758 20135 2760
rect 14273 2755 14339 2758
rect 20069 2755 20135 2758
rect 20294 2756 20300 2820
rect 20364 2818 20370 2820
rect 20713 2818 20779 2821
rect 20364 2816 20779 2818
rect 20364 2760 20718 2816
rect 20774 2760 20779 2816
rect 20364 2758 20779 2760
rect 20364 2756 20370 2758
rect 20713 2755 20779 2758
rect 20897 2818 20963 2821
rect 23105 2818 23171 2821
rect 20897 2816 23171 2818
rect 20897 2760 20902 2816
rect 20958 2760 23110 2816
rect 23166 2760 23171 2816
rect 20897 2758 23171 2760
rect 20897 2755 20963 2758
rect 23105 2755 23171 2758
rect 57881 2818 57947 2821
rect 59200 2818 60000 2848
rect 57881 2816 60000 2818
rect 57881 2760 57886 2816
rect 57942 2760 60000 2816
rect 57881 2758 60000 2760
rect 57881 2755 57947 2758
rect 4210 2752 4526 2753
rect 0 2682 800 2712
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 1761 2682 1827 2685
rect 0 2680 1827 2682
rect 0 2624 1766 2680
rect 1822 2624 1827 2680
rect 0 2622 1827 2624
rect 0 2592 800 2622
rect 1761 2619 1827 2622
rect 12065 2682 12131 2685
rect 12617 2682 12683 2685
rect 12065 2680 12683 2682
rect 12065 2624 12070 2680
rect 12126 2624 12622 2680
rect 12678 2624 12683 2680
rect 12065 2622 12683 2624
rect 12065 2619 12131 2622
rect 12617 2619 12683 2622
rect 13261 2684 13327 2685
rect 13261 2680 13308 2684
rect 13372 2682 13378 2684
rect 18689 2682 18755 2685
rect 20621 2682 20687 2685
rect 13261 2624 13266 2680
rect 13261 2620 13308 2624
rect 13372 2622 13418 2682
rect 18689 2680 20687 2682
rect 18689 2624 18694 2680
rect 18750 2624 20626 2680
rect 20682 2624 20687 2680
rect 18689 2622 20687 2624
rect 13372 2620 13378 2622
rect 13261 2619 13327 2620
rect 18689 2619 18755 2622
rect 20621 2619 20687 2622
rect 20897 2682 20963 2685
rect 21030 2682 21036 2684
rect 20897 2680 21036 2682
rect 20897 2624 20902 2680
rect 20958 2624 21036 2680
rect 20897 2622 21036 2624
rect 20897 2619 20963 2622
rect 21030 2620 21036 2622
rect 21100 2620 21106 2684
rect 21766 2620 21772 2684
rect 21836 2682 21842 2684
rect 22001 2682 22067 2685
rect 21836 2680 22067 2682
rect 21836 2624 22006 2680
rect 22062 2624 22067 2680
rect 21836 2622 22067 2624
rect 21836 2620 21842 2622
rect 22001 2619 22067 2622
rect 22870 2620 22876 2684
rect 22940 2682 22946 2684
rect 23013 2682 23079 2685
rect 22940 2680 23079 2682
rect 22940 2624 23018 2680
rect 23074 2624 23079 2680
rect 22940 2622 23079 2624
rect 22940 2620 22946 2622
rect 23013 2619 23079 2622
rect 39430 2620 39436 2684
rect 39500 2682 39506 2684
rect 40217 2682 40283 2685
rect 41321 2684 41387 2685
rect 41270 2682 41276 2684
rect 39500 2680 40283 2682
rect 39500 2624 40222 2680
rect 40278 2624 40283 2680
rect 39500 2622 40283 2624
rect 41230 2622 41276 2682
rect 41340 2680 41387 2684
rect 41382 2624 41387 2680
rect 39500 2620 39506 2622
rect 40217 2619 40283 2622
rect 41270 2620 41276 2622
rect 41340 2620 41387 2624
rect 41321 2619 41387 2620
rect 42793 2682 42859 2685
rect 42926 2682 42932 2684
rect 42793 2680 42932 2682
rect 42793 2624 42798 2680
rect 42854 2624 42932 2680
rect 42793 2622 42932 2624
rect 42793 2619 42859 2622
rect 42926 2620 42932 2622
rect 42996 2620 43002 2684
rect 8753 2546 8819 2549
rect 19977 2546 20043 2549
rect 30557 2546 30623 2549
rect 8753 2544 30623 2546
rect 8753 2488 8758 2544
rect 8814 2488 19982 2544
rect 20038 2488 30562 2544
rect 30618 2488 30623 2544
rect 8753 2486 30623 2488
rect 8753 2483 8819 2486
rect 19977 2483 20043 2486
rect 30557 2483 30623 2486
rect 11789 2410 11855 2413
rect 17125 2410 17191 2413
rect 11789 2408 17191 2410
rect 11789 2352 11794 2408
rect 11850 2352 17130 2408
rect 17186 2352 17191 2408
rect 11789 2350 17191 2352
rect 11789 2347 11855 2350
rect 17125 2347 17191 2350
rect 17953 2410 18019 2413
rect 43529 2410 43595 2413
rect 17953 2408 22110 2410
rect 17953 2352 17958 2408
rect 18014 2352 22110 2408
rect 17953 2350 22110 2352
rect 17953 2347 18019 2350
rect 22050 2274 22110 2350
rect 26190 2408 43595 2410
rect 26190 2352 43534 2408
rect 43590 2352 43595 2408
rect 26190 2350 43595 2352
rect 26190 2274 26250 2350
rect 43529 2347 43595 2350
rect 22050 2214 26250 2274
rect 56225 2274 56291 2277
rect 59200 2274 60000 2304
rect 56225 2272 60000 2274
rect 56225 2216 56230 2272
rect 56286 2216 60000 2272
rect 56225 2214 60000 2216
rect 56225 2211 56291 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 59200 2184 60000 2214
rect 50290 2143 50606 2144
rect 0 2002 800 2032
rect 1853 2002 1919 2005
rect 0 2000 1919 2002
rect 0 1944 1858 2000
rect 1914 1944 1919 2000
rect 0 1942 1919 1944
rect 0 1912 800 1942
rect 1853 1939 1919 1942
rect 8937 2002 9003 2005
rect 30281 2002 30347 2005
rect 8937 2000 30347 2002
rect 8937 1944 8942 2000
rect 8998 1944 30286 2000
rect 30342 1944 30347 2000
rect 8937 1942 30347 1944
rect 8937 1939 9003 1942
rect 30281 1939 30347 1942
rect 20437 1866 20503 1869
rect 25129 1866 25195 1869
rect 20437 1864 25195 1866
rect 20437 1808 20442 1864
rect 20498 1808 25134 1864
rect 25190 1808 25195 1864
rect 20437 1806 25195 1808
rect 20437 1803 20503 1806
rect 25129 1803 25195 1806
rect 18045 1730 18111 1733
rect 27061 1730 27127 1733
rect 18045 1728 27127 1730
rect 18045 1672 18050 1728
rect 18106 1672 27066 1728
rect 27122 1672 27127 1728
rect 18045 1670 27127 1672
rect 18045 1667 18111 1670
rect 27061 1667 27127 1670
rect 57237 1730 57303 1733
rect 59200 1730 60000 1760
rect 57237 1728 60000 1730
rect 57237 1672 57242 1728
rect 57298 1672 60000 1728
rect 57237 1670 60000 1672
rect 57237 1667 57303 1670
rect 59200 1640 60000 1670
rect 17217 1594 17283 1597
rect 25405 1594 25471 1597
rect 17217 1592 25471 1594
rect 17217 1536 17222 1592
rect 17278 1536 25410 1592
rect 25466 1536 25471 1592
rect 17217 1534 25471 1536
rect 17217 1531 17283 1534
rect 25405 1531 25471 1534
rect 14549 1458 14615 1461
rect 25681 1458 25747 1461
rect 14549 1456 25747 1458
rect 14549 1400 14554 1456
rect 14610 1400 25686 1456
rect 25742 1400 25747 1456
rect 14549 1398 25747 1400
rect 14549 1395 14615 1398
rect 25681 1395 25747 1398
rect 17493 1322 17559 1325
rect 29085 1322 29151 1325
rect 17493 1320 29151 1322
rect 17493 1264 17498 1320
rect 17554 1264 29090 1320
rect 29146 1264 29151 1320
rect 17493 1262 29151 1264
rect 17493 1259 17559 1262
rect 29085 1259 29151 1262
rect 15653 1186 15719 1189
rect 36077 1186 36143 1189
rect 15653 1184 36143 1186
rect 15653 1128 15658 1184
rect 15714 1128 36082 1184
rect 36138 1128 36143 1184
rect 15653 1126 36143 1128
rect 15653 1123 15719 1126
rect 36077 1123 36143 1126
rect 56501 1186 56567 1189
rect 59200 1186 60000 1216
rect 56501 1184 60000 1186
rect 56501 1128 56506 1184
rect 56562 1128 60000 1184
rect 56501 1126 60000 1128
rect 56501 1123 56567 1126
rect 59200 1096 60000 1126
rect 15101 1050 15167 1053
rect 27797 1050 27863 1053
rect 15101 1048 27863 1050
rect 15101 992 15106 1048
rect 15162 992 27802 1048
rect 27858 992 27863 1048
rect 15101 990 27863 992
rect 15101 987 15167 990
rect 27797 987 27863 990
rect 3693 914 3759 917
rect 33317 914 33383 917
rect 3693 912 33383 914
rect 3693 856 3698 912
rect 3754 856 33322 912
rect 33378 856 33383 912
rect 3693 854 33383 856
rect 3693 851 3759 854
rect 33317 851 33383 854
rect 19374 716 19380 780
rect 19444 778 19450 780
rect 24669 778 24735 781
rect 19444 776 24735 778
rect 19444 720 24674 776
rect 24730 720 24735 776
rect 19444 718 24735 720
rect 19444 716 19450 718
rect 24669 715 24735 718
rect 54477 98 54543 101
rect 56501 98 56567 101
rect 54477 96 56567 98
rect 54477 40 54482 96
rect 54538 40 56506 96
rect 56562 40 56567 96
rect 54477 38 56567 40
rect 54477 35 54543 38
rect 56501 35 56567 38
<< via3 >>
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 39252 61100 39316 61164
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 12940 60752 13004 60756
rect 12940 60696 12954 60752
rect 12954 60696 13004 60752
rect 12940 60692 13004 60696
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 18460 59392 18524 59396
rect 18460 59336 18510 59392
rect 18510 59336 18524 59392
rect 18460 59332 18524 59336
rect 23060 59332 23124 59396
rect 42380 59332 42444 59396
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 21956 58788 22020 58852
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 40356 58032 40420 58036
rect 40356 57976 40406 58032
rect 40406 57976 40420 58032
rect 40356 57972 40420 57976
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 43484 57292 43548 57356
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 33916 56612 33980 56676
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 36124 53076 36188 53140
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 31156 52532 31220 52596
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 32812 51716 32876 51780
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 36860 50356 36924 50420
rect 38516 50220 38580 50284
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 41828 47636 41892 47700
rect 30236 47500 30300 47564
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 34652 42876 34716 42940
rect 42932 42604 42996 42668
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 29868 41516 29932 41580
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 23796 38524 23860 38588
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 23244 35940 23308 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 22692 34444 22756 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 17540 30636 17604 30700
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 16068 28460 16132 28524
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 16436 26964 16500 27028
rect 34100 26828 34164 26892
rect 36676 26828 36740 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 36308 26284 36372 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 22140 24788 22204 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 20116 24244 20180 24308
rect 39436 24108 39500 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 23980 23428 24044 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 40724 22748 40788 22812
rect 41276 22612 41340 22676
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20300 22068 20364 22132
rect 14412 21932 14476 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 40540 20708 40604 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 39804 19000 39868 19004
rect 39804 18944 39854 19000
rect 39854 18944 39868 19000
rect 39804 18940 39868 18944
rect 13308 18668 13372 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 17356 17988 17420 18052
rect 22692 18048 22756 18052
rect 22692 17992 22742 18048
rect 22742 17992 22756 18048
rect 22692 17988 22756 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 20668 17852 20732 17916
rect 21772 17716 21836 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 17908 17172 17972 17236
rect 18460 16900 18524 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 33732 16220 33796 16284
rect 37228 15948 37292 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 17172 15540 17236 15604
rect 20484 15404 20548 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 21036 14860 21100 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 18644 14588 18708 14652
rect 22876 14316 22940 14380
rect 24716 14180 24780 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 35572 13772 35636 13836
rect 43852 13772 43916 13836
rect 16988 13636 17052 13700
rect 27108 13636 27172 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19380 13500 19444 13564
rect 34284 13500 34348 13564
rect 37228 13500 37292 13564
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 18460 12820 18524 12884
rect 19196 12684 19260 12748
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 27108 12684 27172 12748
rect 33548 12608 33612 12612
rect 33548 12552 33598 12608
rect 33598 12552 33612 12608
rect 33548 12548 33612 12552
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 16068 11460 16132 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 34468 11324 34532 11388
rect 40356 11324 40420 11388
rect 39252 11052 39316 11116
rect 40172 11052 40236 11116
rect 17908 10916 17972 10980
rect 36308 10916 36372 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 22140 10704 22204 10708
rect 22140 10648 22190 10704
rect 22190 10648 22204 10704
rect 22140 10644 22204 10648
rect 34652 10432 34716 10436
rect 34652 10376 34702 10432
rect 34702 10376 34716 10432
rect 34652 10372 34716 10376
rect 40724 10432 40788 10436
rect 40724 10376 40738 10432
rect 40738 10376 40788 10432
rect 40724 10372 40788 10376
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 34468 10236 34532 10300
rect 39988 10236 40052 10300
rect 19380 10024 19444 10028
rect 19380 9968 19430 10024
rect 19430 9968 19444 10024
rect 19380 9964 19444 9968
rect 20116 9964 20180 10028
rect 22324 9964 22388 10028
rect 23980 9828 24044 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 39804 9692 39868 9756
rect 33548 9556 33612 9620
rect 34284 9616 34348 9620
rect 34284 9560 34298 9616
rect 34298 9560 34348 9616
rect 34284 9556 34348 9560
rect 34468 9556 34532 9620
rect 35388 9556 35452 9620
rect 36124 9556 36188 9620
rect 38516 9556 38580 9620
rect 16068 9420 16132 9484
rect 20300 9420 20364 9484
rect 20852 9420 20916 9484
rect 38700 9480 38764 9484
rect 38700 9424 38714 9480
rect 38714 9424 38764 9480
rect 38700 9420 38764 9424
rect 23060 9284 23124 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 17356 9208 17420 9212
rect 17356 9152 17406 9208
rect 17406 9152 17420 9208
rect 17356 9148 17420 9152
rect 34468 9284 34532 9348
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 16436 8876 16500 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 20116 8604 20180 8668
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 23796 8528 23860 8532
rect 23796 8472 23810 8528
rect 23810 8472 23860 8528
rect 23796 8468 23860 8472
rect 35388 8604 35452 8668
rect 35572 8468 35636 8532
rect 36676 8468 36740 8532
rect 22324 8332 22388 8396
rect 33548 8332 33612 8396
rect 33732 8332 33796 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12940 7924 13004 7988
rect 23244 8060 23308 8124
rect 30236 8196 30300 8260
rect 33916 8256 33980 8260
rect 33916 8200 33930 8256
rect 33930 8200 33980 8256
rect 33916 8196 33980 8200
rect 34652 8256 34716 8260
rect 34652 8200 34666 8256
rect 34666 8200 34716 8256
rect 34652 8196 34716 8200
rect 39988 8196 40052 8260
rect 40172 8196 40236 8260
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 38700 7984 38764 7988
rect 38700 7928 38750 7984
rect 38750 7928 38764 7984
rect 38700 7924 38764 7928
rect 14412 7652 14476 7716
rect 16988 7652 17052 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 19380 7576 19444 7580
rect 19380 7520 19430 7576
rect 19430 7520 19444 7576
rect 19380 7516 19444 7520
rect 21956 7576 22020 7580
rect 21956 7520 22006 7576
rect 22006 7520 22020 7576
rect 21956 7516 22020 7520
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 18460 6896 18524 6900
rect 18460 6840 18474 6896
rect 18474 6840 18524 6896
rect 18460 6836 18524 6840
rect 20852 6836 20916 6900
rect 22324 6836 22388 6900
rect 29868 6836 29932 6900
rect 31156 6896 31220 6900
rect 31156 6840 31170 6896
rect 31170 6840 31220 6896
rect 31156 6836 31220 6840
rect 32812 6836 32876 6900
rect 43852 6896 43916 6900
rect 43852 6840 43866 6896
rect 43866 6840 43916 6896
rect 43852 6836 43916 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 19196 6428 19260 6492
rect 19380 6488 19444 6492
rect 19380 6432 19394 6488
rect 19394 6432 19444 6488
rect 19380 6428 19444 6432
rect 19380 6292 19444 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 34652 5884 34716 5948
rect 17540 5808 17604 5812
rect 17540 5752 17590 5808
rect 17590 5752 17604 5808
rect 17540 5748 17604 5752
rect 35756 5748 35820 5812
rect 42380 5536 42444 5540
rect 42380 5480 42394 5536
rect 42394 5480 42444 5536
rect 42380 5476 42444 5480
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 20300 5400 20364 5404
rect 20300 5344 20314 5400
rect 20314 5344 20364 5400
rect 20300 5340 20364 5344
rect 24716 5068 24780 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 34468 4720 34532 4724
rect 34468 4664 34482 4720
rect 34482 4664 34532 4720
rect 34468 4660 34532 4664
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 20116 4252 20180 4316
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 17172 4040 17236 4044
rect 17172 3984 17186 4040
rect 17186 3984 17236 4040
rect 17172 3980 17236 3984
rect 18644 3980 18708 4044
rect 20484 3980 20548 4044
rect 22324 3980 22388 4044
rect 36860 3980 36924 4044
rect 40540 4040 40604 4044
rect 40540 3984 40590 4040
rect 40590 3984 40604 4040
rect 40540 3980 40604 3984
rect 41828 3980 41892 4044
rect 43484 3980 43548 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19380 3708 19444 3772
rect 20668 3768 20732 3772
rect 20668 3712 20682 3768
rect 20682 3712 20732 3768
rect 20668 3708 20732 3712
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 19380 3224 19444 3228
rect 19380 3168 19430 3224
rect 19430 3168 19444 3224
rect 19380 3164 19444 3168
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 20300 2756 20364 2820
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 13308 2680 13372 2684
rect 13308 2624 13322 2680
rect 13322 2624 13372 2680
rect 13308 2620 13372 2624
rect 21036 2620 21100 2684
rect 21772 2620 21836 2684
rect 22876 2620 22940 2684
rect 39436 2620 39500 2684
rect 41276 2680 41340 2684
rect 41276 2624 41326 2680
rect 41326 2624 41340 2680
rect 41276 2620 41340 2624
rect 42932 2620 42996 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 19380 716 19444 780
<< metal4 >>
rect 4208 61504 4528 61520
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 19568 60960 19888 61520
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 12939 60756 13005 60757
rect 12939 60692 12940 60756
rect 13004 60692 13005 60756
rect 12939 60691 13005 60692
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 12942 7989 13002 60691
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 18459 59396 18525 59397
rect 18459 59332 18460 59396
rect 18524 59332 18525 59396
rect 18459 59331 18525 59332
rect 17539 30700 17605 30701
rect 17539 30636 17540 30700
rect 17604 30636 17605 30700
rect 17539 30635 17605 30636
rect 16067 28524 16133 28525
rect 16067 28460 16068 28524
rect 16132 28460 16133 28524
rect 16067 28459 16133 28460
rect 14411 21996 14477 21997
rect 14411 21932 14412 21996
rect 14476 21932 14477 21996
rect 14411 21931 14477 21932
rect 13307 18732 13373 18733
rect 13307 18668 13308 18732
rect 13372 18668 13373 18732
rect 13307 18667 13373 18668
rect 12939 7988 13005 7989
rect 12939 7924 12940 7988
rect 13004 7924 13005 7988
rect 12939 7923 13005 7924
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 13310 2685 13370 18667
rect 14414 7717 14474 21931
rect 16070 11525 16130 28459
rect 16435 27028 16501 27029
rect 16435 26964 16436 27028
rect 16500 26964 16501 27028
rect 16435 26963 16501 26964
rect 16067 11524 16133 11525
rect 16067 11460 16068 11524
rect 16132 11460 16133 11524
rect 16067 11459 16133 11460
rect 16070 9485 16130 11459
rect 16067 9484 16133 9485
rect 16067 9420 16068 9484
rect 16132 9420 16133 9484
rect 16067 9419 16133 9420
rect 16438 8941 16498 26963
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 17171 15604 17237 15605
rect 17171 15540 17172 15604
rect 17236 15540 17237 15604
rect 17171 15539 17237 15540
rect 16987 13700 17053 13701
rect 16987 13636 16988 13700
rect 17052 13636 17053 13700
rect 16987 13635 17053 13636
rect 16435 8940 16501 8941
rect 16435 8876 16436 8940
rect 16500 8876 16501 8940
rect 16435 8875 16501 8876
rect 16990 7717 17050 13635
rect 14411 7716 14477 7717
rect 14411 7652 14412 7716
rect 14476 7652 14477 7716
rect 14411 7651 14477 7652
rect 16987 7716 17053 7717
rect 16987 7652 16988 7716
rect 17052 7652 17053 7716
rect 16987 7651 17053 7652
rect 17174 4045 17234 15539
rect 17358 9213 17418 17987
rect 17355 9212 17421 9213
rect 17355 9148 17356 9212
rect 17420 9148 17421 9212
rect 17355 9147 17421 9148
rect 17542 5813 17602 30635
rect 17907 17236 17973 17237
rect 17907 17172 17908 17236
rect 17972 17172 17973 17236
rect 17907 17171 17973 17172
rect 17910 10981 17970 17171
rect 18462 16965 18522 59331
rect 19568 58784 19888 59808
rect 34928 61504 35248 61520
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 39251 61164 39317 61165
rect 39251 61100 39252 61164
rect 39316 61100 39317 61164
rect 39251 61099 39317 61100
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 23059 59396 23125 59397
rect 23059 59332 23060 59396
rect 23124 59332 23125 59396
rect 23059 59331 23125 59332
rect 21955 58852 22021 58853
rect 21955 58788 21956 58852
rect 22020 58788 22021 58852
rect 21955 58787 22021 58788
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 20115 24308 20181 24309
rect 20115 24244 20116 24308
rect 20180 24244 20181 24308
rect 20115 24243 20181 24244
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 18459 16964 18525 16965
rect 18459 16900 18460 16964
rect 18524 16900 18525 16964
rect 18459 16899 18525 16900
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 18643 14652 18709 14653
rect 18643 14588 18644 14652
rect 18708 14588 18709 14652
rect 18643 14587 18709 14588
rect 18459 12884 18525 12885
rect 18459 12820 18460 12884
rect 18524 12820 18525 12884
rect 18459 12819 18525 12820
rect 17907 10980 17973 10981
rect 17907 10916 17908 10980
rect 17972 10916 17973 10980
rect 17907 10915 17973 10916
rect 18462 6901 18522 12819
rect 18459 6900 18525 6901
rect 18459 6836 18460 6900
rect 18524 6836 18525 6900
rect 18459 6835 18525 6836
rect 17539 5812 17605 5813
rect 17539 5748 17540 5812
rect 17604 5748 17605 5812
rect 17539 5747 17605 5748
rect 18646 4045 18706 14587
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19195 12748 19261 12749
rect 19195 12684 19196 12748
rect 19260 12684 19261 12748
rect 19195 12683 19261 12684
rect 19198 6493 19258 12683
rect 19382 10029 19442 13499
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 10028 19445 10029
rect 19379 9964 19380 10028
rect 19444 9964 19445 10028
rect 19379 9963 19445 9964
rect 19568 9824 19888 10848
rect 20118 10029 20178 24243
rect 20299 22132 20365 22133
rect 20299 22068 20300 22132
rect 20364 22068 20365 22132
rect 20299 22067 20365 22068
rect 20115 10028 20181 10029
rect 20115 9964 20116 10028
rect 20180 9964 20181 10028
rect 20115 9963 20181 9964
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 20302 9485 20362 22067
rect 20667 17916 20733 17917
rect 20667 17852 20668 17916
rect 20732 17852 20733 17916
rect 20667 17851 20733 17852
rect 20483 15468 20549 15469
rect 20483 15404 20484 15468
rect 20548 15404 20549 15468
rect 20483 15403 20549 15404
rect 20299 9484 20365 9485
rect 20299 9420 20300 9484
rect 20364 9420 20365 9484
rect 20299 9419 20365 9420
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 20115 8668 20181 8669
rect 20115 8604 20116 8668
rect 20180 8604 20181 8668
rect 20115 8603 20181 8604
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19379 7580 19445 7581
rect 19379 7516 19380 7580
rect 19444 7516 19445 7580
rect 19379 7515 19445 7516
rect 19382 6493 19442 7515
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19195 6492 19261 6493
rect 19195 6428 19196 6492
rect 19260 6428 19261 6492
rect 19195 6427 19261 6428
rect 19379 6492 19445 6493
rect 19379 6428 19380 6492
rect 19444 6428 19445 6492
rect 19379 6427 19445 6428
rect 19379 6356 19445 6357
rect 19379 6292 19380 6356
rect 19444 6292 19445 6356
rect 19379 6291 19445 6292
rect 17171 4044 17237 4045
rect 17171 3980 17172 4044
rect 17236 3980 17237 4044
rect 17171 3979 17237 3980
rect 18643 4044 18709 4045
rect 18643 3980 18644 4044
rect 18708 3980 18709 4044
rect 18643 3979 18709 3980
rect 19382 3773 19442 6291
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 3772 19445 3773
rect 19379 3708 19380 3772
rect 19444 3708 19445 3772
rect 19379 3707 19445 3708
rect 19568 3296 19888 4320
rect 20118 4317 20178 8603
rect 20299 5404 20365 5405
rect 20299 5340 20300 5404
rect 20364 5340 20365 5404
rect 20299 5339 20365 5340
rect 20115 4316 20181 4317
rect 20115 4252 20116 4316
rect 20180 4252 20181 4316
rect 20115 4251 20181 4252
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 3228 19445 3229
rect 19379 3164 19380 3228
rect 19444 3164 19445 3228
rect 19379 3163 19445 3164
rect 13307 2684 13373 2685
rect 13307 2620 13308 2684
rect 13372 2620 13373 2684
rect 13307 2619 13373 2620
rect 19382 781 19442 3163
rect 19568 2208 19888 3232
rect 20302 2821 20362 5339
rect 20486 4045 20546 15403
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 20670 3773 20730 17851
rect 21771 17780 21837 17781
rect 21771 17716 21772 17780
rect 21836 17716 21837 17780
rect 21771 17715 21837 17716
rect 21035 14924 21101 14925
rect 21035 14860 21036 14924
rect 21100 14860 21101 14924
rect 21035 14859 21101 14860
rect 20851 9484 20917 9485
rect 20851 9420 20852 9484
rect 20916 9420 20917 9484
rect 20851 9419 20917 9420
rect 20854 6901 20914 9419
rect 20851 6900 20917 6901
rect 20851 6836 20852 6900
rect 20916 6836 20917 6900
rect 20851 6835 20917 6836
rect 20667 3772 20733 3773
rect 20667 3708 20668 3772
rect 20732 3708 20733 3772
rect 20667 3707 20733 3708
rect 20299 2820 20365 2821
rect 20299 2756 20300 2820
rect 20364 2756 20365 2820
rect 20299 2755 20365 2756
rect 21038 2685 21098 14859
rect 21774 2685 21834 17715
rect 21958 7581 22018 58787
rect 22691 34508 22757 34509
rect 22691 34444 22692 34508
rect 22756 34444 22757 34508
rect 22691 34443 22757 34444
rect 22139 24852 22205 24853
rect 22139 24788 22140 24852
rect 22204 24788 22205 24852
rect 22139 24787 22205 24788
rect 22142 10709 22202 24787
rect 22694 18053 22754 34443
rect 22691 18052 22757 18053
rect 22691 17988 22692 18052
rect 22756 17988 22757 18052
rect 22691 17987 22757 17988
rect 22875 14380 22941 14381
rect 22875 14316 22876 14380
rect 22940 14316 22941 14380
rect 22875 14315 22941 14316
rect 22139 10708 22205 10709
rect 22139 10644 22140 10708
rect 22204 10644 22205 10708
rect 22139 10643 22205 10644
rect 22323 10028 22389 10029
rect 22323 9964 22324 10028
rect 22388 9964 22389 10028
rect 22323 9963 22389 9964
rect 22326 8397 22386 9963
rect 22323 8396 22389 8397
rect 22323 8332 22324 8396
rect 22388 8332 22389 8396
rect 22323 8331 22389 8332
rect 21955 7580 22021 7581
rect 21955 7516 21956 7580
rect 22020 7516 22021 7580
rect 21955 7515 22021 7516
rect 22326 6901 22386 8331
rect 22323 6900 22389 6901
rect 22323 6836 22324 6900
rect 22388 6836 22389 6900
rect 22323 6835 22389 6836
rect 22326 4045 22386 6835
rect 22323 4044 22389 4045
rect 22323 3980 22324 4044
rect 22388 3980 22389 4044
rect 22323 3979 22389 3980
rect 22878 2685 22938 14315
rect 23062 9349 23122 59331
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 33915 56676 33981 56677
rect 33915 56612 33916 56676
rect 33980 56612 33981 56676
rect 33915 56611 33981 56612
rect 31155 52596 31221 52597
rect 31155 52532 31156 52596
rect 31220 52532 31221 52596
rect 31155 52531 31221 52532
rect 30235 47564 30301 47565
rect 30235 47500 30236 47564
rect 30300 47500 30301 47564
rect 30235 47499 30301 47500
rect 29867 41580 29933 41581
rect 29867 41516 29868 41580
rect 29932 41516 29933 41580
rect 29867 41515 29933 41516
rect 23795 38588 23861 38589
rect 23795 38524 23796 38588
rect 23860 38524 23861 38588
rect 23795 38523 23861 38524
rect 23243 36004 23309 36005
rect 23243 35940 23244 36004
rect 23308 35940 23309 36004
rect 23243 35939 23309 35940
rect 23059 9348 23125 9349
rect 23059 9284 23060 9348
rect 23124 9284 23125 9348
rect 23059 9283 23125 9284
rect 23246 8125 23306 35939
rect 23798 8533 23858 38523
rect 23979 23492 24045 23493
rect 23979 23428 23980 23492
rect 24044 23428 24045 23492
rect 23979 23427 24045 23428
rect 23982 9893 24042 23427
rect 24715 14244 24781 14245
rect 24715 14180 24716 14244
rect 24780 14180 24781 14244
rect 24715 14179 24781 14180
rect 23979 9892 24045 9893
rect 23979 9828 23980 9892
rect 24044 9828 24045 9892
rect 23979 9827 24045 9828
rect 23795 8532 23861 8533
rect 23795 8468 23796 8532
rect 23860 8468 23861 8532
rect 23795 8467 23861 8468
rect 23243 8124 23309 8125
rect 23243 8060 23244 8124
rect 23308 8060 23309 8124
rect 23243 8059 23309 8060
rect 24718 5133 24778 14179
rect 27107 13700 27173 13701
rect 27107 13636 27108 13700
rect 27172 13636 27173 13700
rect 27107 13635 27173 13636
rect 27110 12749 27170 13635
rect 27107 12748 27173 12749
rect 27107 12684 27108 12748
rect 27172 12684 27173 12748
rect 27107 12683 27173 12684
rect 29870 6901 29930 41515
rect 30238 8261 30298 47499
rect 30235 8260 30301 8261
rect 30235 8196 30236 8260
rect 30300 8196 30301 8260
rect 30235 8195 30301 8196
rect 31158 6901 31218 52531
rect 32811 51780 32877 51781
rect 32811 51716 32812 51780
rect 32876 51716 32877 51780
rect 32811 51715 32877 51716
rect 32814 6901 32874 51715
rect 33731 16284 33797 16285
rect 33731 16220 33732 16284
rect 33796 16220 33797 16284
rect 33731 16219 33797 16220
rect 33547 12612 33613 12613
rect 33547 12548 33548 12612
rect 33612 12548 33613 12612
rect 33547 12547 33613 12548
rect 33550 9621 33610 12547
rect 33547 9620 33613 9621
rect 33547 9556 33548 9620
rect 33612 9556 33613 9620
rect 33547 9555 33613 9556
rect 33550 8397 33610 9555
rect 33734 8397 33794 16219
rect 33547 8396 33613 8397
rect 33547 8332 33548 8396
rect 33612 8332 33613 8396
rect 33547 8331 33613 8332
rect 33731 8396 33797 8397
rect 33731 8332 33732 8396
rect 33796 8332 33797 8396
rect 33731 8331 33797 8332
rect 33918 8261 33978 56611
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 36123 53140 36189 53141
rect 36123 53076 36124 53140
rect 36188 53076 36189 53140
rect 36123 53075 36189 53076
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34651 42940 34717 42941
rect 34651 42876 34652 42940
rect 34716 42876 34717 42940
rect 34651 42875 34717 42876
rect 34099 26892 34165 26893
rect 34099 26828 34100 26892
rect 34164 26828 34165 26892
rect 34099 26827 34165 26828
rect 34102 9618 34162 26827
rect 34283 13564 34349 13565
rect 34283 13500 34284 13564
rect 34348 13500 34349 13564
rect 34283 13499 34349 13500
rect 34286 9890 34346 13499
rect 34467 11388 34533 11389
rect 34467 11324 34468 11388
rect 34532 11324 34533 11388
rect 34467 11323 34533 11324
rect 34470 10301 34530 11323
rect 34654 10437 34714 42875
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 35571 13836 35637 13837
rect 35571 13772 35572 13836
rect 35636 13772 35637 13836
rect 35571 13771 35637 13772
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34651 10436 34717 10437
rect 34651 10372 34652 10436
rect 34716 10372 34717 10436
rect 34651 10371 34717 10372
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34467 10300 34533 10301
rect 34467 10236 34468 10300
rect 34532 10236 34533 10300
rect 34467 10235 34533 10236
rect 34286 9830 34530 9890
rect 34470 9621 34530 9830
rect 34283 9620 34349 9621
rect 34283 9618 34284 9620
rect 34102 9558 34284 9618
rect 34283 9556 34284 9558
rect 34348 9556 34349 9620
rect 34283 9555 34349 9556
rect 34467 9620 34533 9621
rect 34467 9556 34468 9620
rect 34532 9556 34533 9620
rect 34467 9555 34533 9556
rect 34467 9348 34533 9349
rect 34467 9284 34468 9348
rect 34532 9284 34533 9348
rect 34467 9283 34533 9284
rect 33915 8260 33981 8261
rect 33915 8196 33916 8260
rect 33980 8196 33981 8260
rect 33915 8195 33981 8196
rect 29867 6900 29933 6901
rect 29867 6836 29868 6900
rect 29932 6836 29933 6900
rect 29867 6835 29933 6836
rect 31155 6900 31221 6901
rect 31155 6836 31156 6900
rect 31220 6836 31221 6900
rect 31155 6835 31221 6836
rect 32811 6900 32877 6901
rect 32811 6836 32812 6900
rect 32876 6836 32877 6900
rect 32811 6835 32877 6836
rect 24715 5132 24781 5133
rect 24715 5068 24716 5132
rect 24780 5068 24781 5132
rect 24715 5067 24781 5068
rect 34470 4725 34530 9283
rect 34928 9280 35248 10304
rect 35387 9620 35453 9621
rect 35387 9556 35388 9620
rect 35452 9556 35453 9620
rect 35387 9555 35453 9556
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34651 8260 34717 8261
rect 34651 8196 34652 8260
rect 34716 8196 34717 8260
rect 34651 8195 34717 8196
rect 34654 5949 34714 8195
rect 34928 8192 35248 9216
rect 35390 8669 35450 9555
rect 35387 8668 35453 8669
rect 35387 8604 35388 8668
rect 35452 8604 35453 8668
rect 35387 8603 35453 8604
rect 35574 8533 35634 13771
rect 36126 9621 36186 53075
rect 36859 50420 36925 50421
rect 36859 50356 36860 50420
rect 36924 50356 36925 50420
rect 36859 50355 36925 50356
rect 36675 26892 36741 26893
rect 36675 26828 36676 26892
rect 36740 26828 36741 26892
rect 36675 26827 36741 26828
rect 36307 26348 36373 26349
rect 36307 26284 36308 26348
rect 36372 26284 36373 26348
rect 36307 26283 36373 26284
rect 36310 10981 36370 26283
rect 36307 10980 36373 10981
rect 36307 10916 36308 10980
rect 36372 10916 36373 10980
rect 36307 10915 36373 10916
rect 36123 9620 36189 9621
rect 36123 9556 36124 9620
rect 36188 9556 36189 9620
rect 36123 9555 36189 9556
rect 36678 8533 36738 26827
rect 35571 8532 35637 8533
rect 35571 8468 35572 8532
rect 35636 8530 35637 8532
rect 36675 8532 36741 8533
rect 35636 8470 35818 8530
rect 35636 8468 35637 8470
rect 35571 8467 35637 8468
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34651 5948 34717 5949
rect 34651 5884 34652 5948
rect 34716 5884 34717 5948
rect 34651 5883 34717 5884
rect 34928 4928 35248 5952
rect 35758 5813 35818 8470
rect 36675 8468 36676 8532
rect 36740 8468 36741 8532
rect 36675 8467 36741 8468
rect 35755 5812 35821 5813
rect 35755 5748 35756 5812
rect 35820 5748 35821 5812
rect 35755 5747 35821 5748
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34467 4724 34533 4725
rect 34467 4660 34468 4724
rect 34532 4660 34533 4724
rect 34467 4659 34533 4660
rect 34928 3840 35248 4864
rect 36862 4045 36922 50355
rect 38515 50284 38581 50285
rect 38515 50220 38516 50284
rect 38580 50220 38581 50284
rect 38515 50219 38581 50220
rect 37227 16012 37293 16013
rect 37227 15948 37228 16012
rect 37292 15948 37293 16012
rect 37227 15947 37293 15948
rect 37230 13565 37290 15947
rect 37227 13564 37293 13565
rect 37227 13500 37228 13564
rect 37292 13500 37293 13564
rect 37227 13499 37293 13500
rect 38518 9621 38578 50219
rect 39254 11117 39314 61099
rect 50288 60960 50608 61520
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 42379 59396 42445 59397
rect 42379 59332 42380 59396
rect 42444 59332 42445 59396
rect 42379 59331 42445 59332
rect 40355 58036 40421 58037
rect 40355 57972 40356 58036
rect 40420 57972 40421 58036
rect 40355 57971 40421 57972
rect 39435 24172 39501 24173
rect 39435 24108 39436 24172
rect 39500 24108 39501 24172
rect 39435 24107 39501 24108
rect 39251 11116 39317 11117
rect 39251 11052 39252 11116
rect 39316 11052 39317 11116
rect 39251 11051 39317 11052
rect 38515 9620 38581 9621
rect 38515 9556 38516 9620
rect 38580 9556 38581 9620
rect 38515 9555 38581 9556
rect 38699 9484 38765 9485
rect 38699 9420 38700 9484
rect 38764 9420 38765 9484
rect 38699 9419 38765 9420
rect 38702 7989 38762 9419
rect 38699 7988 38765 7989
rect 38699 7924 38700 7988
rect 38764 7924 38765 7988
rect 38699 7923 38765 7924
rect 36859 4044 36925 4045
rect 36859 3980 36860 4044
rect 36924 3980 36925 4044
rect 36859 3979 36925 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 21035 2684 21101 2685
rect 21035 2620 21036 2684
rect 21100 2620 21101 2684
rect 21035 2619 21101 2620
rect 21771 2684 21837 2685
rect 21771 2620 21772 2684
rect 21836 2620 21837 2684
rect 21771 2619 21837 2620
rect 22875 2684 22941 2685
rect 22875 2620 22876 2684
rect 22940 2620 22941 2684
rect 22875 2619 22941 2620
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 39438 2685 39498 24107
rect 39803 19004 39869 19005
rect 39803 18940 39804 19004
rect 39868 18940 39869 19004
rect 39803 18939 39869 18940
rect 39806 9757 39866 18939
rect 40358 11389 40418 57971
rect 41827 47700 41893 47701
rect 41827 47636 41828 47700
rect 41892 47636 41893 47700
rect 41827 47635 41893 47636
rect 40723 22812 40789 22813
rect 40723 22748 40724 22812
rect 40788 22748 40789 22812
rect 40723 22747 40789 22748
rect 40539 20772 40605 20773
rect 40539 20708 40540 20772
rect 40604 20708 40605 20772
rect 40539 20707 40605 20708
rect 40355 11388 40421 11389
rect 40355 11324 40356 11388
rect 40420 11324 40421 11388
rect 40355 11323 40421 11324
rect 40171 11116 40237 11117
rect 40171 11052 40172 11116
rect 40236 11052 40237 11116
rect 40171 11051 40237 11052
rect 39987 10300 40053 10301
rect 39987 10236 39988 10300
rect 40052 10236 40053 10300
rect 39987 10235 40053 10236
rect 39803 9756 39869 9757
rect 39803 9692 39804 9756
rect 39868 9692 39869 9756
rect 39803 9691 39869 9692
rect 39990 8261 40050 10235
rect 40174 8261 40234 11051
rect 39987 8260 40053 8261
rect 39987 8196 39988 8260
rect 40052 8196 40053 8260
rect 39987 8195 40053 8196
rect 40171 8260 40237 8261
rect 40171 8196 40172 8260
rect 40236 8196 40237 8260
rect 40171 8195 40237 8196
rect 40542 4045 40602 20707
rect 40726 10437 40786 22747
rect 41275 22676 41341 22677
rect 41275 22612 41276 22676
rect 41340 22612 41341 22676
rect 41275 22611 41341 22612
rect 40723 10436 40789 10437
rect 40723 10372 40724 10436
rect 40788 10372 40789 10436
rect 40723 10371 40789 10372
rect 40539 4044 40605 4045
rect 40539 3980 40540 4044
rect 40604 3980 40605 4044
rect 40539 3979 40605 3980
rect 41278 2685 41338 22611
rect 41830 4045 41890 47635
rect 42382 5541 42442 59331
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 43483 57356 43549 57357
rect 43483 57292 43484 57356
rect 43548 57292 43549 57356
rect 43483 57291 43549 57292
rect 42931 42668 42997 42669
rect 42931 42604 42932 42668
rect 42996 42604 42997 42668
rect 42931 42603 42997 42604
rect 42379 5540 42445 5541
rect 42379 5476 42380 5540
rect 42444 5476 42445 5540
rect 42379 5475 42445 5476
rect 41827 4044 41893 4045
rect 41827 3980 41828 4044
rect 41892 3980 41893 4044
rect 41827 3979 41893 3980
rect 42934 2685 42994 42603
rect 43486 4045 43546 57291
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 43851 13836 43917 13837
rect 43851 13772 43852 13836
rect 43916 13772 43917 13836
rect 43851 13771 43917 13772
rect 43854 6901 43914 13771
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 43851 6900 43917 6901
rect 43851 6836 43852 6900
rect 43916 6836 43917 6900
rect 43851 6835 43917 6836
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 43483 4044 43549 4045
rect 43483 3980 43484 4044
rect 43548 3980 43549 4044
rect 43483 3979 43549 3980
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 39435 2684 39501 2685
rect 39435 2620 39436 2684
rect 39500 2620 39501 2684
rect 39435 2619 39501 2620
rect 41275 2684 41341 2685
rect 41275 2620 41276 2684
rect 41340 2620 41341 2684
rect 41275 2619 41341 2620
rect 42931 2684 42997 2685
rect 42931 2620 42932 2684
rect 42996 2620 42997 2684
rect 42931 2619 42997 2620
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 19379 780 19445 781
rect 19379 716 19380 780
rect 19444 716 19445 780
rect 19379 715 19445 716
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 32752 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 34868 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 33120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 34224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 35604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 20148 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 26404 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 28888 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 35880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 23000 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 17940 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 38180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 2300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 2300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 2300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 30636 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 29072 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 56580 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 40112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1676037725
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_144
timestamp 1676037725
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 1676037725
transform 1 0 14720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1676037725
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1676037725
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1676037725
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_292
timestamp 1676037725
transform 1 0 27968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1676037725
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1676037725
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1676037725
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1676037725
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_463
timestamp 1676037725
transform 1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 1676037725
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_490
timestamp 1676037725
transform 1 0 46184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1676037725
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1676037725
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_547
timestamp 1676037725
transform 1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1676037725
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 1676037725
transform 1 0 54372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_597
timestamp 1676037725
transform 1 0 56028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_607
timestamp 1676037725
transform 1 0 56948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1676037725
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1676037725
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1676037725
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1676037725
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1676037725
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1676037725
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1676037725
transform 1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1676037725
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1676037725
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_242
timestamp 1676037725
transform 1 0 23368 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1676037725
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_274
timestamp 1676037725
transform 1 0 26312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1676037725
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_303
timestamp 1676037725
transform 1 0 28980 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_311
timestamp 1676037725
transform 1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_322
timestamp 1676037725
transform 1 0 30728 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1676037725
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1676037725
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1676037725
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_383
timestamp 1676037725
transform 1 0 36340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_401
timestamp 1676037725
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1676037725
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_421
timestamp 1676037725
transform 1 0 39836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1676037725
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1676037725
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_481
timestamp 1676037725
transform 1 0 45356 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_489
timestamp 1676037725
transform 1 0 46092 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1676037725
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_513
timestamp 1676037725
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_523
timestamp 1676037725
transform 1 0 49220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_531
timestamp 1676037725
transform 1 0 49956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_539
timestamp 1676037725
transform 1 0 50692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_547
timestamp 1676037725
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1676037725
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_577
timestamp 1676037725
transform 1 0 54188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_587
timestamp 1676037725
transform 1 0 55108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_597
timestamp 1676037725
transform 1 0 56028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_607
timestamp 1676037725
transform 1 0 56948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1676037725
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1676037725
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1676037725
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1676037725
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1676037725
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1676037725
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1676037725
transform 1 0 20056 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1676037725
transform 1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1676037725
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1676037725
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1676037725
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_327
timestamp 1676037725
transform 1 0 31188 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_335
timestamp 1676037725
transform 1 0 31924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_352
timestamp 1676037725
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1676037725
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1676037725
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_405
timestamp 1676037725
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_437
timestamp 1676037725
transform 1 0 41308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1676037725
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1676037725
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_483
timestamp 1676037725
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_491
timestamp 1676037725
transform 1 0 46276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_495
timestamp 1676037725
transform 1 0 46644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_502
timestamp 1676037725
transform 1 0 47288 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1676037725
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_518
timestamp 1676037725
transform 1 0 48760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_526
timestamp 1676037725
transform 1 0 49496 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_539
timestamp 1676037725
transform 1 0 50692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1676037725
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1676037725
transform 1 0 52164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1676037725
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1676037725
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1676037725
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_595
timestamp 1676037725
transform 1 0 55844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_602
timestamp 1676037725
transform 1 0 56488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1676037725
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1676037725
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1676037725
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1676037725
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1676037725
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1676037725
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1676037725
transform 1 0 14536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_175
timestamp 1676037725
transform 1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1676037725
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1676037725
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1676037725
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1676037725
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_292
timestamp 1676037725
transform 1 0 27968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1676037725
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1676037725
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_348
timestamp 1676037725
transform 1 0 33120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_369
timestamp 1676037725
transform 1 0 35052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1676037725
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1676037725
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_399
timestamp 1676037725
transform 1 0 37812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1676037725
transform 1 0 38916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_419
timestamp 1676037725
transform 1 0 39652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_427
timestamp 1676037725
transform 1 0 40388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_435
timestamp 1676037725
transform 1 0 41124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1676037725
transform 1 0 41860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_465
timestamp 1676037725
transform 1 0 43884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_481
timestamp 1676037725
transform 1 0 45356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1676037725
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_511
timestamp 1676037725
transform 1 0 48116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_537
timestamp 1676037725
transform 1 0 50508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_542
timestamp 1676037725
transform 1 0 50968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_546
timestamp 1676037725
transform 1 0 51336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_551
timestamp 1676037725
transform 1 0 51796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_567
timestamp 1676037725
transform 1 0 53268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_575
timestamp 1676037725
transform 1 0 54004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_583
timestamp 1676037725
transform 1 0 54740 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_591
timestamp 1676037725
transform 1 0 55476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_603
timestamp 1676037725
transform 1 0 56580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_607
timestamp 1676037725
transform 1 0 56948 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1676037725
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1676037725
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1676037725
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1676037725
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1676037725
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_105
timestamp 1676037725
transform 1 0 10764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1676037725
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1676037725
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1676037725
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1676037725
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1676037725
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1676037725
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1676037725
transform 1 0 20056 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1676037725
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1676037725
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_240
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_290
timestamp 1676037725
transform 1 0 27784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_296
timestamp 1676037725
transform 1 0 28336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1676037725
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_341
timestamp 1676037725
transform 1 0 32476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1676037725
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1676037725
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_387
timestamp 1676037725
transform 1 0 36708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1676037725
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1676037725
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_411
timestamp 1676037725
transform 1 0 38916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_427
timestamp 1676037725
transform 1 0 40388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_435
timestamp 1676037725
transform 1 0 41124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_443
timestamp 1676037725
transform 1 0 41860 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_447
timestamp 1676037725
transform 1 0 42228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_468
timestamp 1676037725
transform 1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_483
timestamp 1676037725
transform 1 0 45540 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1676037725
transform 1 0 48668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 1676037725
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_579
timestamp 1676037725
transform 1 0 54372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1676037725
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_86
timestamp 1676037725
transform 1 0 9016 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_99
timestamp 1676037725
transform 1 0 10212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1676037725
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1676037725
transform 1 0 12880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1676037725
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1676037725
transform 1 0 14352 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_154
timestamp 1676037725
transform 1 0 15272 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1676037725
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp 1676037725
transform 1 0 18124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1676037725
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_239
timestamp 1676037725
transform 1 0 23092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1676037725
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_298
timestamp 1676037725
transform 1 0 28520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_325
timestamp 1676037725
transform 1 0 31004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1676037725
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_345
timestamp 1676037725
transform 1 0 32844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_355
timestamp 1676037725
transform 1 0 33764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_365
timestamp 1676037725
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_375
timestamp 1676037725
transform 1 0 35604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1676037725
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_399
timestamp 1676037725
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_407
timestamp 1676037725
transform 1 0 38548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_415
timestamp 1676037725
transform 1 0 39284 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_423
timestamp 1676037725
transform 1 0 40020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_431
timestamp 1676037725
transform 1 0 40756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_439
timestamp 1676037725
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_455
timestamp 1676037725
transform 1 0 42964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_463
timestamp 1676037725
transform 1 0 43700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_471
timestamp 1676037725
transform 1 0 44436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_479
timestamp 1676037725
transform 1 0 45172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_487
timestamp 1676037725
transform 1 0 45908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_612
timestamp 1676037725
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1676037725
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_107
timestamp 1676037725
transform 1 0 10948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1676037725
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_129
timestamp 1676037725
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1676037725
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_154
timestamp 1676037725
transform 1 0 15272 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_162
timestamp 1676037725
transform 1 0 16008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1676037725
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1676037725
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_216
timestamp 1676037725
transform 1 0 20976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_224
timestamp 1676037725
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1676037725
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1676037725
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_278
timestamp 1676037725
transform 1 0 26680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_282
timestamp 1676037725
transform 1 0 27048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_299
timestamp 1676037725
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_326
timestamp 1676037725
transform 1 0 31096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_334
timestamp 1676037725
transform 1 0 31832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_355
timestamp 1676037725
transform 1 0 33764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1676037725
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_384
timestamp 1676037725
transform 1 0 36432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1676037725
transform 1 0 37260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_397
timestamp 1676037725
transform 1 0 37628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_407
timestamp 1676037725
transform 1 0 38548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_415
timestamp 1676037725
transform 1 0 39284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_443
timestamp 1676037725
transform 1 0 41860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_458
timestamp 1676037725
transform 1 0 43240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_466
timestamp 1676037725
transform 1 0 43976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_482
timestamp 1676037725
transform 1 0 45448 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_494
timestamp 1676037725
transform 1 0 46552 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_506
timestamp 1676037725
transform 1 0 47656 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_518
timestamp 1676037725
transform 1 0 48760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_530
timestamp 1676037725
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_605
timestamp 1676037725
transform 1 0 56764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_622
timestamp 1676037725
transform 1 0 58328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_99
timestamp 1676037725
transform 1 0 10212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1676037725
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_119
timestamp 1676037725
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_131
timestamp 1676037725
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_143
timestamp 1676037725
transform 1 0 14260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_155
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_177
timestamp 1676037725
transform 1 0 17388 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_199
timestamp 1676037725
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_236
timestamp 1676037725
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_260
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_288
timestamp 1676037725
transform 1 0 27600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1676037725
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_313
timestamp 1676037725
transform 1 0 29900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_324
timestamp 1676037725
transform 1 0 30912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1676037725
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_356
timestamp 1676037725
transform 1 0 33856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_364
timestamp 1676037725
transform 1 0 34592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_376
timestamp 1676037725
transform 1 0 35696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1676037725
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_411
timestamp 1676037725
transform 1 0 38916 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_419
timestamp 1676037725
transform 1 0 39652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_431
timestamp 1676037725
transform 1 0 40756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_443
timestamp 1676037725
transform 1 0 41860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_453
timestamp 1676037725
transform 1 0 42780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_468
timestamp 1676037725
transform 1 0 44160 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_480
timestamp 1676037725
transform 1 0 45264 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_492
timestamp 1676037725
transform 1 0 46368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_593
timestamp 1676037725
transform 1 0 55660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_598
timestamp 1676037725
transform 1 0 56120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_611
timestamp 1676037725
transform 1 0 57316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1676037725
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1676037725
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1676037725
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1676037725
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1676037725
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_166
timestamp 1676037725
transform 1 0 16376 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_182
timestamp 1676037725
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_220
timestamp 1676037725
transform 1 0 21344 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1676037725
transform 1 0 23276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_262
timestamp 1676037725
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_282
timestamp 1676037725
transform 1 0 27048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1676037725
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_322
timestamp 1676037725
transform 1 0 30728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_347
timestamp 1676037725
transform 1 0 33028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1676037725
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_376
timestamp 1676037725
transform 1 0 35696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_386
timestamp 1676037725
transform 1 0 36616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_396
timestamp 1676037725
transform 1 0 37536 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_405
timestamp 1676037725
transform 1 0 38364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1676037725
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_426
timestamp 1676037725
transform 1 0 40296 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_432
timestamp 1676037725
transform 1 0 40848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_438
timestamp 1676037725
transform 1 0 41400 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_448
timestamp 1676037725
transform 1 0 42320 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_452
timestamp 1676037725
transform 1 0 42688 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_460
timestamp 1676037725
transform 1 0 43424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_470
timestamp 1676037725
transform 1 0 44344 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_605
timestamp 1676037725
transform 1 0 56764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 1676037725
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1676037725
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_94
timestamp 1676037725
transform 1 0 9752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_177
timestamp 1676037725
transform 1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1676037725
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_204
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_247
timestamp 1676037725
transform 1 0 23828 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_255
timestamp 1676037725
transform 1 0 24564 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_292
timestamp 1676037725
transform 1 0 27968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1676037725
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_319
timestamp 1676037725
transform 1 0 30452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_325
timestamp 1676037725
transform 1 0 31004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1676037725
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_348
timestamp 1676037725
transform 1 0 33120 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1676037725
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_377
timestamp 1676037725
transform 1 0 35788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1676037725
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_412
timestamp 1676037725
transform 1 0 39008 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_424
timestamp 1676037725
transform 1 0 40112 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_436
timestamp 1676037725
transform 1 0 41216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_454
timestamp 1676037725
transform 1 0 42872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_467
timestamp 1676037725
transform 1 0 44068 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1676037725
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1676037725
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_604
timestamp 1676037725
transform 1 0 56672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1676037725
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_622
timestamp 1676037725
transform 1 0 58328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1676037725
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_112
timestamp 1676037725
transform 1 0 11408 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1676037725
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1676037725
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1676037725
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_211
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_228
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1676037725
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1676037725
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_268
timestamp 1676037725
transform 1 0 25760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_285
timestamp 1676037725
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_298
timestamp 1676037725
transform 1 0 28520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1676037725
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_319
timestamp 1676037725
transform 1 0 30452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_347
timestamp 1676037725
transform 1 0 33028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_390
timestamp 1676037725
transform 1 0 36984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1676037725
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_414
timestamp 1676037725
transform 1 0 39192 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_426
timestamp 1676037725
transform 1 0 40296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_449
timestamp 1676037725
transform 1 0 42412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_470
timestamp 1676037725
transform 1 0 44344 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_597
timestamp 1676037725
transform 1 0 56028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1676037725
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_622
timestamp 1676037725
transform 1 0 58328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1676037725
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_179
timestamp 1676037725
transform 1 0 17572 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_239
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1676037725
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_292
timestamp 1676037725
transform 1 0 27968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_311
timestamp 1676037725
transform 1 0 29716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_328
timestamp 1676037725
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_346
timestamp 1676037725
transform 1 0 32936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_350
timestamp 1676037725
transform 1 0 33304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_358
timestamp 1676037725
transform 1 0 34040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_371
timestamp 1676037725
transform 1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1676037725
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1676037725
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_418
timestamp 1676037725
transform 1 0 39560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_422
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_431
timestamp 1676037725
transform 1 0 40756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_443
timestamp 1676037725
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_458
timestamp 1676037725
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_468
timestamp 1676037725
transform 1 0 44160 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_478
timestamp 1676037725
transform 1 0 45080 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_490
timestamp 1676037725
transform 1 0 46184 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_605
timestamp 1676037725
transform 1 0 56764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1676037725
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1676037725
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1676037725
transform 1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_179
timestamp 1676037725
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1676037725
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1676037725
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1676037725
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1676037725
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_298
timestamp 1676037725
transform 1 0 28520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_302
timestamp 1676037725
transform 1 0 28888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_341
timestamp 1676037725
transform 1 0 32476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_352
timestamp 1676037725
transform 1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1676037725
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_373
timestamp 1676037725
transform 1 0 35420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1676037725
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_409
timestamp 1676037725
transform 1 0 38732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_426
timestamp 1676037725
transform 1 0 40296 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_468
timestamp 1676037725
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_601
timestamp 1676037725
transform 1 0 56396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_607
timestamp 1676037725
transform 1 0 56948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_611
timestamp 1676037725
transform 1 0 57316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_623
timestamp 1676037725
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_121
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1676037725
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1676037725
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1676037725
transform 1 0 19412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_243
timestamp 1676037725
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1676037725
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_299
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_312
timestamp 1676037725
transform 1 0 29808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_323
timestamp 1676037725
transform 1 0 30820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_345
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_353
timestamp 1676037725
transform 1 0 33580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_372
timestamp 1676037725
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_383
timestamp 1676037725
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_397
timestamp 1676037725
transform 1 0 37628 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_407
timestamp 1676037725
transform 1 0 38548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_415
timestamp 1676037725
transform 1 0 39284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_427
timestamp 1676037725
transform 1 0 40388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1676037725
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_468
timestamp 1676037725
transform 1 0 44160 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_481
timestamp 1676037725
transform 1 0 45356 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_493
timestamp 1676037725
transform 1 0 46460 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_501
timestamp 1676037725
transform 1 0 47196 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_597
timestamp 1676037725
transform 1 0 56028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1676037725
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1676037725
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1676037725
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_117
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1676037725
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_157
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1676037725
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1676037725
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1676037725
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1676037725
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_320
timestamp 1676037725
transform 1 0 30544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_354
timestamp 1676037725
transform 1 0 33672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_374
timestamp 1676037725
transform 1 0 35512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_378
timestamp 1676037725
transform 1 0 35880 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_386
timestamp 1676037725
transform 1 0 36616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_390
timestamp 1676037725
transform 1 0 36984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_407
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1676037725
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_425
timestamp 1676037725
transform 1 0 40204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_434
timestamp 1676037725
transform 1 0 41032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_463
timestamp 1676037725
transform 1 0 43700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1676037725
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1676037725
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1676037725
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1676037725
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1676037725
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1676037725
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1676037725
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1676037725
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_601
timestamp 1676037725
transform 1 0 56396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_605
timestamp 1676037725
transform 1 0 56764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_622
timestamp 1676037725
transform 1 0 58328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1676037725
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_239
timestamp 1676037725
transform 1 0 23092 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_272
timestamp 1676037725
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_287
timestamp 1676037725
transform 1 0 27508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_346
timestamp 1676037725
transform 1 0 32936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_350
timestamp 1676037725
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_358
timestamp 1676037725
transform 1 0 34040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_377
timestamp 1676037725
transform 1 0 35788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_404
timestamp 1676037725
transform 1 0 38272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_413
timestamp 1676037725
transform 1 0 39100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_420
timestamp 1676037725
transform 1 0 39744 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_434
timestamp 1676037725
transform 1 0 41032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1676037725
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_460
timestamp 1676037725
transform 1 0 43424 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1676037725
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_545
timestamp 1676037725
transform 1 0 51244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_557
timestamp 1676037725
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1676037725
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1676037725
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1676037725
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_609
timestamp 1676037725
transform 1 0 57132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_613
timestamp 1676037725
transform 1 0 57500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1676037725
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1676037725
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_354
timestamp 1676037725
transform 1 0 33672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_386
timestamp 1676037725
transform 1 0 36616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1676037725
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_404
timestamp 1676037725
transform 1 0 38272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_434
timestamp 1676037725
transform 1 0 41032 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_440
timestamp 1676037725
transform 1 0 41584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_461
timestamp 1676037725
transform 1 0 43516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1676037725
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1676037725
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1676037725
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_557
timestamp 1676037725
transform 1 0 52348 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_567
timestamp 1676037725
transform 1 0 53268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_579
timestamp 1676037725
transform 1 0 54372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1676037725
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1676037725
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1676037725
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_613
timestamp 1676037725
transform 1 0 57500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_623
timestamp 1676037725
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_122
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_134
timestamp 1676037725
transform 1 0 13432 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1676037725
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1676037725
transform 1 0 18768 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_243
timestamp 1676037725
transform 1 0 23460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1676037725
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1676037725
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1676037725
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1676037725
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1676037725
transform 1 0 32844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_354
timestamp 1676037725
transform 1 0 33672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_367
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_377
timestamp 1676037725
transform 1 0 35788 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_411
timestamp 1676037725
transform 1 0 38916 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_418
timestamp 1676037725
transform 1 0 39560 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_440
timestamp 1676037725
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_468
timestamp 1676037725
transform 1 0 44160 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_480
timestamp 1676037725
transform 1 0 45264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_492
timestamp 1676037725
transform 1 0 46368 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1676037725
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1676037725
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1676037725
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1676037725
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1676037725
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1676037725
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1676037725
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1676037725
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1676037725
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1676037725
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_617
timestamp 1676037725
transform 1 0 57868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1676037725
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1676037725
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp 1676037725
transform 1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_281
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1676037725
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_343
timestamp 1676037725
transform 1 0 32660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_347
timestamp 1676037725
transform 1 0 33028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_386
timestamp 1676037725
transform 1 0 36616 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_394
timestamp 1676037725
transform 1 0 37352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_405
timestamp 1676037725
transform 1 0 38364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_414
timestamp 1676037725
transform 1 0 39192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_430
timestamp 1676037725
transform 1 0 40664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_438
timestamp 1676037725
transform 1 0 41400 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_458
timestamp 1676037725
transform 1 0 43240 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_470
timestamp 1676037725
transform 1 0 44344 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1676037725
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1676037725
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1676037725
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1676037725
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1676037725
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1676037725
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1676037725
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1676037725
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1676037725
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1676037725
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1676037725
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1676037725
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1676037725
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_188
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1676037725
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_320
timestamp 1676037725
transform 1 0 30544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1676037725
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_346
timestamp 1676037725
transform 1 0 32936 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_354
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_414
timestamp 1676037725
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_426
timestamp 1676037725
transform 1 0 40296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_437
timestamp 1676037725
transform 1 0 41308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1676037725
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_460
timestamp 1676037725
transform 1 0 43424 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_472
timestamp 1676037725
transform 1 0 44528 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_484
timestamp 1676037725
transform 1 0 45632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_496
timestamp 1676037725
transform 1 0 46736 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1676037725
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1676037725
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1676037725
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1676037725
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1676037725
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1676037725
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1676037725
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1676037725
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1676037725
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1676037725
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1676037725
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1676037725
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_152
timestamp 1676037725
transform 1 0 15088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_216
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_320
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_326
timestamp 1676037725
transform 1 0 31096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_347
timestamp 1676037725
transform 1 0 33028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_358
timestamp 1676037725
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_369
timestamp 1676037725
transform 1 0 35052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_396
timestamp 1676037725
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_404
timestamp 1676037725
transform 1 0 38272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_414
timestamp 1676037725
transform 1 0 39192 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_430
timestamp 1676037725
transform 1 0 40664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_441
timestamp 1676037725
transform 1 0 41676 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_448
timestamp 1676037725
transform 1 0 42320 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_460
timestamp 1676037725
transform 1 0 43424 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1676037725
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1676037725
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1676037725
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1676037725
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1676037725
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1676037725
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1676037725
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1676037725
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1676037725
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_601
timestamp 1676037725
transform 1 0 56396 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1676037725
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1676037725
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1676037725
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1676037725
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_190
timestamp 1676037725
transform 1 0 18584 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_248
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_309
timestamp 1676037725
transform 1 0 29532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_364
timestamp 1676037725
transform 1 0 34592 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_401
timestamp 1676037725
transform 1 0 37996 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_409
timestamp 1676037725
transform 1 0 38732 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_427
timestamp 1676037725
transform 1 0 40388 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_435
timestamp 1676037725
transform 1 0 41124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1676037725
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_457
timestamp 1676037725
transform 1 0 43148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_462
timestamp 1676037725
transform 1 0 43608 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_475
timestamp 1676037725
transform 1 0 44804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1676037725
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_512
timestamp 1676037725
transform 1 0 48208 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_524
timestamp 1676037725
transform 1 0 49312 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_536
timestamp 1676037725
transform 1 0 50416 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_548
timestamp 1676037725
transform 1 0 51520 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1676037725
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1676037725
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1676037725
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1676037725
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1676037725
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1676037725
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1676037725
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1676037725
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_216
timestamp 1676037725
transform 1 0 20976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_302
timestamp 1676037725
transform 1 0 28888 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1676037725
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_347
timestamp 1676037725
transform 1 0 33028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_376
timestamp 1676037725
transform 1 0 35696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_396
timestamp 1676037725
transform 1 0 37536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_400
timestamp 1676037725
transform 1 0 37904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_431
timestamp 1676037725
transform 1 0 40756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_440
timestamp 1676037725
transform 1 0 41584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_444
timestamp 1676037725
transform 1 0 41952 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_454
timestamp 1676037725
transform 1 0 42872 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_462
timestamp 1676037725
transform 1 0 43608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_497
timestamp 1676037725
transform 1 0 46828 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_517
timestamp 1676037725
transform 1 0 48668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_529
timestamp 1676037725
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1676037725
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1676037725
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1676037725
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1676037725
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1676037725
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1676037725
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1676037725
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1676037725
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1676037725
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1676037725
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1676037725
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_192
timestamp 1676037725
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1676037725
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_370
timestamp 1676037725
transform 1 0 35144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1676037725
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_400
timestamp 1676037725
transform 1 0 37904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_408
timestamp 1676037725
transform 1 0 38640 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_419
timestamp 1676037725
transform 1 0 39652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_427
timestamp 1676037725
transform 1 0 40388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_457
timestamp 1676037725
transform 1 0 43148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_467
timestamp 1676037725
transform 1 0 44068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_487
timestamp 1676037725
transform 1 0 45908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_513
timestamp 1676037725
transform 1 0 48300 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_531
timestamp 1676037725
transform 1 0 49956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_543
timestamp 1676037725
transform 1 0 51060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_555
timestamp 1676037725
transform 1 0 52164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1676037725
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1676037725
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1676037725
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1676037725
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1676037725
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1676037725
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1676037725
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1676037725
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1676037725
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1676037725
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1676037725
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1676037725
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1676037725
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_326
timestamp 1676037725
transform 1 0 31096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_346
timestamp 1676037725
transform 1 0 32936 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1676037725
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1676037725
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_390
timestamp 1676037725
transform 1 0 36984 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_404
timestamp 1676037725
transform 1 0 38272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1676037725
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_428
timestamp 1676037725
transform 1 0 40480 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_460
timestamp 1676037725
transform 1 0 43424 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1676037725
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_486
timestamp 1676037725
transform 1 0 45816 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_494
timestamp 1676037725
transform 1 0 46552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_528
timestamp 1676037725
transform 1 0 49680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_533
timestamp 1676037725
transform 1 0 50140 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_540
timestamp 1676037725
transform 1 0 50784 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_552
timestamp 1676037725
transform 1 0 51888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_564
timestamp 1676037725
transform 1 0 52992 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_576
timestamp 1676037725
transform 1 0 54096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1676037725
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1676037725
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1676037725
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1676037725
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1676037725
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_136
timestamp 1676037725
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1676037725
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_356
timestamp 1676037725
transform 1 0 33856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_376
timestamp 1676037725
transform 1 0 35696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1676037725
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_412
timestamp 1676037725
transform 1 0 39008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_421
timestamp 1676037725
transform 1 0 39836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_430
timestamp 1676037725
transform 1 0 40664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_436
timestamp 1676037725
transform 1 0 41216 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1676037725
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_453
timestamp 1676037725
transform 1 0 42780 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_482
timestamp 1676037725
transform 1 0 45448 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_495
timestamp 1676037725
transform 1 0 46644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_518
timestamp 1676037725
transform 1 0 48760 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_527
timestamp 1676037725
transform 1 0 49588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_539
timestamp 1676037725
transform 1 0 50692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_551
timestamp 1676037725
transform 1 0 51796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1676037725
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1676037725
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1676037725
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1676037725
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1676037725
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1676037725
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1676037725
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1676037725
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1676037725
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1676037725
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1676037725
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_272
timestamp 1676037725
transform 1 0 26128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_327
timestamp 1676037725
transform 1 0 31188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1676037725
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_376
timestamp 1676037725
transform 1 0 35696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_380
timestamp 1676037725
transform 1 0 36064 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 1676037725
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_411
timestamp 1676037725
transform 1 0 38916 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_434
timestamp 1676037725
transform 1 0 41032 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_443
timestamp 1676037725
transform 1 0 41860 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_451
timestamp 1676037725
transform 1 0 42596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_459
timestamp 1676037725
transform 1 0 43332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_470
timestamp 1676037725
transform 1 0 44344 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_484
timestamp 1676037725
transform 1 0 45632 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_496
timestamp 1676037725
transform 1 0 46736 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_509
timestamp 1676037725
transform 1 0 47932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_530
timestamp 1676037725
transform 1 0 49864 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1676037725
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1676037725
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1676037725
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1676037725
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1676037725
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1676037725
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1676037725
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_601
timestamp 1676037725
transform 1 0 56396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1676037725
transform 1 0 57500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_623
timestamp 1676037725
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1676037725
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1676037725
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_263
timestamp 1676037725
transform 1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_288
timestamp 1676037725
transform 1 0 27600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_318
timestamp 1676037725
transform 1 0 30360 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_324
timestamp 1676037725
transform 1 0 30912 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_341
timestamp 1676037725
transform 1 0 32476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_368
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_381
timestamp 1676037725
transform 1 0 36156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1676037725
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_400
timestamp 1676037725
transform 1 0 37904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_422
timestamp 1676037725
transform 1 0 39928 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_435
timestamp 1676037725
transform 1 0 41124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1676037725
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_459
timestamp 1676037725
transform 1 0 43332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_467
timestamp 1676037725
transform 1 0 44068 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_513
timestamp 1676037725
transform 1 0 48300 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_532
timestamp 1676037725
transform 1 0 50048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_544
timestamp 1676037725
transform 1 0 51152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_556
timestamp 1676037725
transform 1 0 52256 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1676037725
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1676037725
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1676037725
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1676037725
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1676037725
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1676037725
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1676037725
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1676037725
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_150
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1676037725
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_216
timestamp 1676037725
transform 1 0 20976 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1676037725
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_292
timestamp 1676037725
transform 1 0 27968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_296
timestamp 1676037725
transform 1 0 28336 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_343
timestamp 1676037725
transform 1 0 32660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_356
timestamp 1676037725
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_373
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1676037725
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1676037725
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_440
timestamp 1676037725
transform 1 0 41584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_444
timestamp 1676037725
transform 1 0 41952 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_450
timestamp 1676037725
transform 1 0 42504 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_471
timestamp 1676037725
transform 1 0 44436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_486
timestamp 1676037725
transform 1 0 45816 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_498
timestamp 1676037725
transform 1 0 46920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_507
timestamp 1676037725
transform 1 0 47748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_528
timestamp 1676037725
transform 1 0 49680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_533
timestamp 1676037725
transform 1 0 50140 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_552
timestamp 1676037725
transform 1 0 51888 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_564
timestamp 1676037725
transform 1 0 52992 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_576
timestamp 1676037725
transform 1 0 54096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1676037725
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1676037725
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1676037725
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_267
timestamp 1676037725
transform 1 0 25668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_291
timestamp 1676037725
transform 1 0 27876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_321
timestamp 1676037725
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_365
timestamp 1676037725
transform 1 0 34684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1676037725
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_408
timestamp 1676037725
transform 1 0 38640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_426
timestamp 1676037725
transform 1 0 40296 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_439
timestamp 1676037725
transform 1 0 41492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1676037725
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_453
timestamp 1676037725
transform 1 0 42780 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_471
timestamp 1676037725
transform 1 0 44436 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_479
timestamp 1676037725
transform 1 0 45172 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_499
timestamp 1676037725
transform 1 0 47012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_528
timestamp 1676037725
transform 1 0 49680 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_537
timestamp 1676037725
transform 1 0 50508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_549
timestamp 1676037725
transform 1 0 51612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_557
timestamp 1676037725
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1676037725
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1676037725
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1676037725
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1676037725
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1676037725
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1676037725
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_617
timestamp 1676037725
transform 1 0 57868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1676037725
transform 1 0 58420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_203
timestamp 1676037725
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_272
timestamp 1676037725
transform 1 0 26128 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_315
timestamp 1676037725
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_325
timestamp 1676037725
transform 1 0 31004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_355
timestamp 1676037725
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1676037725
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_372
timestamp 1676037725
transform 1 0 35328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_376
timestamp 1676037725
transform 1 0 35696 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1676037725
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_416
timestamp 1676037725
transform 1 0 39376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_426
timestamp 1676037725
transform 1 0 40296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_458
timestamp 1676037725
transform 1 0 43240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_486
timestamp 1676037725
transform 1 0 45816 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_498
timestamp 1676037725
transform 1 0 46920 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_506
timestamp 1676037725
transform 1 0 47656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_515
timestamp 1676037725
transform 1 0 48484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_526
timestamp 1676037725
transform 1 0 49496 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1676037725
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1676037725
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1676037725
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1676037725
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1676037725
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1676037725
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1676037725
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1676037725
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1676037725
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1676037725
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_248
timestamp 1676037725
transform 1 0 23920 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1676037725
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_378
timestamp 1676037725
transform 1 0 35880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_421
timestamp 1676037725
transform 1 0 39836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_426
timestamp 1676037725
transform 1 0 40296 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_437
timestamp 1676037725
transform 1 0 41308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1676037725
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_457
timestamp 1676037725
transform 1 0 43148 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_469
timestamp 1676037725
transform 1 0 44252 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_481
timestamp 1676037725
transform 1 0 45356 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_493
timestamp 1676037725
transform 1 0 46460 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_501
timestamp 1676037725
transform 1 0 47196 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_515
timestamp 1676037725
transform 1 0 48484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_524
timestamp 1676037725
transform 1 0 49312 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_536
timestamp 1676037725
transform 1 0 50416 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_548
timestamp 1676037725
transform 1 0 51520 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1676037725
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1676037725
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1676037725
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1676037725
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1676037725
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1676037725
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_617
timestamp 1676037725
transform 1 0 57868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1676037725
transform 1 0 58420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1676037725
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_220
timestamp 1676037725
transform 1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_263
timestamp 1676037725
transform 1 0 25300 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_271
timestamp 1676037725
transform 1 0 26036 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1676037725
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_354
timestamp 1676037725
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_383
timestamp 1676037725
transform 1 0 36340 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1676037725
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1676037725
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_427
timestamp 1676037725
transform 1 0 40388 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_509
timestamp 1676037725
transform 1 0 47932 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_516
timestamp 1676037725
transform 1 0 48576 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_528
timestamp 1676037725
transform 1 0 49680 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1676037725
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1676037725
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1676037725
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1676037725
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1676037725
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1676037725
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1676037725
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1676037725
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1676037725
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_623
timestamp 1676037725
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1676037725
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_194
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp 1676037725
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_270
timestamp 1676037725
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_290
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_296
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_314
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_344
timestamp 1676037725
transform 1 0 32752 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_356
timestamp 1676037725
transform 1 0 33856 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_368
timestamp 1676037725
transform 1 0 34960 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_380
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_412
timestamp 1676037725
transform 1 0 39008 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_424
timestamp 1676037725
transform 1 0 40112 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_436
timestamp 1676037725
transform 1 0 41216 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1676037725
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1676037725
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1676037725
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1676037725
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1676037725
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1676037725
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1676037725
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1676037725
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1676037725
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1676037725
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1676037725
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_205
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1676037725
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1676037725
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_283
timestamp 1676037725
transform 1 0 27140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1676037725
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_320
timestamp 1676037725
transform 1 0 30544 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_324
timestamp 1676037725
transform 1 0 30912 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_336
timestamp 1676037725
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_348
timestamp 1676037725
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1676037725
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1676037725
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1676037725
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1676037725
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1676037725
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1676037725
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1676037725
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1676037725
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1676037725
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1676037725
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1676037725
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_213
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1676037725
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1676037725
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_308
timestamp 1676037725
transform 1 0 29440 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_320
timestamp 1676037725
transform 1 0 30544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1676037725
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1676037725
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1676037725
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1676037725
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1676037725
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1676037725
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1676037725
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1676037725
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1676037725
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1676037725
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1676037725
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1676037725
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_11
timestamp 1676037725
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1676037725
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_184
timestamp 1676037725
transform 1 0 18032 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1676037725
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1676037725
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1676037725
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1676037725
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1676037725
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1676037725
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1676037725
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1676037725
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1676037725
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1676037725
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1676037725
transform 1 0 57500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_623
timestamp 1676037725
transform 1 0 58420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_11
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_23
timestamp 1676037725
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1676037725
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_184
timestamp 1676037725
transform 1 0 18032 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_196
timestamp 1676037725
transform 1 0 19136 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_208
timestamp 1676037725
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_233
timestamp 1676037725
transform 1 0 22540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1676037725
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1676037725
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_288
timestamp 1676037725
transform 1 0 27600 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_300
timestamp 1676037725
transform 1 0 28704 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_312
timestamp 1676037725
transform 1 0 29808 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_324
timestamp 1676037725
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1676037725
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1676037725
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1676037725
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1676037725
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1676037725
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1676037725
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1676037725
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1676037725
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1676037725
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1676037725
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1676037725
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1676037725
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1676037725
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_183
timestamp 1676037725
transform 1 0 17940 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1676037725
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1676037725
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_280
timestamp 1676037725
transform 1 0 26864 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_292
timestamp 1676037725
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1676037725
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1676037725
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1676037725
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1676037725
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1676037725
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1676037725
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1676037725
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1676037725
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1676037725
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1676037725
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_623
timestamp 1676037725
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_176
timestamp 1676037725
transform 1 0 17296 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_200
timestamp 1676037725
transform 1 0 19504 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1676037725
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1676037725
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1676037725
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1676037725
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1676037725
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1676037725
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1676037725
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1676037725
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1676037725
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1676037725
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1676037725
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_11
timestamp 1676037725
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1676037725
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_36
timestamp 1676037725
transform 1 0 4416 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_48
timestamp 1676037725
transform 1 0 5520 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_60
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_72
timestamp 1676037725
transform 1 0 7728 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1676037725
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1676037725
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1676037725
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1676037725
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1676037725
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1676037725
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1676037725
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1676037725
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1676037725
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1676037725
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1676037725
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1676037725
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1676037725
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_23
timestamp 1676037725
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_35
timestamp 1676037725
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1676037725
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1676037725
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1676037725
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1676037725
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1676037725
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1676037725
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1676037725
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1676037725
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1676037725
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1676037725
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1676037725
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1676037725
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1676037725
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1676037725
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1676037725
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1676037725
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1676037725
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1676037725
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1676037725
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1676037725
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1676037725
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1676037725
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1676037725
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1676037725
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1676037725
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1676037725
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1676037725
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1676037725
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1676037725
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1676037725
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1676037725
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1676037725
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1676037725
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1676037725
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1676037725
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1676037725
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1676037725
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_189
timestamp 1676037725
transform 1 0 18492 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_201
timestamp 1676037725
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1676037725
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1676037725
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1676037725
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1676037725
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1676037725
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1676037725
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1676037725
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1676037725
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1676037725
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1676037725
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1676037725
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1676037725
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1676037725
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1676037725
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1676037725
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1676037725
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1676037725
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1676037725
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1676037725
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1676037725
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1676037725
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1676037725
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1676037725
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1676037725
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1676037725
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_601
timestamp 1676037725
transform 1 0 56396 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1676037725
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1676037725
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1676037725
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1676037725
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1676037725
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1676037725
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1676037725
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1676037725
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1676037725
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1676037725
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1676037725
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1676037725
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1676037725
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1676037725
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1676037725
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1676037725
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1676037725
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1676037725
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1676037725
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1676037725
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1676037725
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_11
timestamp 1676037725
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1676037725
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1676037725
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1676037725
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1676037725
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1676037725
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1676037725
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1676037725
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1676037725
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1676037725
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1676037725
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1676037725
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_11
timestamp 1676037725
transform 1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1676037725
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1676037725
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1676037725
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1676037725
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1676037725
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1676037725
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1676037725
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1676037725
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1676037725
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1676037725
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1676037725
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1676037725
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1676037725
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_617
timestamp 1676037725
transform 1 0 57868 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1676037725
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_11
timestamp 1676037725
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1676037725
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1676037725
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1676037725
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1676037725
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1676037725
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1676037725
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1676037725
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1676037725
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1676037725
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1676037725
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1676037725
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1676037725
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_177
timestamp 1676037725
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_187
timestamp 1676037725
transform 1 0 18308 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_199
timestamp 1676037725
transform 1 0 19412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_211
timestamp 1676037725
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_265
timestamp 1676037725
transform 1 0 25484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1676037725
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1676037725
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1676037725
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1676037725
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1676037725
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1676037725
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1676037725
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1676037725
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1676037725
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1676037725
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1676037725
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1676037725
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_11
timestamp 1676037725
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1676037725
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_241
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1676037725
transform 1 0 25208 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_275
timestamp 1676037725
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_287
timestamp 1676037725
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_299
timestamp 1676037725
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1676037725
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1676037725
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1676037725
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1676037725
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1676037725
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1676037725
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1676037725
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1676037725
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_601
timestamp 1676037725
transform 1 0 56396 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1676037725
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1676037725
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_11
timestamp 1676037725
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_23
timestamp 1676037725
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1676037725
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1676037725
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_250
timestamp 1676037725
transform 1 0 24104 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_258
timestamp 1676037725
transform 1 0 24840 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_268
timestamp 1676037725
transform 1 0 25760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1676037725
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1676037725
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1676037725
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1676037725
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1676037725
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1676037725
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1676037725
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1676037725
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1676037725
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1676037725
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1676037725
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1676037725
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1676037725
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_207
timestamp 1676037725
transform 1 0 20148 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_219
timestamp 1676037725
transform 1 0 21252 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_231
timestamp 1676037725
transform 1 0 22356 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1676037725
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1676037725
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1676037725
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1676037725
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1676037725
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1676037725
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1676037725
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1676037725
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1676037725
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1676037725
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1676037725
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_9
timestamp 1676037725
transform 1 0 1932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1676037725
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1676037725
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1676037725
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1676037725
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1676037725
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1676037725
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1676037725
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1676037725
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1676037725
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1676037725
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1676037725
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1676037725
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 1676037725
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1676037725
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_261
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_270
timestamp 1676037725
transform 1 0 25944 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_282
timestamp 1676037725
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_294
timestamp 1676037725
transform 1 0 28152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1676037725
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1676037725
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1676037725
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1676037725
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1676037725
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1676037725
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1676037725
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1676037725
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1676037725
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1676037725
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1676037725
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1676037725
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1676037725
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1676037725
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1676037725
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1676037725
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1676037725
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1676037725
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1676037725
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1676037725
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1676037725
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1676037725
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1676037725
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1676037725
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1676037725
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1676037725
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1676037725
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_229
timestamp 1676037725
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1676037725
transform 1 0 23276 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1676037725
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_287
timestamp 1676037725
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1676037725
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1676037725
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1676037725
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1676037725
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1676037725
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1676037725
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1676037725
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1676037725
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1676037725
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_601
timestamp 1676037725
transform 1 0 56396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1676037725
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1676037725
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1676037725
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_236
timestamp 1676037725
transform 1 0 22816 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_248
timestamp 1676037725
transform 1 0 23920 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_260
timestamp 1676037725
transform 1 0 25024 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_272
timestamp 1676037725
transform 1 0 26128 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1676037725
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1676037725
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1676037725
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1676037725
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1676037725
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1676037725
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1676037725
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1676037725
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1676037725
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1676037725
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1676037725
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_213
timestamp 1676037725
transform 1 0 20700 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1676037725
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_236
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1676037725
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1676037725
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1676037725
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1676037725
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1676037725
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1676037725
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1676037725
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1676037725
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1676037725
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1676037725
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1676037725
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1676037725
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_236
timestamp 1676037725
transform 1 0 22816 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_240
timestamp 1676037725
transform 1 0 23184 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_261
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_269
timestamp 1676037725
transform 1 0 25852 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1676037725
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1676037725
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1676037725
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1676037725
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1676037725
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1676037725
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1676037725
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1676037725
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1676037725
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1676037725
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1676037725
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1676037725
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1676037725
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1676037725
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_207
timestamp 1676037725
transform 1 0 20148 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_211
timestamp 1676037725
transform 1 0 20516 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_232
timestamp 1676037725
transform 1 0 22448 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 1676037725
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_391
timestamp 1676037725
transform 1 0 37076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_403
timestamp 1676037725
transform 1 0 38180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_415
timestamp 1676037725
transform 1 0 39284 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_430
timestamp 1676037725
transform 1 0 40664 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_442
timestamp 1676037725
transform 1 0 41768 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_454
timestamp 1676037725
transform 1 0 42872 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_466
timestamp 1676037725
transform 1 0 43976 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_474
timestamp 1676037725
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1676037725
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1676037725
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1676037725
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1676037725
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1676037725
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1676037725
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1676037725
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1676037725
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1676037725
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1676037725
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1676037725
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_9
timestamp 1676037725
transform 1 0 1932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_21
timestamp 1676037725
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1676037725
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1676037725
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_207
timestamp 1676037725
transform 1 0 20148 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1676037725
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_243
timestamp 1676037725
transform 1 0 23460 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_253
timestamp 1676037725
transform 1 0 24380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_265
timestamp 1676037725
transform 1 0 25484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1676037725
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1676037725
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1676037725
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1676037725
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1676037725
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1676037725
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1676037725
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1676037725
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1676037725
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1676037725
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1676037725
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1676037725
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_9
timestamp 1676037725
transform 1 0 1932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 1676037725
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_60
timestamp 1676037725
transform 1 0 6624 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_72
timestamp 1676037725
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_185
timestamp 1676037725
transform 1 0 18124 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_213
timestamp 1676037725
transform 1 0 20700 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_226
timestamp 1676037725
transform 1 0 21896 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_239
timestamp 1676037725
transform 1 0 23092 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_425
timestamp 1676037725
transform 1 0 40204 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1676037725
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1676037725
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1676037725
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1676037725
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_577
timestamp 1676037725
transform 1 0 54188 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_585
timestamp 1676037725
transform 1 0 54924 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1676037725
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1676037725
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1676037725
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1676037725
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_9
timestamp 1676037725
transform 1 0 1932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1676037725
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_25
timestamp 1676037725
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_37
timestamp 1676037725
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1676037725
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_67
timestamp 1676037725
transform 1 0 7268 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_79
timestamp 1676037725
transform 1 0 8372 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_91
timestamp 1676037725
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1676037725
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_188
timestamp 1676037725
transform 1 0 18400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_199
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1676037725
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_241
timestamp 1676037725
transform 1 0 23276 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_254
timestamp 1676037725
transform 1 0 24472 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_266
timestamp 1676037725
transform 1 0 25576 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1676037725
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1676037725
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1676037725
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1676037725
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1676037725
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_561
timestamp 1676037725
transform 1 0 52716 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_569
timestamp 1676037725
transform 1 0 53452 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1676037725
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1676037725
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1676037725
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1676037725
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1676037725
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1676037725
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_17
timestamp 1676037725
transform 1 0 2668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1676037725
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_185
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1676037725
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_215
timestamp 1676037725
transform 1 0 20884 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_227
timestamp 1676037725
transform 1 0 21988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_239
timestamp 1676037725
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1676037725
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1676037725
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1676037725
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1676037725
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1676037725
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1676037725
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1676037725
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1676037725
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1676037725
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1676037725
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1676037725
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_9
timestamp 1676037725
transform 1 0 1932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_21
timestamp 1676037725
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_45
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 1676037725
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_209
timestamp 1676037725
transform 1 0 20332 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1676037725
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1676037725
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1676037725
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1676037725
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1676037725
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1676037725
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1676037725
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1676037725
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1676037725
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1676037725
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1676037725
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1676037725
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_617
timestamp 1676037725
transform 1 0 57868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1676037725
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_9
timestamp 1676037725
transform 1 0 1932 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_243
timestamp 1676037725
transform 1 0 23460 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1676037725
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1676037725
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1676037725
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1676037725
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1676037725
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1676037725
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1676037725
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1676037725
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1676037725
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1676037725
transform 1 0 57500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1676037725
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1676037725
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1676037725
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1676037725
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1676037725
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1676037725
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_357
timestamp 1676037725
transform 1 0 33948 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_366
timestamp 1676037725
transform 1 0 34776 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_378
timestamp 1676037725
transform 1 0 35880 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1676037725
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1676037725
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1676037725
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1676037725
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1676037725
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1676037725
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1676037725
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1676037725
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1676037725
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1676037725
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1676037725
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1676037725
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_9
timestamp 1676037725
transform 1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_219
timestamp 1676037725
transform 1 0 21252 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_231
timestamp 1676037725
transform 1 0 22356 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_243
timestamp 1676037725
transform 1 0 23460 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1676037725
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1676037725
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1676037725
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1676037725
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1676037725
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1676037725
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1676037725
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1676037725
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_601
timestamp 1676037725
transform 1 0 56396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_613
timestamp 1676037725
transform 1 0 57500 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1676037725
transform 1 0 58420 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1676037725
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1676037725
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1676037725
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1676037725
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1676037725
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1676037725
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1676037725
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1676037725
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1676037725
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1676037725
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1676037725
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_9
timestamp 1676037725
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1676037725
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1676037725
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1676037725
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1676037725
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1676037725
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1676037725
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1676037725
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1676037725
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1676037725
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1676037725
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1676037725
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1676037725
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1676037725
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_601
timestamp 1676037725
transform 1 0 56396 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1676037725
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1676037725
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1676037725
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1676037725
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1676037725
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1676037725
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1676037725
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1676037725
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1676037725
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1676037725
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1676037725
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1676037725
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1676037725
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1676037725
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_11
timestamp 1676037725
transform 1 0 2116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_23
timestamp 1676037725
transform 1 0 3220 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_269
timestamp 1676037725
transform 1 0 25852 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_281
timestamp 1676037725
transform 1 0 26956 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_293
timestamp 1676037725
transform 1 0 28060 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_305
timestamp 1676037725
transform 1 0 29164 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1676037725
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1676037725
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1676037725
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1676037725
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1676037725
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1676037725
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1676037725
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1676037725
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_601
timestamp 1676037725
transform 1 0 56396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1676037725
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1676037725
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_9
timestamp 1676037725
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1676037725
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_33
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1676037725
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1676037725
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1676037725
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1676037725
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1676037725
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1676037725
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1676037725
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1676037725
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1676037725
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1676037725
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1676037725
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1676037725
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1676037725
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1676037725
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1676037725
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_362
timestamp 1676037725
transform 1 0 34408 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_396
timestamp 1676037725
transform 1 0 37536 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_408
timestamp 1676037725
transform 1 0 38640 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1676037725
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1676037725
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1676037725
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1676037725
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1676037725
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1676037725
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1676037725
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1676037725
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_601
timestamp 1676037725
transform 1 0 56396 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1676037725
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1676037725
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1676037725
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1676037725
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1676037725
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_349
timestamp 1676037725
transform 1 0 33212 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_365
timestamp 1676037725
transform 1 0 34684 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_377
timestamp 1676037725
transform 1 0 35788 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_389
timestamp 1676037725
transform 1 0 36892 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1676037725
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1676037725
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1676037725
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1676037725
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1676037725
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1676037725
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1676037725
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1676037725
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1676037725
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1676037725
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1676037725
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_9
timestamp 1676037725
transform 1 0 1932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1676037725
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1676037725
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1676037725
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_375
timestamp 1676037725
transform 1 0 35604 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_379
timestamp 1676037725
transform 1 0 35972 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_391
timestamp 1676037725
transform 1 0 37076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_403
timestamp 1676037725
transform 1 0 38180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_415
timestamp 1676037725
transform 1 0 39284 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1676037725
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1676037725
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1676037725
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1676037725
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1676037725
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1676037725
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1676037725
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1676037725
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1676037725
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1676037725
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1676037725
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1676037725
transform 1 0 1932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1676037725
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1676037725
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1676037725
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1676037725
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1676037725
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1676037725
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1676037725
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1676037725
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1676037725
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1676037725
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1676037725
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1676037725
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1676037725
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1676037725
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1676037725
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1676037725
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1676037725
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1676037725
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_11
timestamp 1676037725
transform 1 0 2116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1676037725
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1676037725
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1676037725
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1676037725
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1676037725
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_389
timestamp 1676037725
transform 1 0 36892 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_405
timestamp 1676037725
transform 1 0 38364 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1676037725
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1676037725
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1676037725
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1676037725
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1676037725
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1676037725
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1676037725
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1676037725
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1676037725
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_601
timestamp 1676037725
transform 1 0 56396 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1676037725
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1676037725
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_177
timestamp 1676037725
transform 1 0 17388 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_188
timestamp 1676037725
transform 1 0 18400 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_200
timestamp 1676037725
transform 1 0 19504 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_212
timestamp 1676037725
transform 1 0 20608 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1676037725
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_381
timestamp 1676037725
transform 1 0 36156 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1676037725
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1676037725
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1676037725
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1676037725
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1676037725
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1676037725
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1676037725
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1676037725
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1676037725
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1676037725
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1676037725
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1676037725
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1676037725
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1676037725
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1676037725
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1676037725
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1676037725
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1676037725
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1676037725
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1676037725
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1676037725
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1676037725
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1676037725
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1676037725
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1676037725
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1676037725
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_9
timestamp 1676037725
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1676037725
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1676037725
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1676037725
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1676037725
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1676037725
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1676037725
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1676037725
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1676037725
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1676037725
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1676037725
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1676037725
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1676037725
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1676037725
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1676037725
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1676037725
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1676037725
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1676037725
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1676037725
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1676037725
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1676037725
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1676037725
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1676037725
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1676037725
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1676037725
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1676037725
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1676037725
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_623
timestamp 1676037725
transform 1 0 58420 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_9
timestamp 1676037725
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1676037725
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1676037725
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1676037725
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1676037725
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1676037725
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1676037725
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1676037725
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1676037725
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1676037725
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1676037725
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1676037725
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1676037725
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1676037725
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1676037725
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1676037725
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1676037725
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1676037725
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1676037725
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1676037725
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_601
timestamp 1676037725
transform 1 0 56396 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_605
timestamp 1676037725
transform 1 0 56764 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1676037725
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1676037725
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1676037725
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1676037725
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1676037725
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1676037725
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1676037725
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1676037725
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1676037725
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1676037725
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1676037725
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1676037725
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1676037725
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1676037725
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1676037725
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1676037725
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1676037725
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1676037725
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_9
timestamp 1676037725
transform 1 0 1932 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1676037725
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1676037725
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1676037725
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1676037725
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1676037725
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1676037725
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1676037725
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1676037725
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1676037725
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1676037725
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1676037725
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_9
timestamp 1676037725
transform 1 0 1932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1676037725
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1676037725
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1676037725
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1676037725
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1676037725
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1676037725
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1676037725
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1676037725
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1676037725
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1676037725
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1676037725
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1676037725
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1676037725
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1676037725
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1676037725
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_21
timestamp 1676037725
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1676037725
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1676037725
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1676037725
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1676037725
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1676037725
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1676037725
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1676037725
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1676037725
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1676037725
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1676037725
transform 1 0 57500 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1676037725
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_36
timestamp 1676037725
transform 1 0 4416 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_48
timestamp 1676037725
transform 1 0 5520 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1676037725
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1676037725
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1676037725
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1676037725
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1676037725
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1676037725
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1676037725
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1676037725
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1676037725
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1676037725
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1676037725
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1676037725
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1676037725
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1676037725
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1676037725
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1676037725
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1676037725
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1676037725
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1676037725
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1676037725
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1676037725
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1676037725
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_613
timestamp 1676037725
transform 1 0 57500 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_619
timestamp 1676037725
transform 1 0 58052 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1676037725
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_9
timestamp 1676037725
transform 1 0 1932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_66
timestamp 1676037725
transform 1 0 7176 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_78
timestamp 1676037725
transform 1 0 8280 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_90
timestamp 1676037725
transform 1 0 9384 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_102
timestamp 1676037725
transform 1 0 10488 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_110
timestamp 1676037725
transform 1 0 11224 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1676037725
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1676037725
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1676037725
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1676037725
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1676037725
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1676037725
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1676037725
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1676037725
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1676037725
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1676037725
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1676037725
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_11
timestamp 1676037725
transform 1 0 2116 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1676037725
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1676037725
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1676037725
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1676037725
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1676037725
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1676037725
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1676037725
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1676037725
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1676037725
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1676037725
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1676037725
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_9
timestamp 1676037725
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_21
timestamp 1676037725
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_33
timestamp 1676037725
transform 1 0 4140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1676037725
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1676037725
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_247
timestamp 1676037725
transform 1 0 23828 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_260
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_272
timestamp 1676037725
transform 1 0 26128 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1676037725
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1676037725
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1676037725
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1676037725
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1676037725
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1676037725
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1676037725
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1676037725
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1676037725
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1676037725
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1676037725
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_617
timestamp 1676037725
transform 1 0 57868 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1676037725
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1676037725
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1676037725
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1676037725
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1676037725
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1676037725
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1676037725
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1676037725
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1676037725
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1676037725
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1676037725
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1676037725
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_437
timestamp 1676037725
transform 1 0 41308 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_449
timestamp 1676037725
transform 1 0 42412 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_461
timestamp 1676037725
transform 1 0 43516 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_473
timestamp 1676037725
transform 1 0 44620 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1676037725
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1676037725
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1676037725
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1676037725
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1676037725
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1676037725
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1676037725
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1676037725
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1676037725
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1676037725
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1676037725
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_21
timestamp 1676037725
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_33
timestamp 1676037725
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_45
timestamp 1676037725
transform 1 0 5244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1676037725
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1676037725
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1676037725
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1676037725
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1676037725
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1676037725
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1676037725
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1676037725
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1676037725
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1676037725
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1676037725
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1676037725
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1676037725
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1676037725
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1676037725
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1676037725
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1676037725
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1676037725
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1676037725
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1676037725
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1676037725
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1676037725
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1676037725
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1676037725
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1676037725
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1676037725
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1676037725
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1676037725
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1676037725
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1676037725
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1676037725
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1676037725
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1676037725
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1676037725
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1676037725
transform 1 0 1380 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_9
timestamp 1676037725
transform 1 0 1932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_21
timestamp 1676037725
transform 1 0 3036 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1676037725
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1676037725
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1676037725
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1676037725
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1676037725
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1676037725
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1676037725
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1676037725
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1676037725
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1676037725
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1676037725
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1676037725
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1676037725
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1676037725
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1676037725
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1676037725
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1676037725
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1676037725
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1676037725
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1676037725
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1676037725
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1676037725
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_233
timestamp 1676037725
transform 1 0 22540 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_250
timestamp 1676037725
transform 1 0 24104 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1676037725
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1676037725
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1676037725
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1676037725
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1676037725
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1676037725
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1676037725
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1676037725
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1676037725
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1676037725
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1676037725
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1676037725
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1676037725
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1676037725
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1676037725
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1676037725
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1676037725
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1676037725
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1676037725
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1676037725
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1676037725
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1676037725
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1676037725
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1676037725
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1676037725
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1676037725
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1676037725
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1676037725
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1676037725
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1676037725
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1676037725
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1676037725
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1676037725
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1676037725
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1676037725
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1676037725
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1676037725
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1676037725
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_613
timestamp 1676037725
transform 1 0 57500 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_619
timestamp 1676037725
transform 1 0 58052 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1676037725
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1676037725
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_9
timestamp 1676037725
transform 1 0 1932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_21
timestamp 1676037725
transform 1 0 3036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_33
timestamp 1676037725
transform 1 0 4140 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_45
timestamp 1676037725
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1676037725
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1676037725
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1676037725
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1676037725
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1676037725
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1676037725
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1676037725
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1676037725
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1676037725
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1676037725
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1676037725
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1676037725
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1676037725
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1676037725
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1676037725
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1676037725
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1676037725
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1676037725
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1676037725
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1676037725
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1676037725
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1676037725
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1676037725
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1676037725
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1676037725
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1676037725
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1676037725
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1676037725
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1676037725
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1676037725
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1676037725
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1676037725
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1676037725
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1676037725
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1676037725
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1676037725
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1676037725
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1676037725
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1676037725
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_417
timestamp 1676037725
transform 1 0 39468 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_421
timestamp 1676037725
transform 1 0 39836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_436
timestamp 1676037725
transform 1 0 41216 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1676037725
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1676037725
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1676037725
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1676037725
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1676037725
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1676037725
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1676037725
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1676037725
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1676037725
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1676037725
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1676037725
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1676037725
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1676037725
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1676037725
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1676037725
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1676037725
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1676037725
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1676037725
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1676037725
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1676037725
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_9
timestamp 1676037725
transform 1 0 1932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_21
timestamp 1676037725
transform 1 0 3036 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1676037725
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1676037725
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1676037725
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1676037725
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1676037725
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1676037725
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1676037725
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1676037725
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1676037725
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1676037725
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1676037725
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1676037725
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1676037725
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1676037725
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1676037725
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1676037725
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1676037725
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1676037725
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1676037725
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1676037725
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1676037725
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1676037725
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1676037725
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1676037725
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1676037725
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1676037725
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1676037725
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_291
timestamp 1676037725
transform 1 0 27876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_303
timestamp 1676037725
transform 1 0 28980 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1676037725
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1676037725
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1676037725
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1676037725
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1676037725
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1676037725
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1676037725
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1676037725
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1676037725
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1676037725
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1676037725
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1676037725
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1676037725
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1676037725
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1676037725
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1676037725
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1676037725
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1676037725
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1676037725
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1676037725
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1676037725
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1676037725
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1676037725
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1676037725
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1676037725
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1676037725
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1676037725
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1676037725
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1676037725
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1676037725
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1676037725
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1676037725
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1676037725
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_613
timestamp 1676037725
transform 1 0 57500 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_619
timestamp 1676037725
transform 1 0 58052 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1676037725
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1676037725
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1676037725
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1676037725
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1676037725
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1676037725
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1676037725
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1676037725
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1676037725
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1676037725
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1676037725
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1676037725
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1676037725
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1676037725
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1676037725
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1676037725
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1676037725
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1676037725
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1676037725
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1676037725
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1676037725
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1676037725
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1676037725
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1676037725
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1676037725
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1676037725
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1676037725
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1676037725
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1676037725
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1676037725
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1676037725
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1676037725
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_293
timestamp 1676037725
transform 1 0 28060 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_313
timestamp 1676037725
transform 1 0 29900 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_325
timestamp 1676037725
transform 1 0 31004 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_333
timestamp 1676037725
transform 1 0 31740 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1676037725
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1676037725
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1676037725
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_373
timestamp 1676037725
transform 1 0 35420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_387
timestamp 1676037725
transform 1 0 36708 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1676037725
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1676037725
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1676037725
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_417
timestamp 1676037725
transform 1 0 39468 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_425
timestamp 1676037725
transform 1 0 40204 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_442
timestamp 1676037725
transform 1 0 41768 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1676037725
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1676037725
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1676037725
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1676037725
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1676037725
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1676037725
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1676037725
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1676037725
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1676037725
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1676037725
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1676037725
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1676037725
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1676037725
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1676037725
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1676037725
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1676037725
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1676037725
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1676037725
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_617
timestamp 1676037725
transform 1 0 57868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1676037725
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1676037725
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_9
timestamp 1676037725
transform 1 0 1932 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_21
timestamp 1676037725
transform 1 0 3036 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1676037725
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1676037725
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1676037725
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1676037725
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1676037725
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1676037725
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1676037725
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1676037725
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1676037725
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1676037725
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1676037725
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1676037725
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1676037725
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1676037725
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1676037725
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1676037725
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1676037725
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1676037725
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1676037725
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1676037725
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1676037725
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1676037725
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1676037725
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1676037725
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1676037725
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1676037725
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1676037725
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1676037725
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1676037725
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1676037725
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1676037725
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1676037725
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1676037725
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1676037725
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_345
timestamp 1676037725
transform 1 0 32844 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_361
timestamp 1676037725
transform 1 0 34316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_365
timestamp 1676037725
transform 1 0 34684 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_369
timestamp 1676037725
transform 1 0 35052 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_387
timestamp 1676037725
transform 1 0 36708 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_399
timestamp 1676037725
transform 1 0 37812 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_411
timestamp 1676037725
transform 1 0 38916 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1676037725
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1676037725
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1676037725
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1676037725
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1676037725
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1676037725
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1676037725
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1676037725
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1676037725
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1676037725
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1676037725
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1676037725
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1676037725
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1676037725
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1676037725
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1676037725
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1676037725
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1676037725
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1676037725
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1676037725
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1676037725
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_613
timestamp 1676037725
transform 1 0 57500 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1676037725
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1676037725
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_9
timestamp 1676037725
transform 1 0 1932 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_21
timestamp 1676037725
transform 1 0 3036 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_33
timestamp 1676037725
transform 1 0 4140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1676037725
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1676037725
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1676037725
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1676037725
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1676037725
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1676037725
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1676037725
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1676037725
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1676037725
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1676037725
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1676037725
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1676037725
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1676037725
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1676037725
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1676037725
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1676037725
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1676037725
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1676037725
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1676037725
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1676037725
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1676037725
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1676037725
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1676037725
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1676037725
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1676037725
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1676037725
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1676037725
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1676037725
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1676037725
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1676037725
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1676037725
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1676037725
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1676037725
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1676037725
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1676037725
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_373
timestamp 1676037725
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1676037725
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1676037725
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1676037725
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1676037725
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1676037725
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1676037725
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1676037725
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1676037725
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1676037725
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1676037725
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1676037725
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1676037725
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1676037725
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1676037725
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1676037725
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1676037725
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1676037725
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1676037725
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1676037725
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1676037725
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1676037725
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1676037725
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1676037725
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1676037725
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1676037725
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1676037725
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1676037725
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_3
timestamp 1676037725
transform 1 0 1380 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_11
timestamp 1676037725
transform 1 0 2116 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_23
timestamp 1676037725
transform 1 0 3220 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1676037725
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1676037725
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1676037725
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1676037725
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1676037725
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1676037725
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1676037725
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1676037725
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1676037725
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1676037725
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1676037725
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1676037725
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1676037725
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1676037725
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1676037725
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1676037725
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1676037725
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1676037725
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1676037725
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1676037725
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1676037725
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1676037725
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1676037725
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1676037725
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1676037725
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1676037725
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1676037725
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1676037725
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1676037725
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1676037725
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1676037725
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1676037725
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1676037725
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1676037725
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1676037725
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1676037725
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1676037725
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_365
timestamp 1676037725
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_377
timestamp 1676037725
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_389
timestamp 1676037725
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_401
timestamp 1676037725
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_413
timestamp 1676037725
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1676037725
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1676037725
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1676037725
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1676037725
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1676037725
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1676037725
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1676037725
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1676037725
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1676037725
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1676037725
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1676037725
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1676037725
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1676037725
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1676037725
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1676037725
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1676037725
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1676037725
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1676037725
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1676037725
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1676037725
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1676037725
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_613
timestamp 1676037725
transform 1 0 57500 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_623
timestamp 1676037725
transform 1 0 58420 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_3
timestamp 1676037725
transform 1 0 1380 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_11
timestamp 1676037725
transform 1 0 2116 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_23
timestamp 1676037725
transform 1 0 3220 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_35
timestamp 1676037725
transform 1 0 4324 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_47
timestamp 1676037725
transform 1 0 5428 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1676037725
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1676037725
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1676037725
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1676037725
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1676037725
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1676037725
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1676037725
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1676037725
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1676037725
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1676037725
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1676037725
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1676037725
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1676037725
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1676037725
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1676037725
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1676037725
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1676037725
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1676037725
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1676037725
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1676037725
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1676037725
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1676037725
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1676037725
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1676037725
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1676037725
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1676037725
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1676037725
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1676037725
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1676037725
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1676037725
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1676037725
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1676037725
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1676037725
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1676037725
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1676037725
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1676037725
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1676037725
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_393
timestamp 1676037725
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_405
timestamp 1676037725
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_417
timestamp 1676037725
transform 1 0 39468 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_423
timestamp 1676037725
transform 1 0 40020 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_438
timestamp 1676037725
transform 1 0 41400 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_446
timestamp 1676037725
transform 1 0 42136 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1676037725
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1676037725
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1676037725
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1676037725
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1676037725
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1676037725
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1676037725
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1676037725
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1676037725
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1676037725
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1676037725
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1676037725
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1676037725
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1676037725
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1676037725
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1676037725
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1676037725
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1676037725
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_617
timestamp 1676037725
transform 1 0 57868 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_623
timestamp 1676037725
transform 1 0 58420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_3
timestamp 1676037725
transform 1 0 1380 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_9
timestamp 1676037725
transform 1 0 1932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_21
timestamp 1676037725
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1676037725
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1676037725
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1676037725
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1676037725
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1676037725
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1676037725
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1676037725
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1676037725
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1676037725
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1676037725
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1676037725
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1676037725
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1676037725
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1676037725
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1676037725
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1676037725
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1676037725
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1676037725
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1676037725
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_197
timestamp 1676037725
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_209
timestamp 1676037725
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_221
timestamp 1676037725
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_233
timestamp 1676037725
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1676037725
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1676037725
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1676037725
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1676037725
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1676037725
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1676037725
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1676037725
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1676037725
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1676037725
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1676037725
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1676037725
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1676037725
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1676037725
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1676037725
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1676037725
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_377
timestamp 1676037725
transform 1 0 35788 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_385
timestamp 1676037725
transform 1 0 36524 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_404
timestamp 1676037725
transform 1 0 38272 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_416
timestamp 1676037725
transform 1 0 39376 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_104_421
timestamp 1676037725
transform 1 0 39836 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_438
timestamp 1676037725
transform 1 0 41400 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_450
timestamp 1676037725
transform 1 0 42504 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_462
timestamp 1676037725
transform 1 0 43608 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_104_474
timestamp 1676037725
transform 1 0 44712 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1676037725
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1676037725
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1676037725
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1676037725
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1676037725
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1676037725
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1676037725
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1676037725
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1676037725
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1676037725
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1676037725
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1676037725
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1676037725
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_601
timestamp 1676037725
transform 1 0 56396 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_613
timestamp 1676037725
transform 1 0 57500 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_623
timestamp 1676037725
transform 1 0 58420 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_3
timestamp 1676037725
transform 1 0 1380 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_9
timestamp 1676037725
transform 1 0 1932 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_17
timestamp 1676037725
transform 1 0 2668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_29
timestamp 1676037725
transform 1 0 3772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_41
timestamp 1676037725
transform 1 0 4876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_53
timestamp 1676037725
transform 1 0 5980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_57
timestamp 1676037725
transform 1 0 6348 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_66
timestamp 1676037725
transform 1 0 7176 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_78
timestamp 1676037725
transform 1 0 8280 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_90
timestamp 1676037725
transform 1 0 9384 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_102
timestamp 1676037725
transform 1 0 10488 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_110
timestamp 1676037725
transform 1 0 11224 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1676037725
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1676037725
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1676037725
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1676037725
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1676037725
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1676037725
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1676037725
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_181
timestamp 1676037725
transform 1 0 17756 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_187
timestamp 1676037725
transform 1 0 18308 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_190
timestamp 1676037725
transform 1 0 18584 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_200
timestamp 1676037725
transform 1 0 19504 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_212
timestamp 1676037725
transform 1 0 20608 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_225
timestamp 1676037725
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_237
timestamp 1676037725
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_249
timestamp 1676037725
transform 1 0 24012 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_105_259
timestamp 1676037725
transform 1 0 24932 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_265
timestamp 1676037725
transform 1 0 25484 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_105_274
timestamp 1676037725
transform 1 0 26312 0 -1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1676037725
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_293
timestamp 1676037725
transform 1 0 28060 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_301
timestamp 1676037725
transform 1 0 28796 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_304
timestamp 1676037725
transform 1 0 29072 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_316
timestamp 1676037725
transform 1 0 30176 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_328
timestamp 1676037725
transform 1 0 31280 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1676037725
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1676037725
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1676037725
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1676037725
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1676037725
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1676037725
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1676037725
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1676037725
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1676037725
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1676037725
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1676037725
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1676037725
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_449
timestamp 1676037725
transform 1 0 42412 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_465
timestamp 1676037725
transform 1 0 43884 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_477
timestamp 1676037725
transform 1 0 44988 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_489
timestamp 1676037725
transform 1 0 46092 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_501
timestamp 1676037725
transform 1 0 47196 0 -1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1676037725
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1676037725
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1676037725
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1676037725
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1676037725
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1676037725
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1676037725
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1676037725
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1676037725
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1676037725
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_609
timestamp 1676037725
transform 1 0 57132 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_614
timestamp 1676037725
transform 1 0 57592 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_617
timestamp 1676037725
transform 1 0 57868 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_623
timestamp 1676037725
transform 1 0 58420 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_3
timestamp 1676037725
transform 1 0 1380 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_11
timestamp 1676037725
transform 1 0 2116 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1676037725
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1676037725
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1676037725
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1676037725
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_61
timestamp 1676037725
transform 1 0 6716 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_73
timestamp 1676037725
transform 1 0 7820 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_81
timestamp 1676037725
transform 1 0 8556 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1676037725
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1676037725
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1676037725
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1676037725
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1676037725
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1676037725
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1676037725
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1676037725
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1676037725
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_177
timestamp 1676037725
transform 1 0 17388 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_106_193
timestamp 1676037725
transform 1 0 18860 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_197
timestamp 1676037725
transform 1 0 19228 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_213
timestamp 1676037725
transform 1 0 20700 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_226
timestamp 1676037725
transform 1 0 21896 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_238
timestamp 1676037725
transform 1 0 23000 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_250
timestamp 1676037725
transform 1 0 24104 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_106_253
timestamp 1676037725
transform 1 0 24380 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_106_273
timestamp 1676037725
transform 1 0 26220 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_277
timestamp 1676037725
transform 1 0 26588 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_288
timestamp 1676037725
transform 1 0 27600 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_300
timestamp 1676037725
transform 1 0 28704 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_306
timestamp 1676037725
transform 1 0 29256 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_309
timestamp 1676037725
transform 1 0 29532 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_319
timestamp 1676037725
transform 1 0 30452 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_323
timestamp 1676037725
transform 1 0 30820 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_335
timestamp 1676037725
transform 1 0 31924 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_343
timestamp 1676037725
transform 1 0 32660 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_346
timestamp 1676037725
transform 1 0 32936 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_362
timestamp 1676037725
transform 1 0 34408 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_365
timestamp 1676037725
transform 1 0 34684 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_369
timestamp 1676037725
transform 1 0 35052 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_381
timestamp 1676037725
transform 1 0 36156 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_393
timestamp 1676037725
transform 1 0 37260 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_405
timestamp 1676037725
transform 1 0 38364 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_417
timestamp 1676037725
transform 1 0 39468 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1676037725
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_447
timestamp 1676037725
transform 1 0 42228 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_465
timestamp 1676037725
transform 1 0 43884 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_473
timestamp 1676037725
transform 1 0 44620 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1676037725
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1676037725
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1676037725
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1676037725
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1676037725
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1676037725
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1676037725
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1676037725
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1676037725
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1676037725
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1676037725
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1676037725
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1676037725
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_605
timestamp 1676037725
transform 1 0 56764 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_613
timestamp 1676037725
transform 1 0 57500 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_623
timestamp 1676037725
transform 1 0 58420 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_3
timestamp 1676037725
transform 1 0 1380 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_107_11
timestamp 1676037725
transform 1 0 2116 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_19
timestamp 1676037725
transform 1 0 2852 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_26
timestamp 1676037725
transform 1 0 3496 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_34
timestamp 1676037725
transform 1 0 4232 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_50
timestamp 1676037725
transform 1 0 5704 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1676037725
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_69
timestamp 1676037725
transform 1 0 7452 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_77
timestamp 1676037725
transform 1 0 8188 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_82
timestamp 1676037725
transform 1 0 8648 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_98
timestamp 1676037725
transform 1 0 10120 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_110
timestamp 1676037725
transform 1 0 11224 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1676037725
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_125
timestamp 1676037725
transform 1 0 12604 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_133
timestamp 1676037725
transform 1 0 13340 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_138
timestamp 1676037725
transform 1 0 13800 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_146
timestamp 1676037725
transform 1 0 14536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_162
timestamp 1676037725
transform 1 0 16008 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1676037725
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1676037725
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_193
timestamp 1676037725
transform 1 0 18860 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_197
timestamp 1676037725
transform 1 0 19228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_202
timestamp 1676037725
transform 1 0 19688 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_214
timestamp 1676037725
transform 1 0 20792 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_222
timestamp 1676037725
transform 1 0 21528 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_225
timestamp 1676037725
transform 1 0 21804 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_236
timestamp 1676037725
transform 1 0 22816 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_244
timestamp 1676037725
transform 1 0 23552 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_252
timestamp 1676037725
transform 1 0 24288 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_258
timestamp 1676037725
transform 1 0 24840 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_270
timestamp 1676037725
transform 1 0 25944 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_278
timestamp 1676037725
transform 1 0 26680 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_281
timestamp 1676037725
transform 1 0 26956 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_285
timestamp 1676037725
transform 1 0 27324 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_290
timestamp 1676037725
transform 1 0 27784 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_306
timestamp 1676037725
transform 1 0 29256 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_322
timestamp 1676037725
transform 1 0 30728 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_334
timestamp 1676037725
transform 1 0 31832 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1676037725
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1676037725
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1676037725
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_373
timestamp 1676037725
transform 1 0 35420 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_381
timestamp 1676037725
transform 1 0 36156 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_386
timestamp 1676037725
transform 1 0 36616 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1676037725
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1676037725
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1676037725
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_429
timestamp 1676037725
transform 1 0 40572 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_437
timestamp 1676037725
transform 1 0 41308 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_442
timestamp 1676037725
transform 1 0 41768 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1676037725
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1676037725
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1676037725
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_485
timestamp 1676037725
transform 1 0 45724 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_493
timestamp 1676037725
transform 1 0 46460 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_498
timestamp 1676037725
transform 1 0 46920 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1676037725
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1676037725
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_529
timestamp 1676037725
transform 1 0 49772 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_533
timestamp 1676037725
transform 1 0 50140 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_538
timestamp 1676037725
transform 1 0 50600 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_550
timestamp 1676037725
transform 1 0 51704 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_558
timestamp 1676037725
transform 1 0 52440 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_561
timestamp 1676037725
transform 1 0 52716 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_567
timestamp 1676037725
transform 1 0 53268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_579
timestamp 1676037725
transform 1 0 54372 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_586
timestamp 1676037725
transform 1 0 55016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_594
timestamp 1676037725
transform 1 0 55752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_602
timestamp 1676037725
transform 1 0 56488 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_107_610
timestamp 1676037725
transform 1 0 57224 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_107_617
timestamp 1676037725
transform 1 0 57868 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_623
timestamp 1676037725
transform 1 0 58420 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_3
timestamp 1676037725
transform 1 0 1380 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_14
timestamp 1676037725
transform 1 0 2392 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_24
timestamp 1676037725
transform 1 0 3312 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_29
timestamp 1676037725
transform 1 0 3772 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_37
timestamp 1676037725
transform 1 0 4508 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_42
timestamp 1676037725
transform 1 0 4968 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_108_54
timestamp 1676037725
transform 1 0 6072 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_57
timestamp 1676037725
transform 1 0 6348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_66
timestamp 1676037725
transform 1 0 7176 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_76
timestamp 1676037725
transform 1 0 8096 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_85
timestamp 1676037725
transform 1 0 8924 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_93
timestamp 1676037725
transform 1 0 9660 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_97
timestamp 1676037725
transform 1 0 10028 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_102
timestamp 1676037725
transform 1 0 10488 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_110
timestamp 1676037725
transform 1 0 11224 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_113
timestamp 1676037725
transform 1 0 11500 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_117
timestamp 1676037725
transform 1 0 11868 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_122
timestamp 1676037725
transform 1 0 12328 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_132
timestamp 1676037725
transform 1 0 13248 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_141
timestamp 1676037725
transform 1 0 14076 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_149
timestamp 1676037725
transform 1 0 14812 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_156
timestamp 1676037725
transform 1 0 15456 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_108_166
timestamp 1676037725
transform 1 0 16376 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_169
timestamp 1676037725
transform 1 0 16652 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_173
timestamp 1676037725
transform 1 0 17020 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_178
timestamp 1676037725
transform 1 0 17480 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_186
timestamp 1676037725
transform 1 0 18216 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_194
timestamp 1676037725
transform 1 0 18952 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_197
timestamp 1676037725
transform 1 0 19228 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_201
timestamp 1676037725
transform 1 0 19596 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_206
timestamp 1676037725
transform 1 0 20056 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_214
timestamp 1676037725
transform 1 0 20792 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_222
timestamp 1676037725
transform 1 0 21528 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_225
timestamp 1676037725
transform 1 0 21804 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_229
timestamp 1676037725
transform 1 0 22172 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_236
timestamp 1676037725
transform 1 0 22816 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_244
timestamp 1676037725
transform 1 0 23552 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_250
timestamp 1676037725
transform 1 0 24104 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_253
timestamp 1676037725
transform 1 0 24380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_261
timestamp 1676037725
transform 1 0 25116 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_268
timestamp 1676037725
transform 1 0 25760 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_276
timestamp 1676037725
transform 1 0 26496 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_281
timestamp 1676037725
transform 1 0 26956 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_289
timestamp 1676037725
transform 1 0 27692 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_293
timestamp 1676037725
transform 1 0 28060 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_300
timestamp 1676037725
transform 1 0 28704 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_309
timestamp 1676037725
transform 1 0 29532 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_317
timestamp 1676037725
transform 1 0 30268 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_325
timestamp 1676037725
transform 1 0 31004 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_332
timestamp 1676037725
transform 1 0 31648 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_337
timestamp 1676037725
transform 1 0 32108 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_345
timestamp 1676037725
transform 1 0 32844 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_353
timestamp 1676037725
transform 1 0 33580 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_361
timestamp 1676037725
transform 1 0 34316 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_365
timestamp 1676037725
transform 1 0 34684 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_371
timestamp 1676037725
transform 1 0 35236 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_379
timestamp 1676037725
transform 1 0 35972 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_387
timestamp 1676037725
transform 1 0 36708 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_391
timestamp 1676037725
transform 1 0 37076 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_393
timestamp 1676037725
transform 1 0 37260 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_399
timestamp 1676037725
transform 1 0 37812 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_407
timestamp 1676037725
transform 1 0 38548 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_415
timestamp 1676037725
transform 1 0 39284 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1676037725
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_421
timestamp 1676037725
transform 1 0 39836 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_427
timestamp 1676037725
transform 1 0 40388 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_435
timestamp 1676037725
transform 1 0 41124 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_443
timestamp 1676037725
transform 1 0 41860 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_447
timestamp 1676037725
transform 1 0 42228 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_449
timestamp 1676037725
transform 1 0 42412 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_457
timestamp 1676037725
transform 1 0 43148 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_465
timestamp 1676037725
transform 1 0 43884 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_473
timestamp 1676037725
transform 1 0 44620 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_477
timestamp 1676037725
transform 1 0 44988 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_483
timestamp 1676037725
transform 1 0 45540 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_491
timestamp 1676037725
transform 1 0 46276 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_499
timestamp 1676037725
transform 1 0 47012 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_503
timestamp 1676037725
transform 1 0 47380 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_505
timestamp 1676037725
transform 1 0 47564 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_511
timestamp 1676037725
transform 1 0 48116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_519
timestamp 1676037725
transform 1 0 48852 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_527
timestamp 1676037725
transform 1 0 49588 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1676037725
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_533
timestamp 1676037725
transform 1 0 50140 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_541
timestamp 1676037725
transform 1 0 50876 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_549
timestamp 1676037725
transform 1 0 51612 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_557
timestamp 1676037725
transform 1 0 52348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_561
timestamp 1676037725
transform 1 0 52716 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_565
timestamp 1676037725
transform 1 0 53084 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_572
timestamp 1676037725
transform 1 0 53728 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_580
timestamp 1676037725
transform 1 0 54464 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_589
timestamp 1676037725
transform 1 0 55292 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_597
timestamp 1676037725
transform 1 0 56028 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_607
timestamp 1676037725
transform 1 0 56948 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_615
timestamp 1676037725
transform 1 0 57684 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_617
timestamp 1676037725
transform 1 0 57868 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_623
timestamp 1676037725
transform 1 0 58420 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1676037725
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1676037725
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1676037725
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1676037725
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1676037725
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1676037725
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1676037725
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1676037725
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1676037725
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1676037725
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1676037725
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1676037725
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1676037725
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1676037725
transform -1 0 58880 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1676037725
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1676037725
transform -1 0 58880 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1676037725
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1676037725
transform -1 0 58880 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1676037725
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1676037725
transform -1 0 58880 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1676037725
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1676037725
transform -1 0 58880 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1676037725
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1676037725
transform -1 0 58880 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1676037725
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1676037725
transform -1 0 58880 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 6256 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 11408 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 16560 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 21712 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 26864 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 32016 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 37168 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 42320 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 47472 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 52624 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 57776 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1676037725
transform 1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0452_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1676037725
transform 1 0 45172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1676037725
transform 1 0 40020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_4  _0459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_4  _0460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _0461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _0463_
timestamp 1676037725
transform 1 0 19596 0 1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20240 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_4  _0468_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0469_
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0470_
timestamp 1676037725
transform 1 0 22724 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0471_
timestamp 1676037725
transform 1 0 17848 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0472_
timestamp 1676037725
transform 1 0 20884 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0473_
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _0474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _0475_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0477_
timestamp 1676037725
transform 1 0 19780 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_2  _0478_
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0480_
timestamp 1676037725
transform 1 0 19780 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0481_
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _0482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _0483_
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _0484_
timestamp 1676037725
transform 1 0 19504 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _0485_
timestamp 1676037725
transform 1 0 16928 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _0486_
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0487_
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _0489_
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33028 0 1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0495_
timestamp 1676037725
transform 1 0 33580 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22724 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0498_
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0501_
timestamp 1676037725
transform 1 0 32292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0502_
timestamp 1676037725
transform 1 0 33948 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0503_
timestamp 1676037725
transform 1 0 43516 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0504_
timestamp 1676037725
transform 1 0 33120 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0505_
timestamp 1676037725
transform 1 0 33672 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0506_
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33488 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0508_
timestamp 1676037725
transform 1 0 34408 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0509_
timestamp 1676037725
transform 1 0 38548 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0510_
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0512_
timestamp 1676037725
transform 1 0 52624 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0513_
timestamp 1676037725
transform 1 0 34868 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0514_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0515_
timestamp 1676037725
transform 1 0 35972 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38916 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0517_
timestamp 1676037725
transform 1 0 35972 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0518_
timestamp 1676037725
transform 1 0 17572 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0519_
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0520_
timestamp 1676037725
transform 1 0 36248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0521_
timestamp 1676037725
transform 1 0 35512 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _0522_
timestamp 1676037725
transform 1 0 36156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0523_
timestamp 1676037725
transform 1 0 37628 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0524_
timestamp 1676037725
transform 1 0 34040 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0525_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0526_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0527_
timestamp 1676037725
transform 1 0 35144 0 1 56576
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _0528_
timestamp 1676037725
transform 1 0 19596 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0530_
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0531_
timestamp 1676037725
transform 1 0 24656 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _0532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0533_
timestamp 1676037725
transform 1 0 36248 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0534_
timestamp 1676037725
transform 1 0 36708 0 1 58752
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0535_
timestamp 1676037725
transform 1 0 25576 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0536_
timestamp 1676037725
transform 1 0 25944 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0537_
timestamp 1676037725
transform 1 0 25300 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0538_
timestamp 1676037725
transform 1 0 26680 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0539_
timestamp 1676037725
transform 1 0 25300 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0540_
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 1676037725
transform 1 0 24288 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0542_
timestamp 1676037725
transform 1 0 24656 0 1 59840
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0543_
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25576 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1676037725
transform 1 0 25576 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0546_
timestamp 1676037725
transform 1 0 18768 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0547_
timestamp 1676037725
transform 1 0 19228 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0548_
timestamp 1676037725
transform 1 0 53452 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20516 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0550_
timestamp 1676037725
transform 1 0 18308 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0551_
timestamp 1676037725
transform 1 0 18768 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0553_
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0554_
timestamp 1676037725
transform 1 0 19504 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0556_
timestamp 1676037725
transform 1 0 53636 0 -1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0557_
timestamp 1676037725
transform 1 0 2024 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0560_
timestamp 1676037725
transform 1 0 5980 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0562_
timestamp 1676037725
transform 1 0 20608 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_4  _0563_
timestamp 1676037725
transform 1 0 19136 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0564_
timestamp 1676037725
transform 1 0 19964 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 1676037725
transform 1 0 19504 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0566_
timestamp 1676037725
transform 1 0 20792 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 1676037725
transform 1 0 40020 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0568_
timestamp 1676037725
transform 1 0 2300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0569_
timestamp 1676037725
transform 1 0 21804 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0573_
timestamp 1676037725
transform 1 0 22264 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0574_
timestamp 1676037725
transform 1 0 22724 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0575_
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0576_
timestamp 1676037725
transform 1 0 22448 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0577_
timestamp 1676037725
transform 1 0 40296 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1676037725
transform 1 0 23828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23460 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0581_
timestamp 1676037725
transform 1 0 20608 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0582_
timestamp 1676037725
transform 1 0 40020 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp 1676037725
transform 1 0 2024 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0584_
timestamp 1676037725
transform 1 0 40940 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a2111o_1  _0585_
timestamp 1676037725
transform 1 0 20056 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0586_
timestamp 1676037725
transform 1 0 21068 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1676037725
transform 1 0 27232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0589_
timestamp 1676037725
transform 1 0 33396 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0590_
timestamp 1676037725
transform 1 0 3680 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0591_
timestamp 1676037725
transform 1 0 5060 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0593_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0594_
timestamp 1676037725
transform 1 0 17940 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1676037725
transform 1 0 35604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp 1676037725
transform 1 0 23368 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0598_
timestamp 1676037725
transform 1 0 22080 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0599_
timestamp 1676037725
transform 1 0 6532 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0600_
timestamp 1676037725
transform 1 0 6532 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0601_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0602_
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_4  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0604_
timestamp 1676037725
transform 1 0 23368 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0605_
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 1676037725
transform 1 0 31096 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0610_
timestamp 1676037725
transform 1 0 23092 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0611_
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1676037725
transform 1 0 23460 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0613_
timestamp 1676037725
transform 1 0 24288 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0614_
timestamp 1676037725
transform 1 0 40020 0 1 53312
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp 1676037725
transform 1 0 40664 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0616_
timestamp 1676037725
transform 1 0 39928 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0617_
timestamp 1676037725
transform 1 0 39652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0618_
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0619_
timestamp 1676037725
transform 1 0 41676 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0620_
timestamp 1676037725
transform 1 0 26772 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0621_
timestamp 1676037725
transform 1 0 22816 0 1 54400
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0622_
timestamp 1676037725
transform 1 0 40020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0623_
timestamp 1676037725
transform 1 0 39928 0 -1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_1  _0624_
timestamp 1676037725
transform 1 0 41032 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0625_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0626_
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0627_
timestamp 1676037725
transform 1 0 27968 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0628_
timestamp 1676037725
transform 1 0 26588 0 1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0629_
timestamp 1676037725
transform 1 0 40480 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp 1676037725
transform 1 0 40296 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0631_
timestamp 1676037725
transform 1 0 40756 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0632_
timestamp 1676037725
transform 1 0 42596 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1676037725
transform 1 0 29716 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0634_
timestamp 1676037725
transform 1 0 28612 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _0635_
timestamp 1676037725
transform 1 0 33580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0637_
timestamp 1676037725
transform 1 0 41308 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0638_
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0639_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0640_
timestamp 1676037725
transform 1 0 42596 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0641_
timestamp 1676037725
transform 1 0 42320 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0642_
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0643_
timestamp 1676037725
transform 1 0 40112 0 1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0644_
timestamp 1676037725
transform 1 0 40020 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0645_
timestamp 1676037725
transform 1 0 41124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0646_
timestamp 1676037725
transform 1 0 40112 0 -1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0647_
timestamp 1676037725
transform 1 0 39652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0648_
timestamp 1676037725
transform 1 0 40296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0649_
timestamp 1676037725
transform 1 0 42596 0 -1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0650_
timestamp 1676037725
transform 1 0 43332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0651_
timestamp 1676037725
transform 1 0 32292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0652_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _0653_
timestamp 1676037725
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0655_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0658_
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0659_
timestamp 1676037725
transform 1 0 28612 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0660_
timestamp 1676037725
transform 1 0 9384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0661_
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1676037725
transform 1 0 17572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0663_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0664_
timestamp 1676037725
transform 1 0 7728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0665_
timestamp 1676037725
transform 1 0 8648 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0667_
timestamp 1676037725
transform 1 0 9200 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1676037725
transform 1 0 7912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 1676037725
transform 1 0 9568 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1676037725
transform 1 0 10212 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0671_
timestamp 1676037725
transform 1 0 9660 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0672_
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0673_
timestamp 1676037725
transform 1 0 10120 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0674_
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0675_
timestamp 1676037725
transform 1 0 10120 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0676_
timestamp 1676037725
transform 1 0 18492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0677_
timestamp 1676037725
transform 1 0 15916 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0678_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11224 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0679_
timestamp 1676037725
transform 1 0 31188 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0680_
timestamp 1676037725
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0681_
timestamp 1676037725
transform 1 0 30176 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0682_
timestamp 1676037725
transform 1 0 15824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0683_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0684_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0685_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1676037725
transform 1 0 11316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0687_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0688_
timestamp 1676037725
transform 1 0 10304 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0689_
timestamp 1676037725
transform 1 0 21620 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0690_
timestamp 1676037725
transform 1 0 12328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0691_
timestamp 1676037725
transform 1 0 23000 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0692_
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0693_
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0694_
timestamp 1676037725
transform 1 0 11316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0695_
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0696_
timestamp 1676037725
transform 1 0 13156 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0697_
timestamp 1676037725
transform 1 0 20424 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0698_
timestamp 1676037725
transform 1 0 10672 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0699_
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0700_
timestamp 1676037725
transform 1 0 12144 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0701_
timestamp 1676037725
transform 1 0 19412 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0702_
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0703_
timestamp 1676037725
transform 1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0704_
timestamp 1676037725
transform 1 0 14720 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0705_
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0706_
timestamp 1676037725
transform 1 0 14720 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0707_
timestamp 1676037725
transform 1 0 20608 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0708_
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0709_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0710_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0711_
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 57040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42412 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1676037725
transform 1 0 35972 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0716_
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1676037725
transform 1 0 28336 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1676037725
transform 1 0 30820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1676037725
transform 1 0 34960 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0720_
timestamp 1676037725
transform 1 0 36800 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1676037725
transform 1 0 37720 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1676037725
transform 1 0 37904 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1676037725
transform 1 0 30268 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1676037725
transform 1 0 35972 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1676037725
transform 1 0 29900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1676037725
transform 1 0 28980 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0730_
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1676037725
transform 1 0 36156 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0733_
timestamp 1676037725
transform 1 0 38548 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0735_
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1676037725
transform 1 0 33120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0737_
timestamp 1676037725
transform 1 0 37076 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1676037725
transform 1 0 34040 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0739_
timestamp 1676037725
transform 1 0 38732 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0741_
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1676037725
transform 1 0 30820 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0743_
timestamp 1676037725
transform 1 0 36156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1676037725
transform 1 0 27416 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1676037725
transform 1 0 36984 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1676037725
transform 1 0 30912 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0749_
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0751_
timestamp 1676037725
transform 1 0 28336 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1676037725
transform 1 0 28060 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0753_
timestamp 1676037725
transform 1 0 26404 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1676037725
transform 1 0 38088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0755_
timestamp 1676037725
transform 1 0 39376 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp 1676037725
transform 1 0 36432 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1676037725
transform 1 0 30820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1676037725
transform 1 0 40296 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1676037725
transform 1 0 41400 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1676037725
transform 1 0 28428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1676037725
transform 1 0 28980 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1676037725
transform 1 0 38548 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1676037725
transform 1 0 38548 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1676037725
transform 1 0 40480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1676037725
transform 1 0 40480 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1676037725
transform 1 0 35052 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0775_
timestamp 1676037725
transform 1 0 36248 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1676037725
transform 1 0 33028 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0779_
timestamp 1676037725
transform 1 0 34868 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1676037725
transform 1 0 48208 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_4  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42872 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1676037725
transform 1 0 35236 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1676037725
transform 1 0 29900 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1676037725
transform 1 0 29808 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1676037725
transform 1 0 27692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1676037725
transform 1 0 27968 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1676037725
transform 1 0 25852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1676037725
transform 1 0 37536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1676037725
transform 1 0 30268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1676037725
transform 1 0 37444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1676037725
transform 1 0 38548 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1676037725
transform 1 0 31004 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1676037725
transform 1 0 38824 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1676037725
transform 1 0 36064 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1676037725
transform 1 0 33580 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1676037725
transform 1 0 42596 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1676037725
transform 1 0 44528 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1676037725
transform 1 0 41308 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1676037725
transform 1 0 42596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1676037725
transform 1 0 26956 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0818_
timestamp 1676037725
transform 1 0 42780 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0824_
timestamp 1676037725
transform 1 0 36984 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1676037725
transform 1 0 55752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1676037725
transform 1 0 58052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1676037725
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0828_
timestamp 1676037725
transform 1 0 33396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1676037725
transform 1 0 40020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0831_
timestamp 1676037725
transform 1 0 56304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1676037725
transform 1 0 57040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0833_
timestamp 1676037725
transform 1 0 35052 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1676037725
transform 1 0 34132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0835_
timestamp 1676037725
transform 1 0 33856 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1676037725
transform 1 0 56120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1676037725
transform 1 0 43332 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0839_
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1676037725
transform 1 0 35052 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1676037725
transform 1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 1676037725
transform 1 0 57224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0844_
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1676037725
transform 1 0 34224 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0846_
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0847_
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0848_
timestamp 1676037725
transform 1 0 56764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0849_
timestamp 1676037725
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0853_
timestamp 1676037725
transform 1 0 44436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41676 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0855_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1676037725
transform 1 0 46644 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1676037725
transform 1 0 47748 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1676037725
transform 1 0 45172 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0860_
timestamp 1676037725
transform 1 0 46184 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform 1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0863_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0864_
timestamp 1676037725
transform 1 0 34960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0867_
timestamp 1676037725
transform 1 0 35052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1676037725
transform 1 0 39284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0870_
timestamp 1676037725
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1676037725
transform 1 0 43976 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0872_
timestamp 1676037725
transform 1 0 44344 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0873_
timestamp 1676037725
transform 1 0 33488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1676037725
transform 1 0 40020 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1676037725
transform 1 0 41124 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0877_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1676037725
transform 1 0 40204 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1676037725
transform 1 0 38640 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1676037725
transform 1 0 41492 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1676037725
transform 1 0 27324 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1676037725
transform 1 0 43700 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1676037725
transform 1 0 45172 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0886_
timestamp 1676037725
transform 1 0 36064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1676037725
transform 1 0 49036 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1676037725
transform 1 0 50324 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0889_
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0890_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1676037725
transform 1 0 42872 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1676037725
transform 1 0 42688 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1676037725
transform 1 0 40204 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0894_
timestamp 1676037725
transform 1 0 42688 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1676037725
transform 1 0 42872 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0896_
timestamp 1676037725
transform 1 0 30176 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0897_
timestamp 1676037725
transform 1 0 47840 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1676037725
transform 1 0 48852 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1676037725
transform 1 0 40664 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1676037725
transform 1 0 43608 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0902_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1676037725
transform 1 0 47840 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1676037725
transform 1 0 48116 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0905_
timestamp 1676037725
transform 1 0 42412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0906_
timestamp 1676037725
transform 1 0 45172 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1676037725
transform 1 0 45356 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0908_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0909_
timestamp 1676037725
transform 1 0 33764 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1676037725
transform 1 0 48852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1676037725
transform 1 0 50048 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0912_
timestamp 1676037725
transform 1 0 35328 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1676037725
transform 1 0 47104 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1676037725
transform 1 0 49128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0916_
timestamp 1676037725
transform 1 0 35512 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1676037725
transform 1 0 48116 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1676037725
transform 1 0 47472 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0919_
timestamp 1676037725
transform 1 0 38640 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1676037725
transform 1 0 43884 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1676037725
transform 1 0 40940 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_2  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34224 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0926_
timestamp 1676037725
transform 1 0 36340 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1676037725
transform 1 0 38640 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1676037725
transform 1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0930_
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0933_
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1676037725
transform 1 0 15364 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0939_
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0940_
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1676037725
transform 1 0 10028 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0946_
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0949_
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0950_
timestamp 1676037725
transform 1 0 13800 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _0951_
timestamp 1676037725
transform 1 0 14352 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0955_
timestamp 1676037725
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0957_
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1676037725
transform 1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1676037725
transform 1 0 20884 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1676037725
transform 1 0 20056 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1676037725
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0964_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0965_
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0967_
timestamp 1676037725
transform 1 0 22448 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0969_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0971_
timestamp 1676037725
transform 1 0 18124 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0972_
timestamp 1676037725
transform 1 0 22172 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0973_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0974_
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0975_
timestamp 1676037725
transform 1 0 23000 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0977_
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0978_
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0979_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0980_
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1676037725
transform 1 0 25576 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0982_
timestamp 1676037725
transform 1 0 26036 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1676037725
transform 1 0 30360 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 31004 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 29808 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 25760 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35880 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0993_
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0994_
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0995_
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0996_
timestamp 1676037725
transform 1 0 30912 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform 1 0 22448 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1676037725
transform 1 0 36156 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1004_
timestamp 1676037725
transform 1 0 35880 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1676037725
transform 1 0 29900 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1008_
timestamp 1676037725
transform 1 0 40020 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1009_
timestamp 1676037725
transform 1 0 28428 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1010_
timestamp 1676037725
transform 1 0 38732 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 30360 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1012_
timestamp 1676037725
transform 1 0 40480 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1013_
timestamp 1676037725
transform 1 0 35052 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1676037725
transform 1 0 31464 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1676037725
transform 1 0 34224 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 56856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 34868 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 32016 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 25760 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 25576 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 29532 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 27140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 27416 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 25852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 27048 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 27600 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1676037725
transform 1 0 31556 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1033_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 27600 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1035_
timestamp 1676037725
transform 1 0 37812 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1037_
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1676037725
transform 1 0 33672 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1039_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 35512 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1041_
timestamp 1676037725
transform 1 0 42596 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1042_
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1043_
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1044_
timestamp 1676037725
transform 1 0 42596 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1047_
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 25208 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 56856 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 56856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 56856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1052_
timestamp 1676037725
transform 1 0 37996 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 56856 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1054_
timestamp 1676037725
transform 1 0 42780 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 45356 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1057_
timestamp 1676037725
transform 1 0 34960 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1058_
timestamp 1676037725
transform 1 0 35144 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 44436 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1060_
timestamp 1676037725
transform 1 0 38824 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1061_
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1676037725
transform 1 0 44160 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1063_
timestamp 1676037725
transform 1 0 48392 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1064_
timestamp 1676037725
transform 1 0 43884 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1676037725
transform 1 0 42872 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1066_
timestamp 1676037725
transform 1 0 48116 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1676037725
transform 1 0 42872 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1068_
timestamp 1676037725
transform 1 0 48116 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1676037725
transform 1 0 45448 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1676037725
transform 1 0 48484 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1676037725
transform 1 0 50324 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1073_
timestamp 1676037725
transform 1 0 41400 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1074_
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1075_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1078_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1079_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1080_
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1081_
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1082_
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1089_
timestamp 1676037725
transform 1 0 17204 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1676037725
transform 1 0 17296 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1094_
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1095_
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1097_
timestamp 1676037725
transform 1 0 19780 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1098_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _1121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1676037725
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1676037725
transform 1 0 38916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1128_
timestamp 1676037725
transform 1 0 38548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1129_
timestamp 1676037725
transform 1 0 40020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1676037725
transform 1 0 38916 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1131_
timestamp 1676037725
transform 1 0 41492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1132_
timestamp 1676037725
transform 1 0 40756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1133_
timestamp 1676037725
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1676037725
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1135_
timestamp 1676037725
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41676 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1676037725
transform 1 0 31188 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1676037725
transform 1 0 31188 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1676037725
transform 1 0 41584 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout413 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 44160 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout414 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout415
timestamp 1676037725
transform 1 0 19504 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout416 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39284 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout417
timestamp 1676037725
transform 1 0 44528 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout418
timestamp 1676037725
transform 1 0 42688 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout419
timestamp 1676037725
transform 1 0 46276 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout420
timestamp 1676037725
transform 1 0 43608 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout421 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout422
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout423
timestamp 1676037725
transform 1 0 43792 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout424
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout425
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout426
timestamp 1676037725
transform 1 0 37352 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout427
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout429 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout430
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout431
timestamp 1676037725
transform 1 0 20516 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout432
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout433 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout434
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout435
timestamp 1676037725
transform 1 0 40664 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout436
timestamp 1676037725
transform 1 0 36064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  fanout437
timestamp 1676037725
transform 1 0 23184 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout438
timestamp 1676037725
transform 1 0 37720 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout439
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout440
timestamp 1676037725
transform 1 0 18584 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout441
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout442
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout443
timestamp 1676037725
transform 1 0 21068 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout444
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout445
timestamp 1676037725
transform 1 0 23644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout446
timestamp 1676037725
transform 1 0 21804 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout447
timestamp 1676037725
transform 1 0 21988 0 -1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout448
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout449
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout450
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout451
timestamp 1676037725
transform 1 0 17020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout452
timestamp 1676037725
transform 1 0 35604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout453
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout454
timestamp 1676037725
transform 1 0 35972 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout455
timestamp 1676037725
transform 1 0 18400 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout456
timestamp 1676037725
transform 1 0 20792 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout457
timestamp 1676037725
transform 1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout458
timestamp 1676037725
transform 1 0 31280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout459
timestamp 1676037725
transform 1 0 13248 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout460
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout461
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout462
timestamp 1676037725
transform 1 0 19412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout463
timestamp 1676037725
transform 1 0 20332 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout464
timestamp 1676037725
transform 1 0 35236 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout465
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout466
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout467
timestamp 1676037725
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout468
timestamp 1676037725
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout469
timestamp 1676037725
transform 1 0 13064 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout470
timestamp 1676037725
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout471
timestamp 1676037725
transform 1 0 15640 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout472
timestamp 1676037725
transform 1 0 27416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout473
timestamp 1676037725
transform 1 0 36156 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout474
timestamp 1676037725
transform 1 0 34868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout475
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout476
timestamp 1676037725
transform 1 0 41768 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout477
timestamp 1676037725
transform 1 0 35972 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout478
timestamp 1676037725
transform 1 0 33856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout479
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout480
timestamp 1676037725
transform 1 0 38640 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout481
timestamp 1676037725
transform 1 0 37904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout482
timestamp 1676037725
transform 1 0 43240 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout483
timestamp 1676037725
transform 1 0 41400 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout484
timestamp 1676037725
transform 1 0 43792 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout485
timestamp 1676037725
transform 1 0 43240 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout486
timestamp 1676037725
transform 1 0 42596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout487
timestamp 1676037725
transform 1 0 56488 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__bufbuf_16  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28796 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold2
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold3
timestamp 1676037725
transform 1 0 31280 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold4
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold5
timestamp 1676037725
transform 1 0 30268 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold6
timestamp 1676037725
transform 1 0 24288 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold7
timestamp 1676037725
transform 1 0 32292 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold8
timestamp 1676037725
transform 1 0 21712 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold9
timestamp 1676037725
transform 1 0 27968 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold10
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold11
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold12
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold13
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold14
timestamp 1676037725
transform 1 0 16560 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold15
timestamp 1676037725
transform 1 0 23736 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold16
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold17
timestamp 1676037725
transform 1 0 25576 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold18
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold19
timestamp 1676037725
transform 1 0 21712 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold20
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold21
timestamp 1676037725
transform 1 0 31832 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold22
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold23
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold24
timestamp 1676037725
transform 1 0 21712 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold25
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold26
timestamp 1676037725
transform 1 0 26864 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold27
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold28
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold29
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold30
timestamp 1676037725
transform 1 0 16560 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold31
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold32
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold33
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold34
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold35
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold36
timestamp 1676037725
transform 1 0 21344 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold37
timestamp 1676037725
transform 1 0 26312 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold38
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold39
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold40
timestamp 1676037725
transform 1 0 28244 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold41
timestamp 1676037725
transform 1 0 24288 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold42
timestamp 1676037725
transform 1 0 24748 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold43
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold44
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold45
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold46
timestamp 1676037725
transform 1 0 19136 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold47
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold48
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold49
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold50
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold51
timestamp 1676037725
transform 1 0 24288 0 -1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold52
timestamp 1676037725
transform 1 0 13984 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold53
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold54
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold55
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold56
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold57
timestamp 1676037725
transform 1 0 26220 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold58
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold59
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold60
timestamp 1676037725
transform 1 0 31372 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold61
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold62
timestamp 1676037725
transform 1 0 32568 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold63
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold64
timestamp 1676037725
transform 1 0 22816 0 -1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold65
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold66
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold67
timestamp 1676037725
transform 1 0 31280 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold68
timestamp 1676037725
transform 1 0 26496 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold69
timestamp 1676037725
transform 1 0 24288 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold70
timestamp 1676037725
transform 1 0 26864 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold71
timestamp 1676037725
transform 1 0 27876 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold72
timestamp 1676037725
transform 1 0 28152 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold73
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold74
timestamp 1676037725
transform 1 0 29440 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1676037725
transform 1 0 40204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 41492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 41124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform 1 0 41492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1676037725
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 46460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 42596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 44344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 44988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 47656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 45172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 46460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1676037725
transform 1 0 40388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1676037725
transform 1 0 44988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1676037725
transform 1 0 40756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1676037725
transform 1 0 43332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1676037725
transform 1 0 39284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 54096 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1676037725
transform 1 0 54648 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input30
timestamp 1676037725
transform 1 0 55476 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1676037725
transform 1 0 56396 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 56856 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1676037725
transform 1 0 58052 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1676037725
transform 1 0 57868 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 57132 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 48392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 50324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 49036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 51796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1676037725
transform 1 0 45540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1676037725
transform 1 0 51796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1676037725
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 50600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1676037725
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1676037725
transform 1 0 51428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1676037725
transform 1 0 52532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 49128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 50324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input57
timestamp 1676037725
transform 1 0 45632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 46552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 46184 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1676037725
transform 1 0 46736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 47748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 13432 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1676037725
transform 1 0 20424 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1676037725
transform 1 0 21160 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1676037725
transform 1 0 22264 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 23184 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 23736 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 24472 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input70
timestamp 1676037725
transform 1 0 25208 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1676037725
transform 1 0 26128 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1676037725
transform 1 0 27140 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 27416 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 14168 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input75
timestamp 1676037725
transform 1 0 28152 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 28888 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1676037725
transform 1 0 29716 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1676037725
transform 1 0 30360 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1676037725
transform 1 0 31096 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1676037725
transform 1 0 32292 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1676037725
transform 1 0 33212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input82
timestamp 1676037725
transform 1 0 14904 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1676037725
transform 1 0 15640 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1676037725
transform 1 0 16008 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1676037725
transform 1 0 17112 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1676037725
transform 1 0 17848 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1676037725
transform 1 0 18584 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1676037725
transform 1 0 19320 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1676037725
transform 1 0 19688 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input95
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1676037725
transform 1 0 1564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1676037725
transform 1 0 1564 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1676037725
transform 1 0 1564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform 1 0 1564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 1564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1676037725
transform 1 0 1564 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 1564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input104
timestamp 1676037725
transform 1 0 1564 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input105
timestamp 1676037725
transform 1 0 1564 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 1564 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input107
timestamp 1676037725
transform 1 0 1564 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input108
timestamp 1676037725
transform 1 0 1564 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input109
timestamp 1676037725
transform 1 0 2760 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input111
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1676037725
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1676037725
transform 1 0 1564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1676037725
transform 1 0 33948 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1676037725
transform 1 0 41492 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1676037725
transform 1 0 41400 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input121
timestamp 1676037725
transform 1 0 42596 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1676037725
transform 1 0 43516 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1676037725
transform 1 0 44252 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1676037725
transform 1 0 45172 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1676037725
transform 1 0 45908 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1676037725
transform 1 0 46644 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1676037725
transform 1 0 46552 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1676037725
transform 1 0 47748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1676037725
transform 1 0 34868 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1676037725
transform 1 0 48484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1676037725
transform 1 0 49220 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input132
timestamp 1676037725
transform 1 0 50324 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1676037725
transform 1 0 50232 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1676037725
transform 1 0 51244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input135
timestamp 1676037725
transform 1 0 51980 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1676037725
transform 1 0 52900 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1676037725
transform 1 0 35604 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input138
timestamp 1676037725
transform 1 0 36340 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1676037725
transform 1 0 36248 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1676037725
transform 1 0 37444 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1676037725
transform 1 0 38180 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input142
timestamp 1676037725
transform 1 0 38916 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input143
timestamp 1676037725
transform 1 0 40020 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input144
timestamp 1676037725
transform 1 0 40756 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1676037725
transform 1 0 58052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input146
timestamp 1676037725
transform 1 0 56120 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input147
timestamp 1676037725
transform 1 0 57224 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input148
timestamp 1676037725
transform 1 0 57868 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input149
timestamp 1676037725
transform 1 0 57868 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input150
timestamp 1676037725
transform 1 0 57868 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input151
timestamp 1676037725
transform 1 0 58052 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1676037725
transform 1 0 58052 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1676037725
transform 1 0 58052 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1676037725
transform 1 0 57132 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input155
timestamp 1676037725
transform 1 0 56396 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1676037725
transform 1 0 55384 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input157
timestamp 1676037725
transform 1 0 6624 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input158
timestamp 1676037725
transform 1 0 7544 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1676037725
transform 1 0 8280 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input160
timestamp 1676037725
transform 1 0 9108 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1676037725
transform 1 0 9752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1676037725
transform 1 0 10120 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1676037725
transform 1 0 10856 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1676037725
transform 1 0 11960 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input166
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input168
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1676037725
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1676037725
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input174
timestamp 1676037725
transform 1 0 1564 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input175
timestamp 1676037725
transform 1 0 2300 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input176
timestamp 1676037725
transform 1 0 2484 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input177
timestamp 1676037725
transform 1 0 3128 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input178
timestamp 1676037725
transform 1 0 3864 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1676037725
transform 1 0 4600 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1676037725
transform 1 0 5336 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input181
timestamp 1676037725
transform 1 0 5520 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1676037725
transform 1 0 38548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input183
timestamp 1676037725
transform 1 0 40020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input184
timestamp 1676037725
transform 1 0 41124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input185
timestamp 1676037725
transform 1 0 39652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input186
timestamp 1676037725
transform 1 0 1564 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input187
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input188
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input189
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1676037725
transform 1 0 1564 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input191
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input192
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input193
timestamp 1676037725
transform 1 0 1564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input194
timestamp 1676037725
transform 1 0 52900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input195
timestamp 1676037725
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input196
timestamp 1676037725
transform 1 0 54004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input197
timestamp 1676037725
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input198
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input199
timestamp 1676037725
transform 1 0 53636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input200
timestamp 1676037725
transform 1 0 54556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input201
timestamp 1676037725
transform 1 0 54372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input202
timestamp 1676037725
transform 1 0 55108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input203
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input204
timestamp 1676037725
transform 1 0 55476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input205
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1676037725
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1676037725
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1676037725
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1676037725
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1676037725
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1676037725
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1676037725
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1676037725
transform 1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1676037725
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1676037725
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1676037725
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1676037725
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input232
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input233
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input234
timestamp 1676037725
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1676037725
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1676037725
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1676037725
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input241
timestamp 1676037725
transform 1 0 12696 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input242
timestamp 1676037725
transform 1 0 1564 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input243
timestamp 1676037725
transform 1 0 53176 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input244
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input245
timestamp 1676037725
transform 1 0 57132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input246
timestamp 1676037725
transform 1 0 57868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input247
timestamp 1676037725
transform 1 0 56948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input248
timestamp 1676037725
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input249
timestamp 1676037725
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input250
timestamp 1676037725
transform 1 0 58052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input251
timestamp 1676037725
transform 1 0 58052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input252
timestamp 1676037725
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input253
timestamp 1676037725
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input254
timestamp 1676037725
transform 1 0 56948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input255
timestamp 1676037725
transform 1 0 58052 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input256
timestamp 1676037725
transform 1 0 56948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input257
timestamp 1676037725
transform 1 0 58052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input258
timestamp 1676037725
transform 1 0 56948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input259
timestamp 1676037725
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input260
timestamp 1676037725
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input261
timestamp 1676037725
transform 1 0 58052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input262
timestamp 1676037725
transform 1 0 58052 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input263
timestamp 1676037725
transform 1 0 56948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input264
timestamp 1676037725
transform 1 0 57868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input265
timestamp 1676037725
transform 1 0 56948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input266
timestamp 1676037725
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input267
timestamp 1676037725
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input268
timestamp 1676037725
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input269
timestamp 1676037725
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input270
timestamp 1676037725
transform 1 0 57040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input271
timestamp 1676037725
transform 1 0 58052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input272
timestamp 1676037725
transform 1 0 58052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input273
timestamp 1676037725
transform 1 0 56948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input274
timestamp 1676037725
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input275
timestamp 1676037725
transform 1 0 56948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input276
timestamp 1676037725
transform 1 0 58052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input277
timestamp 1676037725
transform 1 0 58052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input278
timestamp 1676037725
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input279
timestamp 1676037725
transform 1 0 58052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  multiplexer_488 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_489
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_490
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_491
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_492
timestamp 1676037725
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_493
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_494
timestamp 1676037725
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_495
timestamp 1676037725
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_496
timestamp 1676037725
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_497
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_498
timestamp 1676037725
transform 1 0 58144 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_499
timestamp 1676037725
transform 1 0 58144 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_500
timestamp 1676037725
transform 1 0 58144 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_501
timestamp 1676037725
transform 1 0 58144 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_502
timestamp 1676037725
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_503
timestamp 1676037725
transform 1 0 36708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_504
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_505
timestamp 1676037725
transform 1 0 34132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_506
timestamp 1676037725
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_507
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output281
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output282
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output283
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output284
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output285
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output286
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output287
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output288
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output289
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output290
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output291
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output292
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output293
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output294
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output295
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output296
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output297
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output298
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output299
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output300
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output301
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output302
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output303
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output304
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output305
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output306
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output307
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output308
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output309
timestamp 1676037725
transform 1 0 18768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output310
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output311
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output312
timestamp 1676037725
transform 1 0 34132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output313
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output314
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output315
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output316
timestamp 1676037725
transform 1 0 27416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output317
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output318
timestamp 1676037725
transform 1 0 28704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output319
timestamp 1676037725
transform 1 0 30084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output320
timestamp 1676037725
transform 1 0 31004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output321
timestamp 1676037725
transform 1 0 31280 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output322
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output323
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output324
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output325
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output326
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output327
timestamp 1676037725
transform 1 0 33856 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output328
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output329
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output330
timestamp 1676037725
transform 1 0 35052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output331
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output332
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output333
timestamp 1676037725
transform 1 0 35052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output334
timestamp 1676037725
transform 1 0 36432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output335
timestamp 1676037725
transform 1 0 37812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output336
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output337
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output338
timestamp 1676037725
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output339
timestamp 1676037725
transform 1 0 10672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output340
timestamp 1676037725
transform 1 0 15640 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output341
timestamp 1676037725
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output342
timestamp 1676037725
transform 1 0 17480 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output343
timestamp 1676037725
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output344
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output345
timestamp 1676037725
transform 1 0 14904 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output346
timestamp 1676037725
transform 1 0 16560 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output347
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output348
timestamp 1676037725
transform 1 0 17572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output349
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output350
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output351
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output352
timestamp 1676037725
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output353
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output354
timestamp 1676037725
transform 1 0 12144 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output355
timestamp 1676037725
transform 1 0 14720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output356
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output357
timestamp 1676037725
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output358
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output359
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output360
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output361
timestamp 1676037725
transform 1 0 18492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output362
timestamp 1676037725
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output363
timestamp 1676037725
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output364
timestamp 1676037725
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output365
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output366
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output367
timestamp 1676037725
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output368
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output369
timestamp 1676037725
transform 1 0 56396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output370
timestamp 1676037725
transform 1 0 56396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output371
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output372
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output373
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output374
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output375
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output376
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output377
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output378
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output379
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output380
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output381
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output382
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output383
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output384
timestamp 1676037725
transform 1 0 55936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output385
timestamp 1676037725
transform 1 0 57868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output386
timestamp 1676037725
transform 1 0 57868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output387
timestamp 1676037725
transform 1 0 57868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output388
timestamp 1676037725
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output389
timestamp 1676037725
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output390
timestamp 1676037725
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output391
timestamp 1676037725
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output392
timestamp 1676037725
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output393
timestamp 1676037725
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output394
timestamp 1676037725
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output395
timestamp 1676037725
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output396
timestamp 1676037725
transform 1 0 57040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output397
timestamp 1676037725
transform 1 0 57868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output398
timestamp 1676037725
transform 1 0 57868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output399
timestamp 1676037725
transform 1 0 56948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output400
timestamp 1676037725
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output401
timestamp 1676037725
transform 1 0 56948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output402
timestamp 1676037725
transform 1 0 57868 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output403
timestamp 1676037725
transform 1 0 56948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output404
timestamp 1676037725
transform 1 0 57868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output405
timestamp 1676037725
transform 1 0 57868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output406
timestamp 1676037725
transform 1 0 57868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output407
timestamp 1676037725
transform 1 0 57868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output408
timestamp 1676037725
transform 1 0 57868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output409
timestamp 1676037725
transform 1 0 57868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output410
timestamp 1676037725
transform 1 0 57868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output411
timestamp 1676037725
transform 1 0 57868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output412
timestamp 1676037725
transform 1 0 57868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire428
timestamp 1676037725
transform 1 0 22448 0 1 32640
box -38 -48 866 592
<< labels >>
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 dsi_all[27]
port 20 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 dsi_all[2]
port 21 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 dsi_all[3]
port 22 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 dsi_all[4]
port 23 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 dsi_all[5]
port 24 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 dsi_all[6]
port 25 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 dsi_all[7]
port 26 nsew signal tristate
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 dsi_all[8]
port 27 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 dsi_all[9]
port 28 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 dso_6502[0]
port 29 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 dso_6502[10]
port 30 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 dso_6502[11]
port 31 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 dso_6502[12]
port 32 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 dso_6502[13]
port 33 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 dso_6502[14]
port 34 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 dso_6502[15]
port 35 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 dso_6502[16]
port 36 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 dso_6502[17]
port 37 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 dso_6502[18]
port 38 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 dso_6502[19]
port 39 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 dso_6502[1]
port 40 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 dso_6502[20]
port 41 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 dso_6502[21]
port 42 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 dso_6502[22]
port 43 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 dso_6502[23]
port 44 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 dso_6502[24]
port 45 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 dso_6502[25]
port 46 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 dso_6502[26]
port 47 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 dso_6502[2]
port 48 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 dso_6502[3]
port 49 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 dso_6502[4]
port 50 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 dso_6502[5]
port 51 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 dso_6502[6]
port 52 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 dso_6502[7]
port 53 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 dso_6502[8]
port 54 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 dso_6502[9]
port 55 nsew signal input
flabel metal2 s 53838 63200 53894 64000 0 FreeSans 224 90 0 0 dso_LCD[0]
port 56 nsew signal input
flabel metal2 s 54574 63200 54630 64000 0 FreeSans 224 90 0 0 dso_LCD[1]
port 57 nsew signal input
flabel metal2 s 55310 63200 55366 64000 0 FreeSans 224 90 0 0 dso_LCD[2]
port 58 nsew signal input
flabel metal2 s 56046 63200 56102 64000 0 FreeSans 224 90 0 0 dso_LCD[3]
port 59 nsew signal input
flabel metal2 s 56782 63200 56838 64000 0 FreeSans 224 90 0 0 dso_LCD[4]
port 60 nsew signal input
flabel metal2 s 57518 63200 57574 64000 0 FreeSans 224 90 0 0 dso_LCD[5]
port 61 nsew signal input
flabel metal2 s 58254 63200 58310 64000 0 FreeSans 224 90 0 0 dso_LCD[6]
port 62 nsew signal input
flabel metal2 s 58990 63200 59046 64000 0 FreeSans 224 90 0 0 dso_LCD[7]
port 63 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 dso_as1802[0]
port 64 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 dso_as1802[10]
port 65 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 dso_as1802[11]
port 66 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 dso_as1802[12]
port 67 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 dso_as1802[13]
port 68 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 dso_as1802[14]
port 69 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 dso_as1802[15]
port 70 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 dso_as1802[16]
port 71 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 dso_as1802[17]
port 72 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 dso_as1802[18]
port 73 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 dso_as1802[19]
port 74 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 dso_as1802[1]
port 75 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 dso_as1802[20]
port 76 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 dso_as1802[21]
port 77 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 dso_as1802[22]
port 78 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 dso_as1802[23]
port 79 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 dso_as1802[24]
port 80 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 dso_as1802[25]
port 81 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 dso_as1802[26]
port 82 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 dso_as1802[2]
port 83 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 dso_as1802[3]
port 84 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 dso_as1802[4]
port 85 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 dso_as1802[5]
port 86 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 dso_as1802[6]
port 87 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 dso_as1802[7]
port 88 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 dso_as1802[8]
port 89 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 dso_as1802[9]
port 90 nsew signal input
flabel metal2 s 13358 63200 13414 64000 0 FreeSans 224 90 0 0 dso_as2650[0]
port 91 nsew signal input
flabel metal2 s 20718 63200 20774 64000 0 FreeSans 224 90 0 0 dso_as2650[10]
port 92 nsew signal input
flabel metal2 s 21454 63200 21510 64000 0 FreeSans 224 90 0 0 dso_as2650[11]
port 93 nsew signal input
flabel metal2 s 22190 63200 22246 64000 0 FreeSans 224 90 0 0 dso_as2650[12]
port 94 nsew signal input
flabel metal2 s 22926 63200 22982 64000 0 FreeSans 224 90 0 0 dso_as2650[13]
port 95 nsew signal input
flabel metal2 s 23662 63200 23718 64000 0 FreeSans 224 90 0 0 dso_as2650[14]
port 96 nsew signal input
flabel metal2 s 24398 63200 24454 64000 0 FreeSans 224 90 0 0 dso_as2650[15]
port 97 nsew signal input
flabel metal2 s 25134 63200 25190 64000 0 FreeSans 224 90 0 0 dso_as2650[16]
port 98 nsew signal input
flabel metal2 s 25870 63200 25926 64000 0 FreeSans 224 90 0 0 dso_as2650[17]
port 99 nsew signal input
flabel metal2 s 26606 63200 26662 64000 0 FreeSans 224 90 0 0 dso_as2650[18]
port 100 nsew signal input
flabel metal2 s 27342 63200 27398 64000 0 FreeSans 224 90 0 0 dso_as2650[19]
port 101 nsew signal input
flabel metal2 s 14094 63200 14150 64000 0 FreeSans 224 90 0 0 dso_as2650[1]
port 102 nsew signal input
flabel metal2 s 28078 63200 28134 64000 0 FreeSans 224 90 0 0 dso_as2650[20]
port 103 nsew signal input
flabel metal2 s 28814 63200 28870 64000 0 FreeSans 224 90 0 0 dso_as2650[21]
port 104 nsew signal input
flabel metal2 s 29550 63200 29606 64000 0 FreeSans 224 90 0 0 dso_as2650[22]
port 105 nsew signal input
flabel metal2 s 30286 63200 30342 64000 0 FreeSans 224 90 0 0 dso_as2650[23]
port 106 nsew signal input
flabel metal2 s 31022 63200 31078 64000 0 FreeSans 224 90 0 0 dso_as2650[24]
port 107 nsew signal input
flabel metal2 s 31758 63200 31814 64000 0 FreeSans 224 90 0 0 dso_as2650[25]
port 108 nsew signal input
flabel metal2 s 32494 63200 32550 64000 0 FreeSans 224 90 0 0 dso_as2650[26]
port 109 nsew signal input
flabel metal2 s 14830 63200 14886 64000 0 FreeSans 224 90 0 0 dso_as2650[2]
port 110 nsew signal input
flabel metal2 s 15566 63200 15622 64000 0 FreeSans 224 90 0 0 dso_as2650[3]
port 111 nsew signal input
flabel metal2 s 16302 63200 16358 64000 0 FreeSans 224 90 0 0 dso_as2650[4]
port 112 nsew signal input
flabel metal2 s 17038 63200 17094 64000 0 FreeSans 224 90 0 0 dso_as2650[5]
port 113 nsew signal input
flabel metal2 s 17774 63200 17830 64000 0 FreeSans 224 90 0 0 dso_as2650[6]
port 114 nsew signal input
flabel metal2 s 18510 63200 18566 64000 0 FreeSans 224 90 0 0 dso_as2650[7]
port 115 nsew signal input
flabel metal2 s 19246 63200 19302 64000 0 FreeSans 224 90 0 0 dso_as2650[8]
port 116 nsew signal input
flabel metal2 s 19982 63200 20038 64000 0 FreeSans 224 90 0 0 dso_as2650[9]
port 117 nsew signal input
flabel metal3 s 0 42712 800 42832 0 FreeSans 480 0 0 0 dso_as512512512[0]
port 118 nsew signal input
flabel metal3 s 0 49512 800 49632 0 FreeSans 480 0 0 0 dso_as512512512[10]
port 119 nsew signal input
flabel metal3 s 0 50192 800 50312 0 FreeSans 480 0 0 0 dso_as512512512[11]
port 120 nsew signal input
flabel metal3 s 0 50872 800 50992 0 FreeSans 480 0 0 0 dso_as512512512[12]
port 121 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 dso_as512512512[13]
port 122 nsew signal input
flabel metal3 s 0 52232 800 52352 0 FreeSans 480 0 0 0 dso_as512512512[14]
port 123 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 dso_as512512512[15]
port 124 nsew signal input
flabel metal3 s 0 53592 800 53712 0 FreeSans 480 0 0 0 dso_as512512512[16]
port 125 nsew signal input
flabel metal3 s 0 54272 800 54392 0 FreeSans 480 0 0 0 dso_as512512512[17]
port 126 nsew signal input
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 dso_as512512512[18]
port 127 nsew signal input
flabel metal3 s 0 55632 800 55752 0 FreeSans 480 0 0 0 dso_as512512512[19]
port 128 nsew signal input
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 dso_as512512512[1]
port 129 nsew signal input
flabel metal3 s 0 56312 800 56432 0 FreeSans 480 0 0 0 dso_as512512512[20]
port 130 nsew signal input
flabel metal3 s 0 56992 800 57112 0 FreeSans 480 0 0 0 dso_as512512512[21]
port 131 nsew signal input
flabel metal3 s 0 57672 800 57792 0 FreeSans 480 0 0 0 dso_as512512512[22]
port 132 nsew signal input
flabel metal3 s 0 58352 800 58472 0 FreeSans 480 0 0 0 dso_as512512512[23]
port 133 nsew signal input
flabel metal3 s 0 59032 800 59152 0 FreeSans 480 0 0 0 dso_as512512512[24]
port 134 nsew signal input
flabel metal3 s 0 59712 800 59832 0 FreeSans 480 0 0 0 dso_as512512512[25]
port 135 nsew signal input
flabel metal3 s 0 60392 800 60512 0 FreeSans 480 0 0 0 dso_as512512512[26]
port 136 nsew signal input
flabel metal3 s 0 61072 800 61192 0 FreeSans 480 0 0 0 dso_as512512512[27]
port 137 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 dso_as512512512[2]
port 138 nsew signal input
flabel metal3 s 0 44752 800 44872 0 FreeSans 480 0 0 0 dso_as512512512[3]
port 139 nsew signal input
flabel metal3 s 0 45432 800 45552 0 FreeSans 480 0 0 0 dso_as512512512[4]
port 140 nsew signal input
flabel metal3 s 0 46112 800 46232 0 FreeSans 480 0 0 0 dso_as512512512[5]
port 141 nsew signal input
flabel metal3 s 0 46792 800 46912 0 FreeSans 480 0 0 0 dso_as512512512[6]
port 142 nsew signal input
flabel metal3 s 0 47472 800 47592 0 FreeSans 480 0 0 0 dso_as512512512[7]
port 143 nsew signal input
flabel metal3 s 0 48152 800 48272 0 FreeSans 480 0 0 0 dso_as512512512[8]
port 144 nsew signal input
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 dso_as512512512[9]
port 145 nsew signal input
flabel metal2 s 33230 63200 33286 64000 0 FreeSans 224 90 0 0 dso_as5401[0]
port 146 nsew signal input
flabel metal2 s 40590 63200 40646 64000 0 FreeSans 224 90 0 0 dso_as5401[10]
port 147 nsew signal input
flabel metal2 s 41326 63200 41382 64000 0 FreeSans 224 90 0 0 dso_as5401[11]
port 148 nsew signal input
flabel metal2 s 42062 63200 42118 64000 0 FreeSans 224 90 0 0 dso_as5401[12]
port 149 nsew signal input
flabel metal2 s 42798 63200 42854 64000 0 FreeSans 224 90 0 0 dso_as5401[13]
port 150 nsew signal input
flabel metal2 s 43534 63200 43590 64000 0 FreeSans 224 90 0 0 dso_as5401[14]
port 151 nsew signal input
flabel metal2 s 44270 63200 44326 64000 0 FreeSans 224 90 0 0 dso_as5401[15]
port 152 nsew signal input
flabel metal2 s 45006 63200 45062 64000 0 FreeSans 224 90 0 0 dso_as5401[16]
port 153 nsew signal input
flabel metal2 s 45742 63200 45798 64000 0 FreeSans 224 90 0 0 dso_as5401[17]
port 154 nsew signal input
flabel metal2 s 46478 63200 46534 64000 0 FreeSans 224 90 0 0 dso_as5401[18]
port 155 nsew signal input
flabel metal2 s 47214 63200 47270 64000 0 FreeSans 224 90 0 0 dso_as5401[19]
port 156 nsew signal input
flabel metal2 s 33966 63200 34022 64000 0 FreeSans 224 90 0 0 dso_as5401[1]
port 157 nsew signal input
flabel metal2 s 47950 63200 48006 64000 0 FreeSans 224 90 0 0 dso_as5401[20]
port 158 nsew signal input
flabel metal2 s 48686 63200 48742 64000 0 FreeSans 224 90 0 0 dso_as5401[21]
port 159 nsew signal input
flabel metal2 s 49422 63200 49478 64000 0 FreeSans 224 90 0 0 dso_as5401[22]
port 160 nsew signal input
flabel metal2 s 50158 63200 50214 64000 0 FreeSans 224 90 0 0 dso_as5401[23]
port 161 nsew signal input
flabel metal2 s 50894 63200 50950 64000 0 FreeSans 224 90 0 0 dso_as5401[24]
port 162 nsew signal input
flabel metal2 s 51630 63200 51686 64000 0 FreeSans 224 90 0 0 dso_as5401[25]
port 163 nsew signal input
flabel metal2 s 52366 63200 52422 64000 0 FreeSans 224 90 0 0 dso_as5401[26]
port 164 nsew signal input
flabel metal2 s 34702 63200 34758 64000 0 FreeSans 224 90 0 0 dso_as5401[2]
port 165 nsew signal input
flabel metal2 s 35438 63200 35494 64000 0 FreeSans 224 90 0 0 dso_as5401[3]
port 166 nsew signal input
flabel metal2 s 36174 63200 36230 64000 0 FreeSans 224 90 0 0 dso_as5401[4]
port 167 nsew signal input
flabel metal2 s 36910 63200 36966 64000 0 FreeSans 224 90 0 0 dso_as5401[5]
port 168 nsew signal input
flabel metal2 s 37646 63200 37702 64000 0 FreeSans 224 90 0 0 dso_as5401[6]
port 169 nsew signal input
flabel metal2 s 38382 63200 38438 64000 0 FreeSans 224 90 0 0 dso_as5401[7]
port 170 nsew signal input
flabel metal2 s 39118 63200 39174 64000 0 FreeSans 224 90 0 0 dso_as5401[8]
port 171 nsew signal input
flabel metal2 s 39854 63200 39910 64000 0 FreeSans 224 90 0 0 dso_as5401[9]
port 172 nsew signal input
flabel metal3 s 59200 56584 60000 56704 0 FreeSans 480 0 0 0 dso_counter[0]
port 173 nsew signal input
flabel metal3 s 59200 62024 60000 62144 0 FreeSans 480 0 0 0 dso_counter[10]
port 174 nsew signal input
flabel metal3 s 59200 62568 60000 62688 0 FreeSans 480 0 0 0 dso_counter[11]
port 175 nsew signal input
flabel metal3 s 59200 57128 60000 57248 0 FreeSans 480 0 0 0 dso_counter[1]
port 176 nsew signal input
flabel metal3 s 59200 57672 60000 57792 0 FreeSans 480 0 0 0 dso_counter[2]
port 177 nsew signal input
flabel metal3 s 59200 58216 60000 58336 0 FreeSans 480 0 0 0 dso_counter[3]
port 178 nsew signal input
flabel metal3 s 59200 58760 60000 58880 0 FreeSans 480 0 0 0 dso_counter[4]
port 179 nsew signal input
flabel metal3 s 59200 59304 60000 59424 0 FreeSans 480 0 0 0 dso_counter[5]
port 180 nsew signal input
flabel metal3 s 59200 59848 60000 59968 0 FreeSans 480 0 0 0 dso_counter[6]
port 181 nsew signal input
flabel metal3 s 59200 60392 60000 60512 0 FreeSans 480 0 0 0 dso_counter[7]
port 182 nsew signal input
flabel metal3 s 59200 60936 60000 61056 0 FreeSans 480 0 0 0 dso_counter[8]
port 183 nsew signal input
flabel metal3 s 59200 61480 60000 61600 0 FreeSans 480 0 0 0 dso_counter[9]
port 184 nsew signal input
flabel metal2 s 6734 63200 6790 64000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 185 nsew signal input
flabel metal2 s 7470 63200 7526 64000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 186 nsew signal input
flabel metal2 s 8206 63200 8262 64000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 187 nsew signal input
flabel metal2 s 8942 63200 8998 64000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 188 nsew signal input
flabel metal2 s 9678 63200 9734 64000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 189 nsew signal input
flabel metal2 s 10414 63200 10470 64000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 190 nsew signal input
flabel metal2 s 11150 63200 11206 64000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 191 nsew signal input
flabel metal2 s 11886 63200 11942 64000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 192 nsew signal input
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 193 nsew signal input
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 194 nsew signal input
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 195 nsew signal input
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 196 nsew signal input
flabel metal3 s 0 33192 800 33312 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 197 nsew signal input
flabel metal3 s 0 33872 800 33992 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 198 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 199 nsew signal input
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 200 nsew signal input
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 201 nsew signal input
flabel metal2 s 846 63200 902 64000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 202 nsew signal input
flabel metal2 s 1582 63200 1638 64000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 203 nsew signal input
flabel metal2 s 2318 63200 2374 64000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 204 nsew signal input
flabel metal2 s 3054 63200 3110 64000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 205 nsew signal input
flabel metal2 s 3790 63200 3846 64000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 206 nsew signal input
flabel metal2 s 4526 63200 4582 64000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 207 nsew signal input
flabel metal2 s 5262 63200 5318 64000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 208 nsew signal input
flabel metal2 s 5998 63200 6054 64000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 209 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 dso_nand
port 210 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 dso_posit[0]
port 211 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 dso_posit[1]
port 212 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 dso_posit[2]
port 213 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 dso_posit[3]
port 214 nsew signal input
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 215 nsew signal input
flabel metal3 s 0 37952 800 38072 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 216 nsew signal input
flabel metal3 s 0 38632 800 38752 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 217 nsew signal input
flabel metal3 s 0 39312 800 39432 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 218 nsew signal input
flabel metal3 s 0 39992 800 40112 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 219 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 220 nsew signal input
flabel metal3 s 0 41352 800 41472 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 221 nsew signal input
flabel metal3 s 0 42032 800 42152 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 222 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 dso_tune
port 223 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 dso_vgatest[0]
port 224 nsew signal input
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 dso_vgatest[1]
port 225 nsew signal input
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 dso_vgatest[2]
port 226 nsew signal input
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 dso_vgatest[3]
port 227 nsew signal input
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 dso_vgatest[4]
port 228 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 dso_vgatest[5]
port 229 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 dso_vgatest[6]
port 230 nsew signal input
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 dso_vgatest[7]
port 231 nsew signal input
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 dso_vgatest[8]
port 232 nsew signal input
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 dso_vgatest[9]
port 233 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 io_in[0]
port 234 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 io_in[10]
port 235 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 io_in[11]
port 236 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 io_in[12]
port 237 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 io_in[13]
port 238 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 io_in[14]
port 239 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 io_in[15]
port 240 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 io_in[16]
port 241 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 io_in[17]
port 242 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 io_in[18]
port 243 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 io_in[19]
port 244 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 io_in[1]
port 245 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_in[20]
port 246 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 io_in[21]
port 247 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 io_in[22]
port 248 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_in[23]
port 249 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 io_in[24]
port 250 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 io_in[25]
port 251 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 io_in[26]
port 252 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_in[27]
port 253 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 io_in[28]
port 254 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 io_in[29]
port 255 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 io_in[2]
port 256 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 io_in[30]
port 257 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 io_in[31]
port 258 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 io_in[32]
port 259 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 io_in[33]
port 260 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 io_in[34]
port 261 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 io_in[35]
port 262 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_in[36]
port 263 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 io_in[37]
port 264 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 io_in[3]
port 265 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 io_in[4]
port 266 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 io_in[5]
port 267 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 io_in[6]
port 268 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 io_in[7]
port 269 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 io_in[8]
port 270 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_in[9]
port 271 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 272 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 273 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 274 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 275 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 276 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 277 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 278 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 279 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 280 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 281 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 282 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 283 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 284 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 285 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 286 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 287 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 288 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 289 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 290 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 291 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 292 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 293 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 294 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 295 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 296 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 297 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 298 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 299 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 300 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 301 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 302 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 303 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 304 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 305 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 306 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 307 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 308 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 309 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 io_out[0]
port 310 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 io_out[10]
port 311 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 io_out[11]
port 312 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 io_out[12]
port 313 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_out[13]
port 314 nsew signal tristate
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 io_out[14]
port 315 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 io_out[15]
port 316 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 io_out[16]
port 317 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 io_out[17]
port 318 nsew signal tristate
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 io_out[18]
port 319 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 io_out[19]
port 320 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_out[1]
port 321 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 io_out[20]
port 322 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 io_out[21]
port 323 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 io_out[22]
port 324 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 io_out[23]
port 325 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 io_out[24]
port 326 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 io_out[25]
port 327 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 io_out[26]
port 328 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 io_out[27]
port 329 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 io_out[28]
port 330 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 io_out[29]
port 331 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 io_out[2]
port 332 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 io_out[30]
port 333 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 io_out[31]
port 334 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 io_out[32]
port 335 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 io_out[33]
port 336 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 io_out[34]
port 337 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 io_out[35]
port 338 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 io_out[36]
port 339 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 io_out[37]
port 340 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 io_out[3]
port 341 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 io_out[4]
port 342 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 io_out[5]
port 343 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 io_out[6]
port 344 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 io_out[7]
port 345 nsew signal tristate
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 io_out[8]
port 346 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 io_out[9]
port 347 nsew signal tristate
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 nand_dsi[0]
port 348 nsew signal tristate
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 nand_dsi[1]
port 349 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 oeb_6502
port 350 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 oeb_as1802
port 351 nsew signal input
flabel metal2 s 12622 63200 12678 64000 0 FreeSans 224 90 0 0 oeb_as2650
port 352 nsew signal input
flabel metal3 s 0 61752 800 61872 0 FreeSans 480 0 0 0 oeb_as512512512
port 353 nsew signal input
flabel metal2 s 53102 63200 53158 64000 0 FreeSans 224 90 0 0 oeb_as5401
port 354 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 oeb_mc14500
port 355 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 rst_6502
port 356 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 rst_LCD
port 357 nsew signal tristate
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 rst_as1802
port 358 nsew signal tristate
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 rst_as2650
port 359 nsew signal tristate
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 rst_as512512512
port 360 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 rst_as5401
port 361 nsew signal tristate
flabel metal3 s 0 25712 800 25832 0 FreeSans 480 0 0 0 rst_counter
port 362 nsew signal tristate
flabel metal3 s 0 26392 800 26512 0 FreeSans 480 0 0 0 rst_diceroll
port 363 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 rst_mc14500
port 364 nsew signal tristate
flabel metal3 s 0 27752 800 27872 0 FreeSans 480 0 0 0 rst_posit
port 365 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 rst_tbb1143
port 366 nsew signal tristate
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 rst_tune
port 367 nsew signal tristate
flabel metal3 s 0 29792 800 29912 0 FreeSans 480 0 0 0 rst_vgatest
port 368 nsew signal tristate
flabel metal4 s 4208 2128 4528 61520 0 FreeSans 1920 90 0 0 vccd1
port 369 nsew power bidirectional
flabel metal4 s 34928 2128 35248 61520 0 FreeSans 1920 90 0 0 vccd1
port 369 nsew power bidirectional
flabel metal4 s 19568 2128 19888 61520 0 FreeSans 1920 90 0 0 vssd1
port 370 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 61520 0 FreeSans 1920 90 0 0 vssd1
port 370 nsew ground bidirectional
flabel metal3 s 59200 1096 60000 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 371 nsew signal input
flabel metal3 s 59200 1640 60000 1760 0 FreeSans 480 0 0 0 wb_rst_i
port 372 nsew signal input
flabel metal3 s 59200 2184 60000 2304 0 FreeSans 480 0 0 0 wbs_ack_o
port 373 nsew signal tristate
flabel metal3 s 59200 4360 60000 4480 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 374 nsew signal input
flabel metal3 s 59200 20680 60000 20800 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 375 nsew signal input
flabel metal3 s 59200 22312 60000 22432 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 376 nsew signal input
flabel metal3 s 59200 23944 60000 24064 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 377 nsew signal input
flabel metal3 s 59200 25576 60000 25696 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 378 nsew signal input
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 379 nsew signal input
flabel metal3 s 59200 28840 60000 28960 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 380 nsew signal input
flabel metal3 s 59200 30472 60000 30592 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 381 nsew signal input
flabel metal3 s 59200 32104 60000 32224 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 382 nsew signal input
flabel metal3 s 59200 33736 60000 33856 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 383 nsew signal input
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 384 nsew signal input
flabel metal3 s 59200 5992 60000 6112 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 385 nsew signal input
flabel metal3 s 59200 37000 60000 37120 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 386 nsew signal input
flabel metal3 s 59200 38632 60000 38752 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 387 nsew signal input
flabel metal3 s 59200 40264 60000 40384 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 388 nsew signal input
flabel metal3 s 59200 41896 60000 42016 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 389 nsew signal input
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 390 nsew signal input
flabel metal3 s 59200 45160 60000 45280 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 391 nsew signal input
flabel metal3 s 59200 46792 60000 46912 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 392 nsew signal input
flabel metal3 s 59200 48424 60000 48544 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 393 nsew signal input
flabel metal3 s 59200 50056 60000 50176 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 394 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 395 nsew signal input
flabel metal3 s 59200 7624 60000 7744 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 396 nsew signal input
flabel metal3 s 59200 53320 60000 53440 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 397 nsew signal input
flabel metal3 s 59200 54952 60000 55072 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 398 nsew signal input
flabel metal3 s 59200 9256 60000 9376 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 399 nsew signal input
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 400 nsew signal input
flabel metal3 s 59200 12520 60000 12640 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 401 nsew signal input
flabel metal3 s 59200 14152 60000 14272 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 402 nsew signal input
flabel metal3 s 59200 15784 60000 15904 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 403 nsew signal input
flabel metal3 s 59200 17416 60000 17536 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 404 nsew signal input
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 405 nsew signal input
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 wbs_cyc_i
port 406 nsew signal input
flabel metal3 s 59200 4904 60000 5024 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 407 nsew signal input
flabel metal3 s 59200 21224 60000 21344 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 408 nsew signal input
flabel metal3 s 59200 22856 60000 22976 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 409 nsew signal input
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 410 nsew signal input
flabel metal3 s 59200 26120 60000 26240 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 411 nsew signal input
flabel metal3 s 59200 27752 60000 27872 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 412 nsew signal input
flabel metal3 s 59200 29384 60000 29504 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 413 nsew signal input
flabel metal3 s 59200 31016 60000 31136 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 414 nsew signal input
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 415 nsew signal input
flabel metal3 s 59200 34280 60000 34400 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 416 nsew signal input
flabel metal3 s 59200 35912 60000 36032 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 417 nsew signal input
flabel metal3 s 59200 6536 60000 6656 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 418 nsew signal input
flabel metal3 s 59200 37544 60000 37664 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 419 nsew signal input
flabel metal3 s 59200 39176 60000 39296 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 420 nsew signal input
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 421 nsew signal input
flabel metal3 s 59200 42440 60000 42560 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 422 nsew signal input
flabel metal3 s 59200 44072 60000 44192 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 423 nsew signal input
flabel metal3 s 59200 45704 60000 45824 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 424 nsew signal input
flabel metal3 s 59200 47336 60000 47456 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 425 nsew signal input
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 426 nsew signal input
flabel metal3 s 59200 50600 60000 50720 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 427 nsew signal input
flabel metal3 s 59200 52232 60000 52352 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 428 nsew signal input
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 429 nsew signal input
flabel metal3 s 59200 53864 60000 53984 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 430 nsew signal input
flabel metal3 s 59200 55496 60000 55616 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 431 nsew signal input
flabel metal3 s 59200 9800 60000 9920 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 432 nsew signal input
flabel metal3 s 59200 11432 60000 11552 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 433 nsew signal input
flabel metal3 s 59200 13064 60000 13184 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 434 nsew signal input
flabel metal3 s 59200 14696 60000 14816 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 435 nsew signal input
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 436 nsew signal input
flabel metal3 s 59200 17960 60000 18080 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 437 nsew signal input
flabel metal3 s 59200 19592 60000 19712 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 438 nsew signal input
flabel metal3 s 59200 5448 60000 5568 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 439 nsew signal tristate
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 440 nsew signal tristate
flabel metal3 s 59200 23400 60000 23520 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 441 nsew signal tristate
flabel metal3 s 59200 25032 60000 25152 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 442 nsew signal tristate
flabel metal3 s 59200 26664 60000 26784 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 443 nsew signal tristate
flabel metal3 s 59200 28296 60000 28416 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 444 nsew signal tristate
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 445 nsew signal tristate
flabel metal3 s 59200 31560 60000 31680 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 446 nsew signal tristate
flabel metal3 s 59200 33192 60000 33312 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 447 nsew signal tristate
flabel metal3 s 59200 34824 60000 34944 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 448 nsew signal tristate
flabel metal3 s 59200 36456 60000 36576 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 449 nsew signal tristate
flabel metal3 s 59200 7080 60000 7200 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 450 nsew signal tristate
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 451 nsew signal tristate
flabel metal3 s 59200 39720 60000 39840 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 452 nsew signal tristate
flabel metal3 s 59200 41352 60000 41472 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 453 nsew signal tristate
flabel metal3 s 59200 42984 60000 43104 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 454 nsew signal tristate
flabel metal3 s 59200 44616 60000 44736 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 455 nsew signal tristate
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 456 nsew signal tristate
flabel metal3 s 59200 47880 60000 48000 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 457 nsew signal tristate
flabel metal3 s 59200 49512 60000 49632 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 458 nsew signal tristate
flabel metal3 s 59200 51144 60000 51264 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 459 nsew signal tristate
flabel metal3 s 59200 52776 60000 52896 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 460 nsew signal tristate
flabel metal3 s 59200 8712 60000 8832 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 461 nsew signal tristate
flabel metal3 s 59200 54408 60000 54528 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 462 nsew signal tristate
flabel metal3 s 59200 56040 60000 56160 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 463 nsew signal tristate
flabel metal3 s 59200 10344 60000 10464 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 464 nsew signal tristate
flabel metal3 s 59200 11976 60000 12096 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 465 nsew signal tristate
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 466 nsew signal tristate
flabel metal3 s 59200 15240 60000 15360 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 467 nsew signal tristate
flabel metal3 s 59200 16872 60000 16992 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 468 nsew signal tristate
flabel metal3 s 59200 18504 60000 18624 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 469 nsew signal tristate
flabel metal3 s 59200 20136 60000 20256 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 470 nsew signal tristate
flabel metal3 s 59200 3272 60000 3392 0 FreeSans 480 0 0 0 wbs_stb_i
port 471 nsew signal input
flabel metal3 s 59200 3816 60000 3936 0 FreeSans 480 0 0 0 wbs_we_i
port 472 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
<< end >>
