* NGSPICE file created from wrapped_6502.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt wrapped_6502 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_in[9] io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1 vssd1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1270_ _1648_/A _1624_/B vssd1 vssd1 vccd1 vccd1 _1653_/B sky130_fd_sc_hd__or2_2
X_1606_ _1803_/D _1626_/C vssd1 vssd1 vccd1 vccd1 _1606_/X sky130_fd_sc_hd__or2_1
X_0985_ _1041_/A _1024_/A vssd1 vssd1 vccd1 vccd1 _0985_/Y sky130_fd_sc_hd__nor2_1
X_1399_ _1752_/Q _1381_/C _1514_/B input7/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1399_/X
+ sky130_fd_sc_hd__a221o_1
X_1537_ _1542_/S _1547_/S _1536_/X _1792_/Q vssd1 vssd1 vccd1 vccd1 _1544_/S sky130_fd_sc_hd__o22a_1
X_1468_ _1723_/Q _1469_/B vssd1 vssd1 vccd1 vccd1 _1468_/X sky130_fd_sc_hd__or2_1
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1322_ _1586_/C _1323_/B vssd1 vssd1 vccd1 vccd1 _1626_/D sky130_fd_sc_hd__nor2_2
X_1253_ _1586_/C _1323_/B vssd1 vssd1 vccd1 vccd1 _1628_/B sky130_fd_sc_hd__and2_4
X_1184_ _1724_/Q _1173_/C _1206_/B _1749_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1184_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_12_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1807_/CLK sky130_fd_sc_hd__clkbuf_8
X_0968_ _0968_/A _1172_/B vssd1 vssd1 vccd1 vccd1 _1557_/S sky130_fd_sc_hd__or2_4
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0899_ _0968_/A _1084_/B vssd1 vssd1 vccd1 vccd1 _1554_/S sky130_fd_sc_hd__nor2_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1236_ _1719_/Q _1173_/D _1206_/X _1814_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1236_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1305_ _1628_/A _1624_/B vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__nand2_2
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1167_ _0952_/A _1166_/X _1165_/Y _1205_/A vssd1 vssd1 vccd1 vccd1 _1167_/X sky130_fd_sc_hd__o211a_1
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1098_ _1098_/A _1098_/B vssd1 vssd1 vccd1 vccd1 _1102_/B sky130_fd_sc_hd__nand2_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1021_ _1733_/Q _0950_/B _0974_/X input4/X vssd1 vssd1 vccd1 vccd1 _1028_/S sky130_fd_sc_hd__a22o_2
X_1785_ _1799_/CLK _1785_/D vssd1 vssd1 vccd1 vccd1 _1785_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1219_ input4/X _1156_/B _1205_/Y _1741_/Q _1218_/X vssd1 vssd1 vccd1 vccd1 _1220_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1570_ input2/X _1763_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1763_/D sky130_fd_sc_hd__mux2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1004_ _1004_/A _1011_/S vssd1 vssd1 vccd1 vccd1 _1004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1768_ _1769_/CLK _1768_/D vssd1 vssd1 vccd1 vccd1 _1768_/Q sky130_fd_sc_hd__dfxtp_1
X_1699_ _1769_/CLK _1699_/D _1693_/Y vssd1 vssd1 vccd1 vccd1 _1699_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput31 _0893_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_4
Xoutput20 _1401_/X vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_4
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1622_ _1802_/D _1613_/Y _1593_/C vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1484_ _1726_/Q _1489_/B _1495_/B vssd1 vssd1 vccd1 vccd1 _1484_/X sky130_fd_sc_hd__or3_1
X_1553_ _1759_/Q _1552_/X _1553_/S vssd1 vssd1 vccd1 vccd1 _1759_/D sky130_fd_sc_hd__mux2_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0984_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0984_/Y sky130_fd_sc_hd__inv_2
X_1605_ _1774_/Q _1604_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1774_/D sky130_fd_sc_hd__mux2_1
X_1536_ _1560_/A _1785_/Q _1549_/D _1536_/D vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__or4_1
X_1398_ _1735_/Q _1381_/X _1396_/X _1397_/X vssd1 vssd1 vccd1 vccd1 _1398_/X sky130_fd_sc_hd__o22a_1
X_1467_ _1703_/Q _1466_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1703_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1252_ _1256_/A _1252_/B vssd1 vssd1 vccd1 vccd1 _1323_/B sky130_fd_sc_hd__nand2_2
X_1321_ _1628_/A _1652_/B _1641_/D vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1183_ _1510_/B _1173_/C _1205_/A vssd1 vssd1 vccd1 vccd1 _1183_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0967_ _0968_/A _1172_/B vssd1 vssd1 vccd1 vccd1 _1542_/S sky130_fd_sc_hd__nor2_4
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0898_ _0968_/A _1083_/B vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__nor2_2
X_1519_ _1746_/Q _1383_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1746_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1235_ _1238_/A _1235_/B vssd1 vssd1 vccd1 vccd1 _1744_/D sky130_fd_sc_hd__and2_1
X_1304_ _1559_/A _1352_/B _1358_/C _1304_/D vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__or4_1
X_1166_ _1166_/A _1166_/B _1166_/C vssd1 vssd1 vccd1 vccd1 _1166_/X sky130_fd_sc_hd__and3_1
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1097_ _1125_/A _1048_/B _1048_/A vssd1 vssd1 vccd1 vccd1 _1098_/B sky130_fd_sc_hd__o21ai_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1829_/CLK sky130_fd_sc_hd__clkbuf_8
X_1020_ _1114_/A _1017_/Y _1019_/Y vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__o21a_2
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1784_ _1788_/CLK _1784_/D vssd1 vssd1 vccd1 vccd1 _1784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1218_ _1724_/Q _1173_/D _1206_/X _1810_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1218_/X
+ sky130_fd_sc_hd__a221o_1
X_1149_ _1759_/Q _1782_/Q vssd1 vssd1 vccd1 vccd1 _1755_/D sky130_fd_sc_hd__and2_1
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1003_ _1734_/Q _0950_/B _0974_/X input5/X vssd1 vssd1 vccd1 vccd1 _1011_/S sky130_fd_sc_hd__a22o_2
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1767_ _1767_/CLK _1767_/D vssd1 vssd1 vccd1 vccd1 _1767_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _1769_/CLK _1698_/D _1692_/Y vssd1 vssd1 vccd1 vccd1 _1698_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput21 _1404_/X vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_4
Xoutput32 _1436_/X vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1621_ _1780_/Q _1585_/Y _1650_/S vssd1 vssd1 vccd1 vccd1 _1780_/D sky130_fd_sc_hd__mux2_1
X_1552_ input4/X _1551_/X _1557_/S vssd1 vssd1 vccd1 vccd1 _1552_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1483_ _1489_/B _1495_/B _1726_/Q vssd1 vssd1 vccd1 vccd1 _1485_/B sky130_fd_sc_hd__o21a_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1819_ _1826_/CLK _1819_/D vssd1 vssd1 vccd1 vccd1 _1819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0983_ _1004_/A _1043_/A vssd1 vssd1 vccd1 vccd1 _0984_/A sky130_fd_sc_hd__and2_1
X_1604_ _1626_/D _1585_/Y _1598_/X _1603_/X vssd1 vssd1 vccd1 vccd1 _1604_/X sky130_fd_sc_hd__a211o_1
X_1535_ _1457_/A _1673_/B _1771_/Q vssd1 vssd1 vccd1 vccd1 _1536_/D sky130_fd_sc_hd__o21a_1
X_1397_ _1445_/B _1368_/Y _1381_/B _1726_/Q vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1466_ input2/X _1479_/S _1463_/X _1465_/Y vssd1 vssd1 vccd1 vccd1 _1466_/X sky130_fd_sc_hd__a22o_2
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1320_ _1641_/C _1320_/B _1320_/C vssd1 vssd1 vccd1 vccd1 _1320_/X sky130_fd_sc_hd__or3_1
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1251_ _1256_/A _1252_/B vssd1 vssd1 vccd1 vccd1 _1267_/B sky130_fd_sc_hd__and2_1
X_1182_ _1182_/A _1182_/B vssd1 vssd1 vccd1 vccd1 _1732_/D sky130_fd_sc_hd__xnor2_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0897_ _0897_/A _0897_/B _0927_/A _0909_/A vssd1 vssd1 vccd1 vccd1 _1083_/B sky130_fd_sc_hd__or4bb_4
X_0966_ input6/X _0950_/X _0965_/X vssd1 vssd1 vccd1 vccd1 _0966_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1518_ _1518_/A _1568_/B _1518_/C vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__and3_2
X_1449_ _1736_/Q _1372_/A _1424_/X _1761_/Q vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1303_ _1359_/A _1303_/B vssd1 vssd1 vccd1 vccd1 _1304_/D sky130_fd_sc_hd__nor2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1234_ _1234_/A _1234_/B vssd1 vssd1 vccd1 vccd1 _1235_/B sky130_fd_sc_hd__or2_1
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1165_ _1406_/C _1165_/B vssd1 vssd1 vccd1 vccd1 _1165_/Y sky130_fd_sc_hd__nand2_1
X_1096_ _1103_/A _1095_/B _1062_/X vssd1 vssd1 vccd1 vccd1 _1102_/A sky130_fd_sc_hd__a21oi_4
X_0949_ _0952_/A _1166_/B vssd1 vssd1 vccd1 vccd1 _0950_/B sky130_fd_sc_hd__nor2_8
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1783_ _1803_/CLK _1783_/D vssd1 vssd1 vccd1 vccd1 _1783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1217_ _1220_/A _1220_/B vssd1 vssd1 vccd1 vccd1 _1740_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1148_ _1145_/X _1146_/Y _1147_/X vssd1 vssd1 vccd1 vccd1 _1718_/D sky130_fd_sc_hd__a21o_1
X_1079_ _1077_/Y _1079_/B vssd1 vssd1 vccd1 vccd1 _1150_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1002_ _1114_/A _0999_/Y _1001_/Y vssd1 vssd1 vccd1 vccd1 _1006_/B sky130_fd_sc_hd__o21a_2
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1697_ _1769_/CLK _1697_/D _1691_/Y vssd1 vssd1 vccd1 vccd1 _1697_/Q sky130_fd_sc_hd__dfrtp_2
X_1766_ _1767_/CLK _1766_/D vssd1 vssd1 vccd1 vccd1 _1766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1826_/CLK sky130_fd_sc_hd__clkbuf_8
Xoutput22 _1408_/X vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_4
Xoutput33 _1439_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_4
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1620_ _1650_/S _1589_/B _1613_/Y _1619_/X vssd1 vssd1 vccd1 vccd1 _1779_/D sky130_fd_sc_hd__a31o_1
X_1551_ _0831_/Y _1724_/Q _1560_/A vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__mux2_1
X_1482_ _1718_/Q _1482_/B vssd1 vssd1 vccd1 vccd1 _1495_/B sky130_fd_sc_hd__nor2_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1818_ _1826_/CLK _1818_/D vssd1 vssd1 vccd1 vccd1 _1818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1749_ _1808_/CLK _1749_/D vssd1 vssd1 vccd1 vccd1 _1749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ _1004_/A _1043_/A vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__or2_2
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1603_ _1580_/Y _1593_/C _1602_/B vssd1 vssd1 vccd1 vccd1 _1603_/X sky130_fd_sc_hd__o21a_1
X_1534_ _1754_/Q _1533_/X _1534_/S vssd1 vssd1 vccd1 vccd1 _1754_/D sky130_fd_sc_hd__mux2_1
X_1465_ _1479_/S _1465_/B vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__nor2_1
X_1396_ _1751_/Q _1381_/C _1514_/B input6/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1396_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1250_ _1256_/A _1250_/B vssd1 vssd1 vccd1 vccd1 _1586_/C sky130_fd_sc_hd__and2_4
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1181_ _1182_/B _1181_/B _1175_/B vssd1 vssd1 vccd1 vccd1 _1187_/A sky130_fd_sc_hd__or3b_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0896_ _0952_/A _1152_/A vssd1 vssd1 vccd1 vccd1 _0896_/X sky130_fd_sc_hd__or2_1
X_0965_ _1812_/Q _1406_/C _0957_/X _1726_/Q _0964_/Y vssd1 vssd1 vccd1 vccd1 _0965_/X
+ sky130_fd_sc_hd__a221o_2
X_1517_ _1517_/A _1517_/B _1517_/C _1163_/Y vssd1 vssd1 vccd1 vccd1 _1518_/C sky130_fd_sc_hd__or4b_1
X_1448_ _1448_/A _1448_/B _1448_/C vssd1 vssd1 vccd1 vccd1 _1448_/X sky130_fd_sc_hd__or3_2
X_1379_ _1721_/Q _1381_/B _1514_/B input1/X vssd1 vssd1 vccd1 vccd1 _1379_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1233_ _1234_/A _1234_/B vssd1 vssd1 vccd1 vccd1 _1238_/A sky130_fd_sc_hd__nand2_1
X_1302_ _1641_/C _1580_/A _1653_/B _1320_/B vssd1 vssd1 vccd1 vccd1 _1303_/B sky130_fd_sc_hd__or4_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1164_ _1756_/Q _1718_/Q vssd1 vssd1 vccd1 vccd1 _1165_/B sky130_fd_sc_hd__xnor2_1
X_1095_ _1062_/X _1095_/B vssd1 vssd1 vccd1 vccd1 _1103_/B sky130_fd_sc_hd__nand2b_2
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0948_ _1114_/A _0948_/B vssd1 vssd1 vccd1 vccd1 _0948_/Y sky130_fd_sc_hd__nor2_1
X_0879_ _0927_/A _0909_/A _0897_/B _0897_/A vssd1 vssd1 vccd1 vccd1 _1084_/B sky130_fd_sc_hd__or4b_4
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1782_ _1799_/CLK _1782_/D vssd1 vssd1 vccd1 vccd1 _1782_/Q sky130_fd_sc_hd__dfxtp_1
X_1216_ input3/X _1156_/B _1205_/Y _1740_/Q _1215_/X vssd1 vssd1 vccd1 vccd1 _1220_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1147_ _1727_/D _1726_/D _1142_/A _1105_/X _1142_/B vssd1 vssd1 vccd1 vccd1 _1147_/X
+ sky130_fd_sc_hd__o2111a_1
X_1078_ _1125_/A _1076_/X _1075_/X _1063_/X vssd1 vssd1 vccd1 vccd1 _1079_/B sky130_fd_sc_hd__o211ai_4
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _1725_/Q _0957_/X _1000_/X vssd1 vssd1 vccd1 vccd1 _1001_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1765_ _1767_/CLK _1765_/D vssd1 vssd1 vccd1 vccd1 _1765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1696_ _1769_/CLK _1696_/D _0836_/Y vssd1 vssd1 vccd1 vccd1 _1696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput12 _0893_/A vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_4
Xoutput23 _1411_/X vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_4
Xoutput34 _1444_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_4
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1550_ _1566_/A2 _1542_/S _1549_/X vssd1 vssd1 vccd1 vccd1 _1553_/S sky130_fd_sc_hd__o21a_1
X_1481_ _1718_/Q _1784_/Q _1755_/Q vssd1 vssd1 vccd1 vccd1 _1489_/B sky130_fd_sc_hd__and3_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1748_ _1808_/CLK _1748_/D vssd1 vssd1 vccd1 vccd1 _1748_/Q sky130_fd_sc_hd__dfxtp_2
X_1817_ _1825_/CLK _1817_/D vssd1 vssd1 vccd1 vccd1 _1817_/Q sky130_fd_sc_hd__dfxtp_1
X_1679_ _1820_/Q _1486_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1820_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0981_ _1789_/Q _1513_/C _0977_/Y vssd1 vssd1 vccd1 vccd1 _1043_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1602_ _1650_/S _1602_/B vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__and2_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1395_ _1734_/Q _1381_/X _1393_/X _1394_/X vssd1 vssd1 vccd1 vccd1 _1395_/X sky130_fd_sc_hd__o22a_1
X_1533_ input1/X _1532_/X _1557_/S vssd1 vssd1 vccd1 vccd1 _1533_/X sky130_fd_sc_hd__mux2_1
X_1464_ _1469_/B _1475_/B _1722_/Q vssd1 vssd1 vccd1 vccd1 _1465_/B sky130_fd_sc_hd__o21a_1
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1180_ _1748_/Q _1206_/B _1178_/X _1179_/X vssd1 vssd1 vccd1 vccd1 _1182_/B sky130_fd_sc_hd__a211oi_4
X_0964_ _1114_/A _1445_/B vssd1 vssd1 vccd1 vccd1 _0964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1516_ _1516_/A _1516_/B _1516_/C _1516_/D vssd1 vssd1 vccd1 vccd1 _1517_/C sky130_fd_sc_hd__or4_1
X_0895_ _1083_/A _1152_/A vssd1 vssd1 vccd1 vccd1 _1105_/B sky130_fd_sc_hd__nor2_2
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1378_ _1298_/A _0925_/B _0887_/D vssd1 vssd1 vccd1 vccd1 _1378_/Y sky130_fd_sc_hd__o21bai_4
X_1447_ _1735_/Q _1372_/A _1369_/B _1743_/Q _1424_/X vssd1 vssd1 vccd1 vccd1 _1448_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout80 _1700_/Q vssd1 vssd1 vccd1 vccd1 _0914_/A sky130_fd_sc_hd__buf_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1232_ input7/X _1156_/B _1205_/Y _1744_/Q _1231_/X vssd1 vssd1 vccd1 vccd1 _1234_/B
+ sky130_fd_sc_hd__a221o_1
X_1301_ _1614_/B _1641_/B vssd1 vssd1 vccd1 vccd1 _1320_/B sky130_fd_sc_hd__or2_2
X_1163_ _1163_/A _1336_/A vssd1 vssd1 vccd1 vccd1 _1163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1094_ _0994_/B _1061_/X _1060_/X _1049_/Y vssd1 vssd1 vccd1 vccd1 _1095_/B sky130_fd_sc_hd__a211o_2
X_0947_ _1829_/Q _1682_/A _1500_/A _1716_/Q _0944_/X vssd1 vssd1 vccd1 vccd1 _0948_/B
+ sky130_fd_sc_hd__a221oi_4
X_0878_ _0878_/A _1510_/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__or2_4
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ _1799_/CLK _1781_/D vssd1 vssd1 vccd1 vccd1 _1781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1215_ _1723_/Q _1173_/D _1206_/X _1809_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1215_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ _1063_/A _1072_/X _1139_/A _1142_/A vssd1 vssd1 vccd1 vccd1 _1146_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ _1063_/X _1075_/X _1076_/X vssd1 vssd1 vccd1 vccd1 _1077_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1000_ input5/X _0950_/X _1406_/C _1811_/Q vssd1 vssd1 vccd1 vccd1 _1000_/X sky130_fd_sc_hd__a22o_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1764_ _1767_/CLK _1764_/D vssd1 vssd1 vccd1 vccd1 _1764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1695_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1129_ _1141_/B _1129_/B vssd1 vssd1 vccd1 vccd1 _1727_/D sky130_fd_sc_hd__and2_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput13 _1429_/X vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_4
Xoutput24 _1432_/X vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_4
Xoutput35 _1448_/X vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_4
XFILLER_8_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1706_/Q _1479_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1706_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1816_ _1826_/CLK _1816_/D vssd1 vssd1 vccd1 vccd1 _1816_/Q sky130_fd_sc_hd__dfxtp_1
X_1678_ _1819_/Q _1479_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1819_/D sky130_fd_sc_hd__mux2_1
X_1747_ _1829_/CLK _1747_/D vssd1 vssd1 vccd1 vccd1 _1747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0980_ _1789_/Q _1513_/C _0977_/Y vssd1 vssd1 vccd1 vccd1 _1024_/A sky130_fd_sc_hd__a21oi_4
X_1601_ _1626_/B _1599_/X _1600_/X vssd1 vssd1 vccd1 vccd1 _1773_/D sky130_fd_sc_hd__a21o_1
X_1532_ _1531_/X _1718_/Q _1532_/S vssd1 vssd1 vccd1 vccd1 _1532_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1463_ _1722_/Q _1469_/B _1475_/B vssd1 vssd1 vccd1 vccd1 _1463_/X sky130_fd_sc_hd__or3_1
X_1394_ _0999_/Y _1368_/Y _1381_/B _1725_/Q vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0894_ _0894_/A _0953_/C vssd1 vssd1 vccd1 vccd1 _1152_/A sky130_fd_sc_hd__or2_4
X_0963_ _1828_/Q _1682_/A _1500_/A _1715_/Q _0962_/X vssd1 vssd1 vccd1 vccd1 _1445_/B
+ sky130_fd_sc_hd__a221oi_4
X_1515_ _1515_/A _1515_/B _1515_/C vssd1 vssd1 vccd1 vccd1 _1516_/D sky130_fd_sc_hd__or3_1
X_1377_ _1510_/A _1406_/B _1377_/C vssd1 vssd1 vccd1 vccd1 _1381_/C sky130_fd_sc_hd__or3_4
X_1446_ _1369_/A _0876_/Y _1726_/Q vssd1 vssd1 vccd1 vccd1 _1448_/B sky130_fd_sc_hd__o21a_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout81 _1700_/Q vssd1 vssd1 vccd1 vccd1 _0933_/A sky130_fd_sc_hd__buf_4
Xfanout70 _1579_/A vssd1 vssd1 vccd1 vccd1 _1256_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1231_ _1727_/Q _1173_/D _1206_/X _1813_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1231_/X
+ sky130_fd_sc_hd__a221o_1
X_1162_ _1162_/A _1162_/B _1162_/C vssd1 vssd1 vccd1 vccd1 _1166_/C sky130_fd_sc_hd__or3_1
X_1300_ _1300_/A vssd1 vssd1 vccd1 vccd1 _1300_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1093_ _1079_/B _1092_/A _1092_/B _1077_/Y vssd1 vssd1 vccd1 vccd1 _1103_/A sky130_fd_sc_hd__a31o_4
X_0877_ _0878_/A _1510_/A vssd1 vssd1 vccd1 vccd1 _1435_/A sky130_fd_sc_hd__nor2_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0946_ _1050_/S _1673_/B vssd1 vssd1 vccd1 vccd1 _1500_/A sky130_fd_sc_hd__nor2_8
X_1429_ _1435_/A _1426_/X _1427_/X _1428_/Y vssd1 vssd1 vccd1 vccd1 _1429_/X sky130_fd_sc_hd__o31a_2
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1780_ _1799_/CLK _1780_/D vssd1 vssd1 vccd1 vccd1 _1780_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1214_ _1220_/A _1214_/B vssd1 vssd1 vccd1 vccd1 _1739_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1145_ _1139_/A _1142_/A _1063_/A _1072_/X vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__a211o_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1076_ _0992_/A _1010_/A _1076_/S vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__mux2_2
X_0929_ _0914_/A _0869_/B _0912_/B _1373_/A vssd1 vssd1 vccd1 vccd1 _0929_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1694_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__inv_2
X_1763_ _1767_/CLK _1763_/D vssd1 vssd1 vccd1 vccd1 _1763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1128_ _1128_/A _1144_/A _1128_/C vssd1 vssd1 vccd1 vccd1 _1129_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1059_ _1004_/A _1061_/S _1063_/B vssd1 vssd1 vccd1 vccd1 _1059_/X sky130_fd_sc_hd__a21bo_1
Xoutput25 _1413_/X vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput36 _1451_/X vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_4
Xoutput14 _1383_/X vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_4
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1815_ _1830_/CLK _1815_/D vssd1 vssd1 vccd1 vccd1 _1815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1677_ _1818_/Q _1477_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1818_/D sky130_fd_sc_hd__mux2_1
X_1746_ _1829_/CLK _1746_/D vssd1 vssd1 vccd1 vccd1 _1746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1600_ _1773_/Q _1549_/D _1292_/B vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__a21o_1
X_1531_ _0837_/Y _1721_/Q _1560_/A vssd1 vssd1 vccd1 vccd1 _1531_/X sky130_fd_sc_hd__mux2_1
X_1462_ _1720_/Q _1482_/B vssd1 vssd1 vccd1 vccd1 _1475_/B sky130_fd_sc_hd__nor2_2
X_1393_ _1750_/Q _1381_/C _1514_/B input5/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1393_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1729_ _1797_/CLK _1729_/D vssd1 vssd1 vccd1 vccd1 _1729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0893_ _0893_/A vssd1 vssd1 vccd1 vccd1 _0893_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0962_ _1820_/Q _1457_/A _1673_/B _0961_/X vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1514_ _1514_/A _1514_/B _1547_/S vssd1 vssd1 vccd1 vccd1 _1516_/C sky130_fd_sc_hd__or3_1
X_1445_ _1445_/A _1445_/B vssd1 vssd1 vccd1 vccd1 _1448_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1376_ _1162_/B _0890_/Y _1173_/D _1513_/B vssd1 vssd1 vccd1 vccd1 _1377_/C sky130_fd_sc_hd__a211o_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout60 _0927_/X vssd1 vssd1 vccd1 vccd1 _1577_/B sky130_fd_sc_hd__buf_6
Xfanout82 _0897_/B vssd1 vssd1 vccd1 vccd1 _1162_/C sky130_fd_sc_hd__buf_4
Xfanout71 _0838_/Y vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__buf_12
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1230_ _1234_/A _1230_/B vssd1 vssd1 vccd1 vccd1 _1743_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1161_ _1730_/Q _1158_/Y _1160_/X vssd1 vssd1 vccd1 vccd1 _1170_/A sky130_fd_sc_hd__a21oi_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1092_ _1092_/A _1092_/B vssd1 vssd1 vccd1 vccd1 _1150_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0876_ _0968_/A _0912_/B vssd1 vssd1 vccd1 vccd1 _0876_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0945_ _1673_/A _1673_/B vssd1 vssd1 vccd1 vccd1 _1682_/A sky130_fd_sc_hd__nor2_8
X_1428_ _1435_/A _1428_/B vssd1 vssd1 vccd1 vccd1 _1428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1359_ _1359_/A _1359_/B vssd1 vssd1 vccd1 vccd1 _1360_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ _1212_/A _1212_/B _1212_/C vssd1 vssd1 vccd1 vccd1 _1214_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1726_/D sky130_fd_sc_hd__and2_1
X_1075_ _1076_/S _1072_/X _1073_/Y _1074_/X _1091_/A vssd1 vssd1 vccd1 vccd1 _1075_/X
+ sky130_fd_sc_hd__a221o_4
X_0859_ _1172_/A _0970_/A vssd1 vssd1 vccd1 vccd1 _1513_/A sky130_fd_sc_hd__nor2_2
X_0928_ _0928_/A _1366_/A _1286_/A _1510_/B vssd1 vssd1 vccd1 vccd1 _0941_/C sky130_fd_sc_hd__nor4_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1693_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1693_/Y sky130_fd_sc_hd__inv_2
X_1762_ _1767_/CLK _1762_/D vssd1 vssd1 vccd1 vccd1 _1762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1127_ _1128_/A _1144_/A _1128_/C vssd1 vssd1 vccd1 vccd1 _1141_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1058_ _1004_/A _1024_/A _1058_/S vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput26 _1415_/X vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_4
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput15 _1386_/X vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput37 _1454_/X vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ _1806_/CLK _1745_/D vssd1 vssd1 vccd1 vccd1 _1745_/Q sky130_fd_sc_hd__dfxtp_2
X_1814_ _1814_/CLK _1814_/D vssd1 vssd1 vccd1 vccd1 _1814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _1817_/Q _1472_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1817_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1530_ _1532_/S _1528_/X _1529_/X _1542_/S vssd1 vssd1 vccd1 vccd1 _1534_/S sky130_fd_sc_hd__o22a_1
X_1392_ _1733_/Q _1381_/X _1390_/X _1391_/X vssd1 vssd1 vccd1 vccd1 _1392_/X sky130_fd_sc_hd__o22a_1
X_1461_ _1784_/Q _1755_/Q vssd1 vssd1 vccd1 vccd1 _1482_/B sky130_fd_sc_hd__nand2b_2
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1728_ _1797_/CLK _1728_/D vssd1 vssd1 vccd1 vccd1 _1728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ _1798_/Q _1648_/B _1644_/Y _1652_/X vssd1 vssd1 vccd1 vccd1 _1798_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0961_ _1707_/Q _1673_/A vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__or2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0892_ _1445_/A _0892_/B vssd1 vssd1 vccd1 vccd1 _0893_/A sky130_fd_sc_hd__nor2_2
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1375_ _1375_/A _1375_/B _1375_/C _1375_/D vssd1 vssd1 vccd1 vccd1 _1381_/B sky130_fd_sc_hd__or4_4
X_1513_ _1513_/A _1513_/B _1513_/C _1513_/D vssd1 vssd1 vccd1 vccd1 _1516_/B sky130_fd_sc_hd__or4_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1444_ _1445_/A _0999_/Y _1443_/X vssd1 vssd1 vccd1 vccd1 _1444_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout83 _1699_/Q vssd1 vssd1 vccd1 vccd1 _0897_/B sky130_fd_sc_hd__buf_4
Xfanout72 _1242_/X vssd1 vssd1 vccd1 vccd1 _1652_/B sky130_fd_sc_hd__buf_4
Xfanout50 _1344_/B vssd1 vssd1 vccd1 vccd1 _1630_/C sky130_fd_sc_hd__buf_4
Xfanout61 _1566_/A2 vssd1 vssd1 vccd1 vccd1 _1650_/S sky130_fd_sc_hd__buf_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _1721_/Q _1173_/C _1206_/B _1746_/Q vssd1 vssd1 vccd1 vccd1 _1160_/X sky130_fd_sc_hd__a22o_1
X_1091_ _1091_/A _1124_/A vssd1 vssd1 vccd1 vccd1 _1092_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0944_ _1821_/Q _1457_/A _1673_/B _0943_/X vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0875_ _0909_/A _0897_/A _0897_/B _0927_/A vssd1 vssd1 vccd1 vccd1 _0912_/B sky130_fd_sc_hd__nand4b_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1358_ _1358_/A _1358_/B _1358_/C _1358_/D vssd1 vssd1 vccd1 vccd1 _1360_/C sky130_fd_sc_hd__or4_1
X_1427_ _1730_/Q _1372_/A _1425_/Y _1721_/Q vssd1 vssd1 vccd1 vccd1 _1427_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1289_ _0869_/B _0970_/B _0918_/Y _0968_/A vssd1 vssd1 vccd1 vccd1 _1290_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ _1212_/A _1212_/B _1212_/C vssd1 vssd1 vccd1 vccd1 _1220_/A sky130_fd_sc_hd__and3_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1143_ _1128_/A _1109_/Y _1240_/A _1014_/A vssd1 vssd1 vccd1 vccd1 _1144_/B sky130_fd_sc_hd__a211o_1
X_1074_ _1024_/A _1076_/S _1072_/X _0984_/A vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__a211o_1
X_0927_ _0927_/A _1162_/A _0952_/A _0953_/C vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__or4_1
X_0858_ _1162_/A _1162_/B _1162_/C _0917_/A vssd1 vssd1 vccd1 vccd1 _0970_/A sky130_fd_sc_hd__or4bb_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1761_ _1803_/CLK _1761_/D vssd1 vssd1 vccd1 vccd1 _1761_/Q sky130_fd_sc_hd__dfxtp_1
X_1830_ _1830_/CLK _1830_/D vssd1 vssd1 vccd1 vccd1 _1830_/Q sky130_fd_sc_hd__dfxtp_1
X_1692_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1692_/Y sky130_fd_sc_hd__inv_2
X_1126_ _1124_/B _1125_/X _1141_/A vssd1 vssd1 vccd1 vccd1 _1128_/C sky130_fd_sc_hd__a21bo_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1057_ _1063_/B _1061_/S vssd1 vssd1 vccd1 vccd1 _1058_/S sky130_fd_sc_hd__and2b_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput27 _1417_/X vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_4
Xoutput16 _1389_/X vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1814_/CLK _1744_/D vssd1 vssd1 vccd1 vccd1 _1744_/Q sky130_fd_sc_hd__dfxtp_2
X_1813_ _1814_/CLK _1813_/D vssd1 vssd1 vccd1 vccd1 _1813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1675_ _1816_/Q _1466_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1816_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1109_ _1125_/A _0995_/X _0996_/B vssd1 vssd1 vccd1 vccd1 _1109_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1460_ _1784_/Q _1755_/Q _1720_/Q vssd1 vssd1 vccd1 vccd1 _1469_/B sky130_fd_sc_hd__and3_1
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1391_ _1017_/Y _1368_/Y _1381_/B _1724_/Q vssd1 vssd1 vccd1 vccd1 _1391_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1658_ _1797_/Q _1648_/B _1602_/X _1655_/X vssd1 vssd1 vccd1 vccd1 _1797_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1727_ _1788_/CLK _1727_/D vssd1 vssd1 vccd1 vccd1 _1727_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1589_/A _1589_/B vssd1 vssd1 vccd1 vccd1 _1589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ _1063_/A _0960_/B vssd1 vssd1 vccd1 vccd1 _0960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0891_ _1284_/B _0890_/Y _1778_/Q vssd1 vssd1 vccd1 vccd1 _0892_/B sky130_fd_sc_hd__o21a_1
X_1512_ _1512_/A _1512_/B _1512_/C _1512_/D vssd1 vssd1 vccd1 vccd1 _1513_/D sky130_fd_sc_hd__or4_1
X_1374_ _1374_/A _1374_/B _1406_/C _1345_/A vssd1 vssd1 vccd1 vccd1 _1375_/D sky130_fd_sc_hd__or4b_1
X_1443_ _1806_/Q input9/X _0860_/X _1442_/Y vssd1 vssd1 vccd1 vccd1 _1443_/X sky130_fd_sc_hd__o31a_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout73 _0862_/Y vssd1 vssd1 vccd1 vccd1 _0968_/A sky130_fd_sc_hd__buf_6
Xfanout62 _1566_/A2 vssd1 vssd1 vccd1 vccd1 _1626_/B sky130_fd_sc_hd__clkbuf_8
Xfanout51 _0870_/X vssd1 vssd1 vccd1 vccd1 _1369_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout40 _1380_/Y vssd1 vssd1 vccd1 vccd1 _1410_/B1 sky130_fd_sc_hd__buf_4
Xfanout84 _0897_/A vssd1 vssd1 vccd1 vccd1 _1162_/B sky130_fd_sc_hd__buf_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1090_ _1090_/A _1090_/B vssd1 vssd1 vccd1 vccd1 _1092_/A sky130_fd_sc_hd__nand2_2
X_0874_ _1162_/A _0932_/B _0953_/C vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__or3_1
X_0943_ _1708_/Q _1673_/A vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__or2_1
XFILLER_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1288_ _1344_/A _1630_/C _1308_/A vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__or3_1
X_1357_ _1357_/A _1456_/A vssd1 vssd1 vccd1 vccd1 _1358_/D sky130_fd_sc_hd__nand2_1
X_1426_ _1738_/Q _1369_/B _1424_/X _1754_/Q vssd1 vssd1 vccd1 vccd1 _1426_/X sky130_fd_sc_hd__a22o_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1211_ input2/X _1156_/B _1205_/Y _1739_/Q _1210_/X vssd1 vssd1 vccd1 vccd1 _1212_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1142_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1719_/D sky130_fd_sc_hd__and2_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1073_ _1076_/S _1072_/X _1004_/A vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__o21ai_1
X_0926_ _0926_/A _0926_/B _0926_/C vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__and3_2
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0857_ _1298_/A _1166_/A _0973_/C vssd1 vssd1 vccd1 vccd1 _0957_/A sky130_fd_sc_hd__o21ai_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1409_ input2/X _1375_/A _1406_/X _1808_/Q vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1691_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1691_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1760_ _1804_/CLK _1760_/D vssd1 vssd1 vccd1 vccd1 _1760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1125_ _1125_/A _1125_/B vssd1 vssd1 vccd1 vccd1 _1125_/X sky130_fd_sc_hd__or2_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1056_ _1731_/Q _0950_/B _0974_/X input2/X vssd1 vssd1 vccd1 vccd1 _1061_/S sky130_fd_sc_hd__a22o_2
Xoutput28 _1419_/X vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_4
X_0909_ _0909_/A _1298_/A _0953_/C vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__nor3_2
Xoutput17 _1392_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_4
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1743_ _1814_/CLK _1743_/D vssd1 vssd1 vccd1 vccd1 _1743_/Q sky130_fd_sc_hd__dfxtp_2
X_1812_ _1814_/CLK _1812_/D vssd1 vssd1 vccd1 vccd1 _1812_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1674_ _1815_/Q _1458_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1815_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1108_ _1239_/B _1239_/C _1239_/A vssd1 vssd1 vccd1 vccd1 _1240_/A sky130_fd_sc_hd__a21oi_4
X_1039_ _1114_/A _1435_/B _1038_/Y vssd1 vssd1 vccd1 vccd1 _1049_/B sky130_fd_sc_hd__o21a_2
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1390_ _1749_/Q _1381_/C _1514_/B input4/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1390_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1588_ _1802_/D _1588_/B vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__nand2_2
X_1657_ _1796_/Q _1648_/B _1602_/X _1652_/X vssd1 vssd1 vccd1 vccd1 _1796_/D sky130_fd_sc_hd__a22o_1
X_1726_ _1788_/CLK _1726_/D vssd1 vssd1 vccd1 vccd1 _1726_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0890_ _1373_/A _0904_/B vssd1 vssd1 vccd1 vccd1 _0890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1511_ _1511_/A _1511_/B vssd1 vssd1 vccd1 vccd1 _1517_/B sky130_fd_sc_hd__nand2_1
X_1442_ _1800_/Q _1369_/A _1441_/X vssd1 vssd1 vccd1 vccd1 _1442_/Y sky130_fd_sc_hd__a21oi_1
X_1373_ _1373_/A _1373_/B vssd1 vssd1 vccd1 vccd1 _1375_/C sky130_fd_sc_hd__nor2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1709_ _1830_/CLK _1709_/D vssd1 vssd1 vccd1 vccd1 _1709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout85 _1698_/Q vssd1 vssd1 vccd1 vccd1 _0897_/A sky130_fd_sc_hd__buf_4
Xfanout74 _0862_/Y vssd1 vssd1 vccd1 vccd1 _0932_/B sky130_fd_sc_hd__buf_6
Xfanout63 _1510_/B vssd1 vssd1 vccd1 vccd1 _1566_/A2 sky130_fd_sc_hd__buf_4
Xfanout52 _1586_/A vssd1 vssd1 vccd1 vccd1 _1655_/A sky130_fd_sc_hd__buf_6
Xfanout41 _1380_/Y vssd1 vssd1 vccd1 vccd1 _1423_/A2 sky130_fd_sc_hd__buf_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0873_ _1698_/Q _1162_/C vssd1 vssd1 vccd1 vccd1 _0953_/C sky130_fd_sc_hd__nand2_4
X_0942_ _1774_/Q _1510_/B _0941_/X _1512_/C _1286_/A vssd1 vssd1 vccd1 vccd1 _1052_/S
+ sky130_fd_sc_hd__a2111o_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1425_ _1800_/Q _1518_/A _1510_/A vssd1 vssd1 vccd1 vccd1 _1425_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1287_ _1366_/B _1339_/C _1287_/C vssd1 vssd1 vccd1 vccd1 _1290_/B sky130_fd_sc_hd__or3_1
X_1356_ _1485_/A _1356_/B _1559_/A vssd1 vssd1 vccd1 vccd1 _1456_/A sky130_fd_sc_hd__nor3_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1210_ _1722_/Q _1173_/D _1206_/X _1808_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1210_/X
+ sky130_fd_sc_hd__a221o_1
X_1141_ _1141_/A _1141_/B _1141_/C vssd1 vssd1 vccd1 vccd1 _1142_/B sky130_fd_sc_hd__nand3_1
X_1072_ _1114_/A _1428_/B _1071_/Y vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__o21a_4
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0856_ _0952_/A _1298_/B vssd1 vssd1 vccd1 vccd1 _0973_/C sky130_fd_sc_hd__or2_4
X_0925_ _1083_/A _0925_/B vssd1 vssd1 vccd1 vccd1 _1286_/A sky130_fd_sc_hd__nor2_4
X_1408_ _1738_/Q _1410_/B1 _1405_/X _1407_/X vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1339_ _1351_/A _1339_/B _1339_/C _1288_/X vssd1 vssd1 vccd1 vccd1 _1340_/D sky130_fd_sc_hd__or4b_1
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _1830_/Q _1498_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1830_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1124_ _1124_/A _1124_/B _1125_/B vssd1 vssd1 vccd1 vccd1 _1141_/A sky130_fd_sc_hd__or3_2
X_1055_ _0924_/Y _1052_/X _1054_/X vssd1 vssd1 vccd1 vccd1 _1063_/B sky130_fd_sc_hd__a21oi_2
X_0839_ input8/X _1769_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1648_/A sky130_fd_sc_hd__mux2_8
Xoutput29 _1421_/X vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_4
X_0908_ _1485_/A _1369_/C vssd1 vssd1 vccd1 vccd1 _0941_/B sky130_fd_sc_hd__nor2_2
Xoutput18 _1395_/X vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_4
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1811_ _1814_/CLK _1811_/D vssd1 vssd1 vccd1 vccd1 _1811_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1742_ _1814_/CLK _1742_/D vssd1 vssd1 vccd1 vccd1 _1742_/Q sky130_fd_sc_hd__dfxtp_2
X_1673_ _1673_/A _1673_/B _1682_/B vssd1 vssd1 vccd1 vccd1 _1681_/S sky130_fd_sc_hd__and3_4
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1107_ _1239_/B _1239_/C vssd1 vssd1 vccd1 vccd1 _1720_/D sky130_fd_sc_hd__nand2_1
X_1038_ _1723_/Q _0957_/X _1037_/X vssd1 vssd1 vccd1 vccd1 _1038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1725_ _1825_/CLK _1725_/D vssd1 vssd1 vccd1 vccd1 _1725_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1587_ _1804_/D _1624_/B _1652_/B vssd1 vssd1 vccd1 vccd1 _1588_/B sky130_fd_sc_hd__and3_1
X_1656_ _1795_/Q _1653_/A _1653_/Y _1655_/X vssd1 vssd1 vccd1 vccd1 _1795_/D sky130_fd_sc_hd__a22o_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1441_ _1734_/Q _1372_/A _1369_/B _1742_/Q _1440_/X vssd1 vssd1 vccd1 vccd1 _1441_/X
+ sky130_fd_sc_hd__a221o_1
X_1510_ _1510_/A _1510_/B vssd1 vssd1 vccd1 vccd1 _1547_/S sky130_fd_sc_hd__or2_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1372_ _1372_/A _1372_/B _1372_/C vssd1 vssd1 vccd1 vccd1 _1375_/B sky130_fd_sc_hd__or3_1
XFILLER_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1708_ _1826_/CLK _1708_/D vssd1 vssd1 vccd1 vccd1 _1708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1639_ _1655_/A _1613_/Y _1630_/X vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__a21o_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout75 _1083_/A vssd1 vssd1 vccd1 vccd1 _0952_/A sky130_fd_sc_hd__buf_8
Xfanout86 _1697_/Q vssd1 vssd1 vccd1 vccd1 _0927_/A sky130_fd_sc_hd__clkbuf_8
Xfanout53 _0952_/Y vssd1 vssd1 vccd1 vccd1 _1406_/C sky130_fd_sc_hd__buf_4
Xfanout64 _0926_/X vssd1 vssd1 vccd1 vccd1 _1510_/B sky130_fd_sc_hd__buf_12
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout42 _1041_/A vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0941_ _1776_/Q _0941_/B _0941_/C _0941_/D vssd1 vssd1 vccd1 vccd1 _0941_/X sky130_fd_sc_hd__and4_1
X_0872_ _0897_/A _0897_/B vssd1 vssd1 vccd1 vccd1 _0926_/C sky130_fd_sc_hd__and2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1355_ _1298_/A _1354_/X _0918_/Y _0933_/A vssd1 vssd1 vccd1 vccd1 _1360_/B sky130_fd_sc_hd__a2bb2o_1
X_1424_ _1800_/Q _1369_/A _0957_/B vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__a21o_2
X_1286_ _1286_/A _1286_/B _1358_/A _1339_/B vssd1 vssd1 vccd1 vccd1 _1287_/C sky130_fd_sc_hd__or4_1
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1071_ _1721_/Q _0957_/X _1070_/X vssd1 vssd1 vccd1 vccd1 _1071_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _1141_/A _1141_/B _1141_/C vssd1 vssd1 vccd1 vccd1 _1142_/A sky130_fd_sc_hd__a21o_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0924_ _1114_/A vssd1 vssd1 vccd1 vccd1 _0924_/Y sky130_fd_sc_hd__inv_2
X_0855_ _1162_/B _0868_/A _0894_/A vssd1 vssd1 vccd1 vccd1 _1298_/B sky130_fd_sc_hd__or3_4
X_1338_ _1085_/A _1261_/X _1327_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1347_/A sky130_fd_sc_hd__a22o_1
X_1407_ input1/X _1375_/A _1406_/X _1807_/Q vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__a22o_1
X_1269_ _1586_/A _1630_/C vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1054_ _1722_/Q _0957_/X _1053_/X vssd1 vssd1 vccd1 vccd1 _1054_/X sky130_fd_sc_hd__a21o_1
X_1123_ _1009_/A _0992_/A _1123_/S vssd1 vssd1 vccd1 vccd1 _1125_/B sky130_fd_sc_hd__mux2_1
X_0907_ _0970_/A _1166_/B _0932_/B vssd1 vssd1 vccd1 vccd1 _1369_/C sky130_fd_sc_hd__a21oi_4
X_0838_ _0829_/Y input9/X _1806_/Q vssd1 vssd1 vccd1 vccd1 _0838_/Y sky130_fd_sc_hd__a21oi_2
Xoutput19 _1398_/X vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_4
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1741_ _1806_/CLK _1741_/D vssd1 vssd1 vccd1 vccd1 _1741_/Q sky130_fd_sc_hd__dfxtp_2
X_1810_ _1814_/CLK _1810_/D vssd1 vssd1 vccd1 vccd1 _1810_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1672_ _1814_/Q _1423_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1814_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1106_ _1723_/D _1722_/D _1241_/B _1105_/X vssd1 vssd1 vccd1 vccd1 _1239_/C sky130_fd_sc_hd__o211ai_4
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1037_ input3/X _0950_/X _1406_/C _1809_/Q vssd1 vssd1 vccd1 vccd1 _1037_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1724_ _1788_/CLK _1724_/D vssd1 vssd1 vccd1 vccd1 _1724_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _1586_/A _1655_/B _1586_/C _1589_/B vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__or4_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _1655_/A _1655_/B _1655_/C vssd1 vssd1 vccd1 vccd1 _1655_/X sky130_fd_sc_hd__and3_2
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1371_ _1701_/Q _1511_/A _1370_/Y vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__o21ai_4
X_1440_ _1369_/A _1510_/A _1725_/Q vssd1 vssd1 vccd1 vccd1 _1440_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1707_ _1826_/CLK _1707_/D vssd1 vssd1 vccd1 vccd1 _1707_/Q sky130_fd_sc_hd__dfxtp_1
X_1638_ _1788_/Q _1650_/S _1636_/X vssd1 vssd1 vccd1 vccd1 _1788_/D sky130_fd_sc_hd__o21a_1
X_1569_ input1/X _1762_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1762_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout87 _1697_/Q vssd1 vssd1 vccd1 vccd1 _0917_/A sky130_fd_sc_hd__clkbuf_2
Xfanout76 _1172_/A vssd1 vssd1 vccd1 vccd1 _1083_/A sky130_fd_sc_hd__clkbuf_16
Xfanout43 _1156_/X vssd1 vssd1 vccd1 vccd1 _1173_/C sky130_fd_sc_hd__buf_6
Xfanout54 _0952_/Y vssd1 vssd1 vccd1 vccd1 _1206_/A sky130_fd_sc_hd__buf_2
Xfanout65 _0876_/Y vssd1 vssd1 vccd1 vccd1 _1510_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0940_ _1065_/B _1065_/C vssd1 vssd1 vccd1 vccd1 _1050_/S sky130_fd_sc_hd__nand2_8
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0871_ _1372_/A _0957_/B _1369_/A _1369_/B vssd1 vssd1 vccd1 vccd1 _0878_/A sky130_fd_sc_hd__or4_4
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1354_ _0897_/A _0954_/B _0869_/B _1282_/B vssd1 vssd1 vccd1 vccd1 _1354_/X sky130_fd_sc_hd__o211a_1
X_1423_ _1745_/Q _1423_/A2 _1406_/X _1814_/Q _1422_/X vssd1 vssd1 vccd1 vccd1 _1423_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1285_ _1351_/C _1512_/D vssd1 vssd1 vccd1 vccd1 _1339_/C sky130_fd_sc_hd__or2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1070_ input1/X _0950_/X _1206_/A _1807_/Q vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0854_ _0917_/A _0909_/A vssd1 vssd1 vccd1 vccd1 _0894_/A sky130_fd_sc_hd__nand2b_2
X_0923_ _0941_/B _0973_/D _0923_/C _0923_/D vssd1 vssd1 vccd1 vccd1 _1114_/A sky130_fd_sc_hd__and4_4
X_1337_ _0850_/X _0933_/X _1353_/A _1374_/B vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__a211o_1
X_1268_ _1626_/C _1641_/C vssd1 vssd1 vccd1 vccd1 _1308_/A sky130_fd_sc_hd__or2_4
X_1406_ _1510_/A _1406_/B _1406_/C vssd1 vssd1 vccd1 vccd1 _1406_/X sky130_fd_sc_hd__or3_4
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1199_ _1199_/A _1199_/B vssd1 vssd1 vccd1 vccd1 _1736_/D sky130_fd_sc_hd__xor2_1
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ _1091_/A _1728_/D _1121_/X vssd1 vssd1 vccd1 vccd1 _1124_/B sky130_fd_sc_hd__a21oi_1
X_1053_ input2/X _0950_/X _1206_/A _1808_/Q vssd1 vssd1 vccd1 vccd1 _1053_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0906_ _0968_/A _1166_/B vssd1 vssd1 vccd1 vccd1 _1512_/B sky130_fd_sc_hd__nor2_1
X_0837_ _1799_/Q vssd1 vssd1 vccd1 vccd1 _0837_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1671_ _1813_/Q _1421_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1813_/D sky130_fd_sc_hd__mux2_1
X_1740_ _1806_/CLK _1740_/D vssd1 vssd1 vccd1 vccd1 _1740_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1105_ _1784_/Q _1105_/B vssd1 vssd1 vccd1 vccd1 _1105_/X sky130_fd_sc_hd__and2_2
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1036_ _1033_/Y _1035_/Y _1673_/B vssd1 vssd1 vccd1 vccd1 _1435_/B sky130_fd_sc_hd__mux2_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1654_ _1794_/Q _1653_/A _1652_/X _1653_/Y vssd1 vssd1 vccd1 vccd1 _1794_/D sky130_fd_sc_hd__a22o_1
X_1723_ _1825_/CLK _1723_/D vssd1 vssd1 vccd1 vccd1 _1723_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1655_/A _1589_/B vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__nor2_1
X_1019_ _1724_/Q _0957_/X _1018_/X vssd1 vssd1 vccd1 vccd1 _1019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1370_ _0933_/A _1336_/A _1163_/A _1515_/C vssd1 vssd1 vccd1 vccd1 _1370_/Y sky130_fd_sc_hd__a211oi_4
X_1637_ _1655_/A _1624_/B _1628_/B _1628_/A vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__o211a_1
X_1706_ _1826_/CLK _1706_/D vssd1 vssd1 vccd1 vccd1 _1706_/Q sky130_fd_sc_hd__dfxtp_1
X_1568_ _1695_/A _1568_/B vssd1 vssd1 vccd1 vccd1 _1576_/S sky130_fd_sc_hd__or2_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1499_ _1709_/Q _1498_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1709_/D sky130_fd_sc_hd__mux2_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout44 _1052_/S vssd1 vssd1 vccd1 vccd1 _1673_/B sky130_fd_sc_hd__buf_12
Xfanout55 _1549_/D vssd1 vssd1 vccd1 vccd1 _1648_/B sky130_fd_sc_hd__buf_4
Xfanout88 _0909_/A vssd1 vssd1 vccd1 vccd1 _1162_/A sky130_fd_sc_hd__buf_4
Xfanout77 _1373_/A vssd1 vssd1 vccd1 vccd1 _1298_/A sky130_fd_sc_hd__buf_6
Xfanout66 _0861_/Y vssd1 vssd1 vccd1 vccd1 _1479_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0870_ _1485_/A _1512_/A vssd1 vssd1 vccd1 vccd1 _0870_/X sky130_fd_sc_hd__or2_2
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1422_ input8/X _1375_/A _1377_/C _1719_/Q vssd1 vssd1 vccd1 vccd1 _1422_/X sky130_fd_sc_hd__a22o_1
X_1353_ _1353_/A _1353_/B _1353_/C _1309_/X vssd1 vssd1 vccd1 vccd1 _1699_/D sky130_fd_sc_hd__or4b_1
X_1284_ _1779_/Q _1284_/B vssd1 vssd1 vccd1 vccd1 _1366_/B sky130_fd_sc_hd__and2_1
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0999_ _1827_/Q _1682_/A _1500_/A _1714_/Q _0998_/X vssd1 vssd1 vccd1 vccd1 _0999_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0853_ _0914_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _1172_/A sky130_fd_sc_hd__or2_4
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0922_ _1512_/A _1512_/C vssd1 vssd1 vccd1 vccd1 _0923_/D sky130_fd_sc_hd__nor2_1
X_1405_ _1721_/Q _1377_/C _1375_/B _1381_/A vssd1 vssd1 vccd1 vccd1 _1405_/X sky130_fd_sc_hd__a211o_1
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_8
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1336_ _1336_/A _1336_/B _1334_/X _1335_/X vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__or4bb_2
X_1267_ _1586_/C _1267_/B vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__or2_2
X_1198_ _1199_/A _1199_/B vssd1 vssd1 vccd1 vccd1 _1203_/A sky130_fd_sc_hd__or2_1
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1052_ _1050_/X _1051_/X _1052_/S vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__mux2_4
X_1121_ _0985_/Y _1119_/X _1120_/X _0903_/Y vssd1 vssd1 vccd1 vccd1 _1121_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0905_ _0917_/A _1162_/C _1162_/B _1162_/A vssd1 vssd1 vccd1 vccd1 _1166_/B sky130_fd_sc_hd__or4bb_4
X_0836_ _1695_/A vssd1 vssd1 vccd1 vccd1 _0836_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1628_/B _1257_/B _1614_/B vssd1 vssd1 vccd1 vccd1 _1319_/Y sky130_fd_sc_hd__o21ai_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _1812_/Q _1419_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1812_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1035_ _1817_/Q _1457_/A _1034_/X vssd1 vssd1 vccd1 vccd1 _1035_/Y sky130_fd_sc_hd__o21ai_1
X_1104_ _1102_/A _1102_/B _1100_/A _1098_/A vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__o211ai_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1799_ _1799_/CLK _1799_/D vssd1 vssd1 vccd1 vccd1 _1799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1584_ _1602_/B _1580_/Y _1583_/Y _1276_/Y vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__a22o_1
X_1653_ _1653_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__nor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1788_/CLK _1722_/D vssd1 vssd1 vccd1 vccd1 _1722_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ input4/X _0950_/X _1206_/A _1810_/Q vssd1 vssd1 vccd1 vccd1 _1018_/X sky130_fd_sc_hd__a22o_1
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1705_ _1826_/CLK _1705_/D vssd1 vssd1 vccd1 vccd1 _1705_/Q sky130_fd_sc_hd__dfxtp_1
X_1636_ _1804_/D _1802_/D _1653_/A _1636_/D vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__or4_1
X_1567_ _1761_/Q _1566_/X _1567_/S vssd1 vssd1 vccd1 vccd1 _1761_/D sky130_fd_sc_hd__mux2_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1498_ input8/X _1373_/A _0970_/A _1496_/Y _1497_/X vssd1 vssd1 vccd1 vccd1 _1498_/X
+ sky130_fd_sc_hd__o32a_4
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 _1696_/Q vssd1 vssd1 vccd1 vccd1 _0909_/A sky130_fd_sc_hd__buf_4
Xfanout78 _0848_/Y vssd1 vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__buf_6
Xfanout56 _1549_/D vssd1 vssd1 vccd1 vccd1 _1653_/A sky130_fd_sc_hd__buf_2
Xfanout67 _0861_/Y vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__clkbuf_4
Xfanout45 _1050_/S vssd1 vssd1 vccd1 vccd1 _1457_/A sky130_fd_sc_hd__buf_6
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1421_ _1744_/Q _1423_/A2 _1406_/X _1813_/Q _1420_/X vssd1 vssd1 vccd1 vccd1 _1421_/X
+ sky130_fd_sc_hd__a221o_1
X_1352_ _1352_/A _1352_/B _1352_/C _1352_/D vssd1 vssd1 vccd1 vccd1 _1353_/C sky130_fd_sc_hd__or4_1
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1283_ _1165_/B _1406_/C vssd1 vssd1 vccd1 vccd1 _1339_/B sky130_fd_sc_hd__and2b_1
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0998_ _1819_/Q _1457_/A _1673_/B _0997_/X vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__o211a_1
X_1619_ _1779_/Q _1653_/A vssd1 vssd1 vccd1 vccd1 _1619_/X sky130_fd_sc_hd__and2_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0914_/A _0925_/B _0896_/X _1780_/Q _1568_/B vssd1 vssd1 vccd1 vccd1 _0923_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0852_ _0914_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _0926_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1335_ _0952_/A _1166_/B _1312_/Y _1165_/Y _0896_/X vssd1 vssd1 vccd1 vccd1 _1335_/X
+ sky130_fd_sc_hd__o311a_1
X_1404_ _1737_/Q _1381_/X _1402_/X _1403_/X vssd1 vssd1 vccd1 vccd1 _1404_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_8
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1266_ _1718_/Q _1778_/Q _1085_/B vssd1 vssd1 vccd1 vccd1 _1358_/B sky130_fd_sc_hd__o21a_1
X_1197_ _1736_/Q _1183_/Y _1196_/X vssd1 vssd1 vccd1 vccd1 _1199_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1051_ _1816_/Q _1703_/Q _1457_/A vssd1 vssd1 vccd1 vccd1 _1051_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ _1004_/A _1123_/S _0960_/B vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__a21bo_1
X_0904_ _0968_/A _0904_/B vssd1 vssd1 vccd1 vccd1 _0973_/B sky130_fd_sc_hd__or2_1
X_0835_ _1787_/Q vssd1 vssd1 vccd1 vccd1 _0835_/Y sky130_fd_sc_hd__inv_2
X_1318_ _1290_/B _1318_/B _1346_/B vssd1 vssd1 vccd1 vccd1 _1697_/D sky130_fd_sc_hd__nand3b_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ input1/X _1762_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1250_/B sky130_fd_sc_hd__mux2_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1103_ _1103_/A _1103_/B vssd1 vssd1 vccd1 vccd1 _1722_/D sky130_fd_sc_hd__xnor2_4
X_1034_ _1065_/B _1065_/C _1704_/Q vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1798_ _1803_/CLK _1798_/D vssd1 vssd1 vccd1 vccd1 _1798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ _1803_/CLK _1721_/D vssd1 vssd1 vccd1 vccd1 _1721_/Q sky130_fd_sc_hd__dfxtp_4
X_1583_ _1583_/A _1589_/B vssd1 vssd1 vccd1 vccd1 _1583_/Y sky130_fd_sc_hd__nor2_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _1802_/D _1652_/B _1655_/C vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__and3_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _1826_/Q _1682_/A _1500_/A _1713_/Q _1016_/X vssd1 vssd1 vccd1 vccd1 _1017_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1704_ _1825_/CLK _1704_/D vssd1 vssd1 vccd1 vccd1 _1704_/Q sky130_fd_sc_hd__dfxtp_1
X_1635_ _1787_/Q _1549_/D _1626_/X _1802_/D vssd1 vssd1 vccd1 vccd1 _1787_/D sky130_fd_sc_hd__a22o_1
X_1497_ _1496_/A _1496_/B _1485_/A vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__a21o_1
X_1566_ input7/X _1566_/A2 _1565_/X vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__o21a_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 _1513_/A vssd1 vssd1 vccd1 vccd1 _1372_/B sky130_fd_sc_hd__clkbuf_4
Xfanout57 _1577_/B vssd1 vssd1 vccd1 vccd1 _1549_/D sky130_fd_sc_hd__buf_4
Xfanout79 _1801_/Q vssd1 vssd1 vccd1 vccd1 _1560_/A sky130_fd_sc_hd__buf_4
Xfanout46 _0903_/Y vssd1 vssd1 vccd1 vccd1 _1063_/A sky130_fd_sc_hd__buf_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1420_ input7/X _1375_/A _1377_/C _1727_/Q vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__a22o_1
X_1351_ _1351_/A _1351_/B _1351_/C _1514_/A vssd1 vssd1 vccd1 vccd1 _1352_/D sky130_fd_sc_hd__or4_1
X_1282_ _1282_/A _1282_/B vssd1 vssd1 vccd1 vccd1 _1512_/D sky130_fd_sc_hd__nor2_1
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1618_ _1778_/Q _1617_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1778_/D sky130_fd_sc_hd__mux2_1
X_0997_ _1706_/Q _1673_/A vssd1 vssd1 vccd1 vccd1 _0997_/X sky130_fd_sc_hd__or2_1
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1549_ _1560_/A _1797_/Q _1796_/Q _1549_/D vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__or4_1
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ _0928_/A _1366_/A vssd1 vssd1 vccd1 vccd1 _1512_/C sky130_fd_sc_hd__or2_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0851_ _1162_/B _0868_/A _0954_/B vssd1 vssd1 vccd1 vccd1 _1166_/A sky130_fd_sc_hd__or3_4
X_1265_ _1718_/Q _1778_/Q _1262_/X _1264_/X vssd1 vssd1 vccd1 vccd1 _1352_/A sky130_fd_sc_hd__o31ai_1
X_1334_ _1298_/B _1084_/B _1166_/C _0932_/B vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__a31o_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1403_ _1114_/B _1368_/Y _1381_/B _1719_/Q vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1196_ _1727_/Q _1156_/X _1206_/B _1752_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1196_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1050_ _1711_/Q _1824_/Q _1050_/S vssd1 vssd1 vccd1 vccd1 _1050_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0834_ _1783_/Q vssd1 vssd1 vccd1 vccd1 _0834_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0903_ _1786_/Q _1513_/C vssd1 vssd1 vccd1 vccd1 _0903_/Y sky130_fd_sc_hd__nand2_2
X_1248_ input2/X _1763_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1252_/B sky130_fd_sc_hd__mux2_1
X_1317_ _1359_/A _1630_/C _1310_/X _1315_/X vssd1 vssd1 vccd1 vccd1 _1346_/B sky130_fd_sc_hd__o31a_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1723_/Q _1173_/C _1158_/Y _1732_/Q vssd1 vssd1 vccd1 vccd1 _1179_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102_ _1102_/A _1102_/B vssd1 vssd1 vccd1 vccd1 _1723_/D sky130_fd_sc_hd__xor2_4
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1033_ _1825_/Q _1457_/A _1032_/X vssd1 vssd1 vccd1 vccd1 _1033_/Y sky130_fd_sc_hd__a21oi_1
X_1797_ _1797_/CLK _1797_/D vssd1 vssd1 vccd1 vccd1 _1797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1651_ _1278_/Y _1588_/Y _1793_/Q _1648_/B vssd1 vssd1 vccd1 vccd1 _1793_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1720_ _1825_/CLK _1720_/D vssd1 vssd1 vccd1 vccd1 _1720_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _1628_/A _1802_/D vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__nor2_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1818_/Q _1050_/S _1052_/S _1015_/X vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__o211a_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1703_ _1825_/CLK _1703_/D vssd1 vssd1 vccd1 vccd1 _1703_/Q sky130_fd_sc_hd__dfxtp_1
X_1634_ _1786_/Q _1633_/Y _1650_/S vssd1 vssd1 vccd1 vccd1 _1786_/D sky130_fd_sc_hd__mux2_1
X_1496_ _1496_/A _1496_/B vssd1 vssd1 vccd1 vccd1 _1496_/Y sky130_fd_sc_hd__nor2_1
X_1565_ _1560_/A _1727_/Q _1560_/Y _1564_/Y _1549_/D vssd1 vssd1 vccd1 vccd1 _1565_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout69 _1513_/A vssd1 vssd1 vccd1 vccd1 _0957_/B sky130_fd_sc_hd__buf_6
Xfanout58 _1344_/A vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__buf_4
Xfanout47 _1277_/B vssd1 vssd1 vccd1 vccd1 _1641_/C sky130_fd_sc_hd__buf_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1281_ _1083_/A _0912_/B _1364_/A vssd1 vssd1 vccd1 vccd1 _1351_/C sky130_fd_sc_hd__o21ai_1
X_1350_ _0869_/B _0970_/B _0973_/C vssd1 vssd1 vccd1 vccd1 _1514_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0996_ _0995_/X _0996_/B vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__nand2b_4
X_1617_ _1628_/B _1300_/Y _1583_/Y vssd1 vssd1 vccd1 vccd1 _1617_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1479_ _1725_/Q input5/X _1479_/S vssd1 vssd1 vccd1 vccd1 _1479_/X sky130_fd_sc_hd__mux2_2
X_1548_ _1758_/Q _1547_/X _1548_/S vssd1 vssd1 vccd1 vccd1 _1758_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ _0897_/A _0897_/B _0927_/A _0909_/A vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__and4b_1
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1402_ _1753_/Q _1381_/C _1378_/Y input8/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1402_/X
+ sky130_fd_sc_hd__a221o_1
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_8
X_1333_ _1342_/B _1333_/B _1359_/B _1333_/D vssd1 vssd1 vccd1 vccd1 _1336_/B sky130_fd_sc_hd__and4_1
X_1264_ _1779_/Q _0888_/Y _1359_/A _1260_/X _1263_/X vssd1 vssd1 vccd1 vccd1 _1264_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1195_ _1195_/A _1195_/B vssd1 vssd1 vccd1 vccd1 _1735_/D sky130_fd_sc_hd__xor2_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0979_ _0993_/S _1004_/A _0966_/Y vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__a21bo_1
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _1780_/Q vssd1 vssd1 vccd1 vccd1 _0833_/Y sky130_fd_sc_hd__inv_2
X_0902_ _1786_/Q _1513_/C vssd1 vssd1 vccd1 vccd1 _1091_/A sky130_fd_sc_hd__and2_2
X_1247_ input3/X _1764_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1256_/B sky130_fd_sc_hd__mux2_4
X_1178_ _0828_/Y _1772_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1178_/X sky130_fd_sc_hd__o21a_2
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1316_ _1341_/A _1340_/B _1309_/X vssd1 vssd1 vccd1 vccd1 _1318_/B sky130_fd_sc_hd__nor3b_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1101_ _1031_/S _1030_/B _1100_/A _1100_/B vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__o22a_2
X_1032_ _1712_/Q _1065_/B _1065_/C vssd1 vssd1 vccd1 vccd1 _1032_/X sky130_fd_sc_hd__and3_1
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1796_ _1799_/CLK _1796_/D vssd1 vssd1 vccd1 vccd1 _1796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1581_ _1804_/D _1624_/B vssd1 vssd1 vccd1 vccd1 _1589_/B sky130_fd_sc_hd__nand2_4
X_1650_ _1792_/Q _1643_/C _1650_/S vssd1 vssd1 vccd1 vccd1 _1792_/D sky130_fd_sc_hd__mux2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1015_ _1705_/Q _1673_/A vssd1 vssd1 vccd1 vccd1 _1015_/X sky130_fd_sc_hd__or2_1
X_1779_ _1799_/CLK _1779_/D vssd1 vssd1 vccd1 vccd1 _1779_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1633_ _1653_/B _1633_/B vssd1 vssd1 vccd1 vccd1 _1633_/Y sky130_fd_sc_hd__nor2_1
X_1702_ _1830_/CLK _1702_/D vssd1 vssd1 vccd1 vccd1 _1702_/Q sky130_fd_sc_hd__dfxtp_1
X_1564_ _1564_/A _1564_/B vssd1 vssd1 vccd1 vccd1 _1564_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1495_ _1719_/Q _1495_/B vssd1 vssd1 vccd1 vccd1 _1496_/B sky130_fd_sc_hd__xnor2_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout59 _1577_/B vssd1 vssd1 vccd1 vccd1 _1344_/A sky130_fd_sc_hd__buf_2
Xfanout48 _0957_/A vssd1 vssd1 vccd1 vccd1 _1372_/A sky130_fd_sc_hd__buf_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1280_ _1344_/A _1655_/B _1344_/C _1641_/B vssd1 vssd1 vccd1 vccd1 _1364_/A sky130_fd_sc_hd__or4_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0995_ _0995_/A _1124_/A vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__or2_2
X_1616_ _1777_/Q _1615_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1777_/D sky130_fd_sc_hd__mux2_1
X_1547_ input8/X _1719_/Q _1547_/S vssd1 vssd1 vccd1 vccd1 _1547_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1478_ _1705_/Q _1477_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1705_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ _1736_/Q _1381_/X _1399_/X _1400_/X vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__o22a_1
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
X_1332_ _1344_/B _1310_/X _1330_/X _1308_/A _1331_/X vssd1 vssd1 vccd1 vccd1 _1333_/D
+ sky130_fd_sc_hd__o221a_1
X_1263_ _1373_/A _0904_/B _1511_/B _0874_/X vssd1 vssd1 vccd1 vccd1 _1263_/X sky130_fd_sc_hd__o211a_1
X_1194_ _1195_/A _1195_/B vssd1 vssd1 vccd1 vccd1 _1199_/A sky130_fd_sc_hd__or2_1
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0978_ _1788_/Q _1513_/C _0977_/Y vssd1 vssd1 vccd1 vccd1 _1041_/A sky130_fd_sc_hd__a21oi_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0832_ _1795_/Q vssd1 vssd1 vccd1 vccd1 _0832_/Y sky130_fd_sc_hd__inv_2
X_0901_ _1105_/B _1406_/B vssd1 vssd1 vccd1 vccd1 _1513_/C sky130_fd_sc_hd__or2_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1315_ _0897_/A _0973_/B _1357_/A _0973_/C vssd1 vssd1 vccd1 vccd1 _1315_/X sky130_fd_sc_hd__o211a_1
X_1246_ _1256_/A _1344_/C vssd1 vssd1 vccd1 vccd1 _1614_/B sky130_fd_sc_hd__nand2_4
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1177_ _1182_/A _1177_/B vssd1 vssd1 vccd1 vccd1 _1731_/D sky130_fd_sc_hd__nor2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1830_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1100_ _1100_/A _1100_/B vssd1 vssd1 vccd1 vccd1 _1100_/Y sky130_fd_sc_hd__nor2_1
X_1031_ _1029_/Y _1030_/X _1031_/S vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__mux2_4
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1795_ _1804_/CLK _1795_/D vssd1 vssd1 vccd1 vccd1 _1795_/Q sky130_fd_sc_hd__dfxtp_1
X_1229_ _1228_/A _1228_/B _1228_/C vssd1 vssd1 vccd1 vccd1 _1230_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1580_ _1580_/A _1589_/A vssd1 vssd1 vccd1 vccd1 _1580_/Y sky130_fd_sc_hd__nor2_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1014_ _1014_/A _1014_/B vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__or2_2
X_1778_ _1794_/CLK _1778_/D vssd1 vssd1 vccd1 vccd1 _1778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1701_ _1806_/CLK _1701_/D _1695_/Y vssd1 vssd1 vccd1 vccd1 _1701_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1632_ _1785_/Q _1648_/B _1602_/X _1631_/X vssd1 vssd1 vccd1 vccd1 _1785_/D sky130_fd_sc_hd__a22o_1
X_1494_ _1485_/B _1488_/X _1489_/Y vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__a21bo_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1719_/Q _1718_/Q vssd1 vssd1 vccd1 vccd1 _1564_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout49 _1378_/Y vssd1 vssd1 vccd1 vccd1 _1514_/B sky130_fd_sc_hd__buf_6
Xfanout38 _1518_/X vssd1 vssd1 vccd1 vccd1 _1666_/S sky130_fd_sc_hd__buf_6
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0994_ _0994_/A _0994_/B vssd1 vssd1 vccd1 vccd1 _1124_/A sky130_fd_sc_hd__nor2_2
X_1615_ _1628_/B _1641_/B _1614_/Y _1613_/Y _1588_/B vssd1 vssd1 vccd1 vccd1 _1615_/X
+ sky130_fd_sc_hd__a32o_1
X_1546_ _1510_/A _1545_/X _1536_/X vssd1 vssd1 vccd1 vccd1 _1548_/S sky130_fd_sc_hd__o21a_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1477_ _1476_/Y input4/X _1479_/S vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__mux2_4
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1331_ _1630_/C _1308_/A _1319_/Y _1260_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1331_/X
+ sky130_fd_sc_hd__o2111a_1
X_1400_ _0948_/B _1368_/Y _1381_/B _1727_/Q vssd1 vssd1 vccd1 vccd1 _1400_/X sky130_fd_sc_hd__a2bb2o_1
Xinput6 io_in[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
X_1262_ _1779_/Q _1083_/A _1083_/B _1084_/B _1298_/A vssd1 vssd1 vccd1 vccd1 _1262_/X
+ sky130_fd_sc_hd__o32a_1
X_1193_ _1735_/Q _1183_/Y _1192_/X vssd1 vssd1 vccd1 vccd1 _1195_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0977_ _0977_/A _1513_/C _1510_/B vssd1 vssd1 vccd1 vccd1 _0977_/Y sky130_fd_sc_hd__nor3_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1529_ _1779_/Q _1549_/D _1510_/A _1783_/Q vssd1 vssd1 vccd1 vccd1 _1529_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _1297_/A _1554_/S vssd1 vssd1 vccd1 vccd1 _1406_/B sky130_fd_sc_hd__or2_4
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0831_ _1797_/Q vssd1 vssd1 vccd1 vccd1 _0831_/Y sky130_fd_sc_hd__inv_2
X_1314_ _1344_/A _1630_/C _1636_/D _1626_/C vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__or4_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1245_ input4/X _1765_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1344_/C sky130_fd_sc_hd__mux2_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1176_ _1175_/B _1181_/B vssd1 vssd1 vccd1 vccd1 _1177_/B sky130_fd_sc_hd__and2b_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1030_ _1125_/A _1030_/B vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__or2_1
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ _1794_/CLK _1794_/D vssd1 vssd1 vccd1 vccd1 _1794_/Q sky130_fd_sc_hd__dfxtp_1
X_1228_ _1228_/A _1228_/B _1228_/C vssd1 vssd1 vccd1 vccd1 _1234_/A sky130_fd_sc_hd__and3_1
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1159_ _1579_/A _1577_/B vssd1 vssd1 vccd1 vccd1 _1206_/B sky130_fd_sc_hd__nor2_8
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1013_ _1125_/A _1012_/B _1012_/A vssd1 vssd1 vccd1 vccd1 _1014_/B sky130_fd_sc_hd__o21a_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1777_ _1794_/CLK _1777_/D vssd1 vssd1 vccd1 vccd1 _1777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1825_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1700_ _1769_/CLK _1700_/D _1694_/Y vssd1 vssd1 vccd1 vccd1 _1700_/Q sky130_fd_sc_hd__dfrtp_1
X_1631_ _1655_/A _1628_/B _1630_/X vssd1 vssd1 vccd1 vccd1 _1631_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1493_ _1708_/Q _1492_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1708_/D sky130_fd_sc_hd__mux2_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1729_/Q _1728_/Q vssd1 vssd1 vccd1 vccd1 _1564_/A sky130_fd_sc_hd__xor2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 _1518_/X vssd1 vssd1 vccd1 vccd1 _1672_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1829_ _1829_/CLK _1829_/D vssd1 vssd1 vccd1 vccd1 _1829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0993_ _1009_/A _0992_/A _0993_/S vssd1 vssd1 vccd1 vccd1 _0995_/A sky130_fd_sc_hd__mux2_1
X_1614_ _1630_/C _1614_/B vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__nand2_1
X_1545_ _1792_/Q _1105_/B _1566_/A2 _1542_/S vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__a211o_1
X_1476_ _1476_/A _1476_/B vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1330_ _1580_/A _1644_/B _1320_/C vssd1 vssd1 vccd1 vccd1 _1330_/X sky130_fd_sc_hd__o21a_1
X_1261_ _1718_/Q _1779_/Q _1778_/Q vssd1 vssd1 vccd1 vccd1 _1261_/X sky130_fd_sc_hd__or3_1
Xinput7 io_in[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_8
X_1192_ _1726_/Q _1173_/C _1206_/B _1751_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1192_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ _0966_/Y _0993_/S vssd1 vssd1 vccd1 vccd1 _0986_/S sky130_fd_sc_hd__and2b_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1528_ _1560_/A _1697_/Q _1799_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__or4_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1459_ _1702_/Q _1458_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1702_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0830_ _0897_/B vssd1 vssd1 vccd1 vccd1 _0868_/A sky130_fd_sc_hd__clkinv_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1244_ _1256_/A _1652_/B vssd1 vssd1 vccd1 vccd1 _1344_/B sky130_fd_sc_hd__nand2_1
X_1313_ _0950_/B _1312_/Y _1512_/B vssd1 vssd1 vccd1 vccd1 _1340_/B sky130_fd_sc_hd__a21o_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ _1181_/B _1175_/B vssd1 vssd1 vccd1 vccd1 _1182_/A sky130_fd_sc_hd__and2b_1
X_0959_ input7/X _0950_/X _0958_/X vssd1 vssd1 vccd1 vccd1 _0960_/B sky130_fd_sc_hd__a21oi_4
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 io_in[9] vssd1 vssd1 vccd1 vccd1 _1805_/D sky130_fd_sc_hd__clkbuf_2
X_1793_ _1799_/CLK _1793_/D vssd1 vssd1 vccd1 vccd1 _1793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1227_ input6/X _1156_/B _1205_/Y _1743_/Q _1226_/X vssd1 vssd1 vccd1 vccd1 _1228_/C
+ sky130_fd_sc_hd__a221o_1
X_1158_ _0957_/B _1510_/B _1173_/C _1205_/A vssd1 vssd1 vccd1 vccd1 _1158_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1089_ _0835_/Y _1082_/X _1088_/X vssd1 vssd1 vccd1 vccd1 _1090_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ _1012_/A _1012_/B vssd1 vssd1 vccd1 vccd1 _1014_/A sky130_fd_sc_hd__nor2_2
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1776_ _1794_/CLK _1776_/D vssd1 vssd1 vccd1 vccd1 _1776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1630_ _1641_/C _1630_/B _1630_/C vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__and3b_1
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1561_ _1560_/A _1782_/Q _1793_/Q _1549_/D _1545_/X vssd1 vssd1 vccd1 vccd1 _1567_/S
+ sky130_fd_sc_hd__o41a_1
X_1492_ _1490_/Y _1491_/X input7/X _1479_/S vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1759_ _1803_/CLK _1759_/D vssd1 vssd1 vccd1 vccd1 _1759_/Q sky130_fd_sc_hd__dfxtp_2
X_1828_ _1829_/CLK _1828_/D vssd1 vssd1 vccd1 vccd1 _1828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0992_ _0992_/A _1125_/A vssd1 vssd1 vccd1 vccd1 _1009_/A sky130_fd_sc_hd__nor2_1
X_1613_ _1641_/B _1633_/B vssd1 vssd1 vccd1 vccd1 _1613_/Y sky130_fd_sc_hd__nor2_2
X_1544_ _1757_/Q _1543_/X _1544_/S vssd1 vssd1 vccd1 vccd1 _1757_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1769_/CLK sky130_fd_sc_hd__clkbuf_8
X_1475_ _1724_/Q _1475_/B vssd1 vssd1 vccd1 vccd1 _1476_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 io_in[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_6
X_1260_ _1655_/B _1636_/D _1630_/B _1259_/X vssd1 vssd1 vccd1 vccd1 _1260_/X sky130_fd_sc_hd__o31a_2
X_1191_ _1191_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1734_/D sky130_fd_sc_hd__xor2_1
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0975_ _1735_/Q _0950_/B _0974_/X input6/X vssd1 vssd1 vccd1 vccd1 _0993_/S sky130_fd_sc_hd__a22o_2
X_1527_ _1782_/Q _1785_/Q _1783_/Q vssd1 vssd1 vccd1 vccd1 _1532_/S sky130_fd_sc_hd__or3_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1389_ _1732_/Q _1381_/X _1387_/X _1388_/X vssd1 vssd1 vccd1 vccd1 _1389_/X sky130_fd_sc_hd__o22a_1
X_1458_ _1721_/Q input1/X _1479_/S vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__mux2_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1243_ _1256_/A _1652_/B vssd1 vssd1 vccd1 vccd1 _1655_/B sky130_fd_sc_hd__and2_4
X_1312_ _1802_/Q _1312_/B vssd1 vssd1 vccd1 vccd1 _1312_/Y sky130_fd_sc_hd__xnor2_2
X_1174_ _1731_/Q _1158_/Y _1206_/B _1747_/Q _1171_/X vssd1 vssd1 vccd1 vccd1 _1175_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0889_ _1162_/C _0894_/A vssd1 vssd1 vccd1 vccd1 _0904_/B sky130_fd_sc_hd__or2_2
X_0958_ _1813_/Q _1406_/C _0957_/X _1727_/Q _0948_/Y vssd1 vssd1 vccd1 vccd1 _0958_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 rst vssd1 vssd1 vccd1 vccd1 _1695_/A sky130_fd_sc_hd__buf_6
X_1792_ _1799_/CLK _1792_/D vssd1 vssd1 vccd1 vccd1 _1792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1226_ _1726_/Q _1173_/D _1206_/X _1812_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1226_/X
+ sky130_fd_sc_hd__a221o_1
X_1157_ _1579_/A _1510_/B vssd1 vssd1 vccd1 vccd1 _1205_/A sky130_fd_sc_hd__nand2_8
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1088_ _1369_/C _1088_/B _1358_/A _0956_/X vssd1 vssd1 vccd1 vccd1 _1088_/X sky130_fd_sc_hd__or4b_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ _1010_/A _0992_/A _1011_/S vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1775_ _1794_/CLK _1775_/D vssd1 vssd1 vccd1 vccd1 _1775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ _1212_/A _1212_/B vssd1 vssd1 vccd1 vccd1 _1738_/D sky130_fd_sc_hd__xor2_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1560_ _1560_/A _1793_/Q vssd1 vssd1 vccd1 vccd1 _1560_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1491_ _1485_/B _1488_/X _1489_/Y _1479_/S vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__a31o_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1827_ _1829_/CLK _1827_/D vssd1 vssd1 vccd1 vccd1 _1827_/Q sky130_fd_sc_hd__dfxtp_1
X_1758_ _1803_/CLK _1758_/D vssd1 vssd1 vccd1 vccd1 _1758_/Q sky130_fd_sc_hd__dfxtp_1
X_1689_ _1829_/Q _1492_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1829_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0991_ _1125_/A vssd1 vssd1 vccd1 vccd1 _0994_/B sky130_fd_sc_hd__inv_2
X_1612_ _1593_/A _1608_/X _1611_/X _1626_/B _1776_/Q vssd1 vssd1 vccd1 vccd1 _1776_/D
+ sky130_fd_sc_hd__o32a_1
X_1543_ _1541_/Y _1542_/X _1543_/S vssd1 vssd1 vccd1 vccd1 _1543_/X sky130_fd_sc_hd__mux2_1
X_1474_ _1465_/B _1468_/X _1469_/Y vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__a21bo_1
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_in[8] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
X_1190_ _1191_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1195_/A sky130_fd_sc_hd__or2_1
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0974_ _1516_/A _0974_/B vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__and2b_4
X_1526_ _1753_/Q _1404_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1753_/D sky130_fd_sc_hd__mux2_1
X_1457_ _1457_/A _1673_/B _1682_/B vssd1 vssd1 vccd1 vccd1 _1499_/S sky130_fd_sc_hd__and3_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1388_ _1435_/B _1368_/Y _1381_/B _1723_/Q vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1804_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ _1758_/Q _1761_/Q _1754_/Q _1757_/Q _1803_/Q _1804_/Q vssd1 vssd1 vccd1 vccd1
+ _1312_/B sky130_fd_sc_hd__mux4_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1242_ input5/X _1766_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1242_/X sky130_fd_sc_hd__mux2_1
X_1173_ _1372_/B _1510_/B _1173_/C _1173_/D vssd1 vssd1 vccd1 vccd1 _1205_/B sky130_fd_sc_hd__or4_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0888_ _1284_/B vssd1 vssd1 vccd1 vccd1 _0888_/Y sky130_fd_sc_hd__inv_2
X_0957_ _0957_/A _0957_/B _0956_/X vssd1 vssd1 vccd1 vccd1 _0957_/X sky130_fd_sc_hd__or3b_4
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1509_ _1166_/B _1373_/B _1701_/Q vssd1 vssd1 vccd1 vccd1 _1517_/A sky130_fd_sc_hd__a21oi_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1791_ _1797_/CLK _1791_/D vssd1 vssd1 vccd1 vccd1 _1791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1225_ _1228_/A _1228_/B vssd1 vssd1 vccd1 vccd1 _1742_/D sky130_fd_sc_hd__xor2_1
X_1156_ _1206_/A _1156_/B vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__or2_2
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1087_ _0925_/B _0912_/B _1373_/A vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__a21oi_2
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1010_ _1010_/A vssd1 vssd1 vccd1 vccd1 _1010_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1774_ _1799_/CLK _1774_/D vssd1 vssd1 vccd1 vccd1 _1774_/Q sky130_fd_sc_hd__dfxtp_1
X_1208_ input1/X _1156_/B _1205_/Y _1738_/Q _1207_/X vssd1 vssd1 vccd1 vccd1 _1212_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ _1139_/A _1139_/B vssd1 vssd1 vccd1 vccd1 _1141_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1490_ _1488_/X _1489_/Y _1485_/B vssd1 vssd1 vccd1 vccd1 _1490_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1826_ _1826_/CLK _1826_/D vssd1 vssd1 vccd1 vccd1 _1826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1757_ _1803_/CLK _1757_/D vssd1 vssd1 vccd1 vccd1 _1757_/Q sky130_fd_sc_hd__dfxtp_1
X_1688_ _1828_/Q _1486_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1828_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1611_ _1300_/Y _1583_/Y _1596_/Y _1602_/B vssd1 vssd1 vccd1 vccd1 _1611_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0990_ _1791_/Q _1513_/C vssd1 vssd1 vccd1 vccd1 _1125_/A sky130_fd_sc_hd__and2_4
X_1542_ _1722_/Q input2/X _1542_/S vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__mux2_1
X_1473_ _1704_/Q _1472_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1704_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1809_ _1814_/CLK _1809_/D vssd1 vssd1 vccd1 vccd1 _1809_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0973_ _0950_/X _0973_/B _0973_/C _0973_/D vssd1 vssd1 vccd1 vccd1 _0974_/B sky130_fd_sc_hd__and4b_1
X_1525_ _1752_/Q _1401_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1752_/D sky130_fd_sc_hd__mux2_1
X_1456_ _1456_/A _1456_/B _1456_/C vssd1 vssd1 vccd1 vccd1 _1682_/B sky130_fd_sc_hd__nand3_4
X_1387_ _1748_/Q _1381_/C _1514_/B input3/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1387_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1310_ _1636_/D _1641_/B _1614_/B vssd1 vssd1 vccd1 vccd1 _1310_/X sky130_fd_sc_hd__a21o_1
X_1241_ _1100_/Y _1241_/B vssd1 vssd1 vccd1 vccd1 _1724_/D sky130_fd_sc_hd__and2b_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1172_ _1172_/A _1172_/B vssd1 vssd1 vccd1 vccd1 _1173_/D sky130_fd_sc_hd__nor2_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0956_ _1345_/A _1363_/A vssd1 vssd1 vccd1 vccd1 _0956_/X sky130_fd_sc_hd__and2_1
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0887_ _1513_/B _0977_/A _1374_/A _0887_/D vssd1 vssd1 vccd1 vccd1 _1284_/B sky130_fd_sc_hd__or4_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ _1717_/Q _1498_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1717_/D sky130_fd_sc_hd__mux2_1
X_1439_ _1445_/A _1017_/Y _1438_/X vssd1 vssd1 vccd1 vccd1 _1439_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _1797_/CLK _1790_/D vssd1 vssd1 vccd1 vccd1 _1790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1224_ input5/X _1156_/B _1205_/Y _1742_/Q _1223_/X vssd1 vssd1 vccd1 vccd1 _1228_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1155_ _0933_/A _1336_/A _1163_/A _1151_/Y vssd1 vssd1 vccd1 vccd1 _1156_/B sky130_fd_sc_hd__a211o_4
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1086_ _1406_/C _1515_/C _1718_/Q vssd1 vssd1 vccd1 vccd1 _1088_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0939_ _1065_/B _1065_/C vssd1 vssd1 vccd1 vccd1 _1673_/A sky130_fd_sc_hd__and2_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1767_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1773_ _1804_/CLK _1773_/D vssd1 vssd1 vccd1 vccd1 _1773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1207_ _1721_/Q _1173_/D _1206_/X _1807_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1207_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1138_ _1125_/A _1137_/B _1137_/A vssd1 vssd1 vccd1 vccd1 _1139_/B sky130_fd_sc_hd__o21ai_1
X_1069_ _1066_/Y _1068_/Y _1673_/B vssd1 vssd1 vccd1 vccd1 _1428_/B sky130_fd_sc_hd__mux2_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1756_ _1807_/CLK input8/X vssd1 vssd1 vccd1 vccd1 _1756_/Q sky130_fd_sc_hd__dfxtp_1
X_1825_ _1825_/CLK _1825_/D vssd1 vssd1 vccd1 vccd1 _1825_/Q sky130_fd_sc_hd__dfxtp_1
X_1687_ _1827_/Q _1479_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1827_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610_ _1775_/Q _1626_/B _1609_/X vssd1 vssd1 vccd1 vccd1 _1775_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1541_ _1541_/A _1541_/B vssd1 vssd1 vccd1 vccd1 _1541_/Y sky130_fd_sc_hd__nor2_1
X_1472_ _1470_/Y _1471_/X input3/X _1479_/S vssd1 vssd1 vccd1 vccd1 _1472_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1739_ _1807_/CLK _1739_/D vssd1 vssd1 vccd1 vccd1 _1739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ _1808_/CLK _1808_/D vssd1 vssd1 vccd1 vccd1 _1808_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0972_ _0972_/A _1351_/B _0912_/X _1557_/S vssd1 vssd1 vccd1 vccd1 _1516_/A sky130_fd_sc_hd__or4bb_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1524_ _1751_/Q _1398_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1751_/D sky130_fd_sc_hd__mux2_1
X_1455_ _1577_/B _1560_/A _1771_/Q vssd1 vssd1 vccd1 vccd1 _1456_/C sky130_fd_sc_hd__or3b_4
X_1386_ _1731_/Q _1381_/X _1384_/X _1385_/X vssd1 vssd1 vccd1 vccd1 _1386_/X sky130_fd_sc_hd__o22a_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1171_ _1772_/Q _0860_/X _1173_/C _1722_/Q vssd1 vssd1 vccd1 vccd1 _1171_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1240_ _1240_/A _1240_/B vssd1 vssd1 vccd1 vccd1 _1725_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0886_ _0954_/B _0968_/A _0953_/C vssd1 vssd1 vccd1 vccd1 _0887_/D sky130_fd_sc_hd__nor3_1
X_0955_ _1166_/A _1282_/B _1172_/B _0932_/B vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__a31o_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1507_ _1716_/Q _1492_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1716_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1369_ _1369_/A _1369_/B _1369_/C vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__or3_4
X_1438_ _1759_/Q _1424_/X _1425_/Y _1724_/Q _1437_/X vssd1 vssd1 vccd1 vccd1 _1438_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1223_ _1725_/Q _1173_/D _1206_/X _1811_/Q _1372_/B vssd1 vssd1 vccd1 vccd1 _1223_/X
+ sky130_fd_sc_hd__a221o_1
X_1154_ _1701_/Q _1172_/B vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__nor2_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _1085_/A _1085_/B vssd1 vssd1 vccd1 vccd1 _1515_/C sky130_fd_sc_hd__or2_4
X_0869_ _1083_/A _0869_/B vssd1 vssd1 vccd1 vccd1 _1512_/A sky130_fd_sc_hd__nor2_2
X_0938_ _1773_/Q _1566_/A2 _0941_/C _0937_/X vssd1 vssd1 vccd1 vccd1 _1065_/C sky130_fd_sc_hd__a211o_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1772_ _1806_/CLK _1772_/D vssd1 vssd1 vccd1 vccd1 _1772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1206_ _1206_/A _1206_/B vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__or2_4
X_1137_ _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _1139_/A sky130_fd_sc_hd__or2_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1068_ _1815_/Q _1457_/A _1067_/X vssd1 vssd1 vccd1 vccd1 _1068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1794_/CLK sky130_fd_sc_hd__clkbuf_8
X_1755_ _1830_/CLK _1755_/D vssd1 vssd1 vccd1 vccd1 _1755_/Q sky130_fd_sc_hd__dfxtp_1
X_1824_ _1825_/CLK _1824_/D vssd1 vssd1 vccd1 vccd1 _1824_/Q sky130_fd_sc_hd__dfxtp_1
X_1686_ _1826_/Q _1477_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1826_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1540_ _1721_/Q _1722_/Q _1723_/Q _1724_/Q vssd1 vssd1 vccd1 vccd1 _1541_/B sky130_fd_sc_hd__or4_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1471_ _1465_/B _1468_/X _1469_/Y _1479_/S vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__a31o_1
XFILLER_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1807_ _1807_/CLK _1807_/D vssd1 vssd1 vccd1 vccd1 _1807_/Q sky130_fd_sc_hd__dfxtp_1
X_1669_ _1811_/Q _1417_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1811_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1738_ _1807_/CLK _1738_/D vssd1 vssd1 vccd1 vccd1 _1738_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0971_ _0850_/X _0933_/X _1286_/B vssd1 vssd1 vccd1 vccd1 _1351_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1523_ _1750_/Q _1395_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1750_/D sky130_fd_sc_hd__mux2_1
X_1454_ _1758_/Q _1424_/X _1452_/X _1453_/X vssd1 vssd1 vccd1 vccd1 _1454_/X sky130_fd_sc_hd__a211o_2
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1385_ _1052_/X _1381_/A _1381_/B _1722_/Q vssd1 vssd1 vccd1 vccd1 _1385_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1170_ _1170_/A _1170_/B vssd1 vssd1 vccd1 vccd1 _1730_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0954_ _1162_/C _0954_/B _1162_/B vssd1 vssd1 vccd1 vccd1 _1172_/B sky130_fd_sc_hd__or3b_4
X_0885_ _1511_/A _0919_/A vssd1 vssd1 vccd1 vccd1 _1374_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1437_ _1733_/Q _1372_/A _1369_/B _1741_/Q vssd1 vssd1 vccd1 vccd1 _1437_/X sky130_fd_sc_hd__a22o_1
X_1506_ _1715_/Q _1486_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1715_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1299_ _1586_/C _1641_/B vssd1 vssd1 vccd1 vccd1 _1300_/A sky130_fd_sc_hd__or2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1368_ _1369_/A _1369_/B _1369_/C vssd1 vssd1 vccd1 vccd1 _1368_/Y sky130_fd_sc_hd__nor3_4
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1222_ _1228_/A _1222_/B vssd1 vssd1 vccd1 vccd1 _1741_/D sky130_fd_sc_hd__nor2_1
X_1153_ _1298_/B _1282_/A vssd1 vssd1 vccd1 vccd1 _1163_/A sky130_fd_sc_hd__nor2_2
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1084_ _1298_/A _1084_/B vssd1 vssd1 vccd1 vccd1 _1085_/B sky130_fd_sc_hd__nor2_1
X_0937_ _0928_/A _1366_/A _1286_/A _1777_/Q vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__o31a_1
X_0868_ _0868_/A _1083_/A _0926_/B vssd1 vssd1 vccd1 vccd1 _1624_/C sky130_fd_sc_hd__or3b_4
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _1799_/CLK _1771_/D vssd1 vssd1 vccd1 vccd1 _1771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1205_ _1205_/A _1205_/B vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1067_ _1065_/B _1065_/C _1702_/Q vssd1 vssd1 vccd1 vccd1 _1067_/X sky130_fd_sc_hd__a21o_1
X_1136_ _1125_/A _1137_/A _1137_/B vssd1 vssd1 vccd1 vccd1 _1729_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1823_ _1830_/CLK _1823_/D vssd1 vssd1 vccd1 vccd1 _1823_/Q sky130_fd_sc_hd__dfxtp_1
X_1754_ _1803_/CLK _1754_/D vssd1 vssd1 vccd1 vccd1 _1754_/Q sky130_fd_sc_hd__dfxtp_2
X_1685_ _1825_/Q _1472_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1825_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1119_ _1004_/A _1024_/A _1119_/S vssd1 vssd1 vccd1 vccd1 _1119_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1470_ _1468_/X _1469_/Y _1465_/B vssd1 vssd1 vccd1 vccd1 _1470_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1806_ _1806_/CLK _1806_/D vssd1 vssd1 vccd1 vccd1 _1806_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _1810_/Q _1415_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1810_/D sky130_fd_sc_hd__mux2_1
X_1737_ _1807_/CLK _1737_/D vssd1 vssd1 vccd1 vccd1 _1737_/Q sky130_fd_sc_hd__dfxtp_2
X_1599_ _1655_/A _1655_/B _1589_/Y _1598_/X vssd1 vssd1 vccd1 vccd1 _1599_/X sky130_fd_sc_hd__a31o_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1803_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0970_ _0970_/A _0970_/B vssd1 vssd1 vccd1 vccd1 _1286_/B sky130_fd_sc_hd__nor2_1
X_1453_ _1445_/A _1114_/B _1425_/Y _1719_/Q vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__a2bb2o_1
X_1522_ _1749_/Q _1392_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1749_/D sky130_fd_sc_hd__mux2_1
X_1384_ _1747_/Q _1381_/C _1514_/B input2/X _1410_/B1 vssd1 vssd1 vccd1 vccd1 _1384_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0953_ _0954_/B _1172_/A _0953_/C vssd1 vssd1 vccd1 vccd1 _1345_/A sky130_fd_sc_hd__or3_4
X_0884_ _0933_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__nand2_2
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1367_ _1367_/A _1372_/C _1367_/C vssd1 vssd1 vccd1 vccd1 _1701_/D sky130_fd_sc_hd__or3_1
X_1436_ _1435_/A _1433_/X _1434_/X _1435_/Y vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__o31a_2
X_1505_ _1714_/Q _1479_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1714_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1298_ _1298_/A _1298_/B vssd1 vssd1 vccd1 vccd1 _1358_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1221_ _1220_/A _1220_/B _1220_/C vssd1 vssd1 vccd1 vccd1 _1222_/B sky130_fd_sc_hd__a21oi_1
X_1152_ _1152_/A _1282_/A vssd1 vssd1 vccd1 vccd1 _1511_/B sky130_fd_sc_hd__or2_1
X_1083_ _1083_/A _1083_/B vssd1 vssd1 vccd1 vccd1 _1085_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0936_ _1775_/Q _0941_/B _0941_/C _0941_/D vssd1 vssd1 vccd1 vccd1 _1065_/B sky130_fd_sc_hd__nand4b_4
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0867_ _0917_/A _0909_/A _0897_/A _0897_/B vssd1 vssd1 vccd1 vccd1 _0869_/B sky130_fd_sc_hd__or4b_4
X_1419_ _1743_/Q _1423_/A2 _1406_/X _1812_/Q _1418_/X vssd1 vssd1 vccd1 vccd1 _1419_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1770_ _1806_/CLK _1770_/D vssd1 vssd1 vccd1 vccd1 _1770_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _1212_/A _1204_/B vssd1 vssd1 vccd1 vccd1 _1737_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1135_ _1010_/A _0992_/A _1135_/S vssd1 vssd1 vccd1 vccd1 _1137_/B sky130_fd_sc_hd__mux2_1
X_1066_ _1823_/Q _1457_/A _1065_/X vssd1 vssd1 vccd1 vccd1 _1066_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0919_ _0919_/A _1373_/B vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1753_ _1808_/CLK _1753_/D vssd1 vssd1 vccd1 vccd1 _1753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1822_ _1830_/CLK _1822_/D vssd1 vssd1 vccd1 vccd1 _1822_/Q sky130_fd_sc_hd__dfxtp_1
X_1684_ _1824_/Q _1466_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1824_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1118_ _0960_/B _1123_/S vssd1 vssd1 vccd1 vccd1 _1119_/S sky130_fd_sc_hd__and2b_1
X_1049_ _1063_/A _1049_/B vssd1 vssd1 vccd1 vccd1 _1049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1805_ _1806_/CLK _1805_/D vssd1 vssd1 vccd1 vccd1 _1805_/Q sky130_fd_sc_hd__dfxtp_1
X_1736_ _1808_/CLK _1736_/D vssd1 vssd1 vccd1 vccd1 _1736_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1809_/Q _1413_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1809_/D sky130_fd_sc_hd__mux2_1
X_1598_ _1582_/Y _1593_/C _1597_/X vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__a21bo_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1452_ _1737_/Q _1372_/A _1369_/B _1745_/Q vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__a22o_1
X_1521_ _1748_/Q _1389_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1748_/D sky130_fd_sc_hd__mux2_1
X_1383_ _1746_/Q _1381_/C _1379_/X _1382_/X vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__a211o_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1719_ _1797_/CLK _1719_/D vssd1 vssd1 vccd1 vccd1 _1719_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ _0952_/A _1282_/B vssd1 vssd1 vccd1 vccd1 _0952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0883_ _0914_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _0970_/B sky130_fd_sc_hd__and2_1
X_1504_ _1713_/Q _1477_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1713_/D sky130_fd_sc_hd__mux2_1
X_1366_ _1366_/A _1366_/B _1366_/C _1365_/X vssd1 vssd1 vccd1 vccd1 _1367_/C sky130_fd_sc_hd__or4b_1
X_1435_ _1435_/A _1435_/B vssd1 vssd1 vccd1 vccd1 _1435_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1297_ _1297_/A _1297_/B _1296_/X vssd1 vssd1 vccd1 vccd1 _1352_/B sky130_fd_sc_hd__or3b_1
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1788_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1151_ _1152_/A _1282_/A vssd1 vssd1 vccd1 vccd1 _1151_/Y sky130_fd_sc_hd__nor2_1
X_1220_ _1220_/A _1220_/B _1220_/C vssd1 vssd1 vccd1 vccd1 _1228_/A sky130_fd_sc_hd__and3_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1082_ _0834_/Y _1781_/Q _1406_/B _1105_/B _1785_/Q vssd1 vssd1 vccd1 vccd1 _1082_/X
+ sky130_fd_sc_hd__a32o_1
X_0866_ _0927_/A _0909_/A vssd1 vssd1 vccd1 vccd1 _0926_/B sky130_fd_sc_hd__nor2_1
X_0935_ _0929_/Y _1515_/B _1346_/A _1518_/A vssd1 vssd1 vccd1 vccd1 _0941_/D sky130_fd_sc_hd__and4bb_2
X_1349_ _1349_/A _1349_/B vssd1 vssd1 vccd1 vccd1 _1353_/B sky130_fd_sc_hd__nor2_1
X_1418_ input6/X _1375_/A _1377_/C _1726_/Q vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1203_ _1203_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1204_/B sky130_fd_sc_hd__and2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1134_ _1091_/A _1092_/A _1131_/Y _1133_/X vssd1 vssd1 vccd1 vccd1 _1137_/A sky130_fd_sc_hd__o2bb2a_1
X_1065_ _1710_/Q _1065_/B _1065_/C vssd1 vssd1 vccd1 vccd1 _1065_/X sky130_fd_sc_hd__and3_1
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0849_ _0927_/A _1162_/A vssd1 vssd1 vccd1 vccd1 _0954_/B sky130_fd_sc_hd__nand2_2
X_0918_ _1373_/B vssd1 vssd1 vccd1 vccd1 _0918_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1752_ _1808_/CLK _1752_/D vssd1 vssd1 vccd1 vccd1 _1752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1821_ _1826_/CLK _1821_/D vssd1 vssd1 vccd1 vccd1 _1821_/Q sky130_fd_sc_hd__dfxtp_1
X_1683_ _1823_/Q _1458_/X _1690_/S vssd1 vssd1 vccd1 vccd1 _1823_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1117_ _1736_/Q _0950_/B _0974_/X input7/X vssd1 vssd1 vccd1 vccd1 _1123_/S sky130_fd_sc_hd__a22o_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1048_ _1048_/A _1048_/B vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__or2_4
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1666_ _1808_/Q _1411_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__mux2_1
X_1804_ _1804_/CLK _1804_/D vssd1 vssd1 vccd1 vccd1 _1804_/Q sky130_fd_sc_hd__dfxtp_1
X_1735_ _1808_/CLK _1735_/D vssd1 vssd1 vccd1 vccd1 _1735_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1652_/B _1641_/B _1641_/C _1589_/B _1655_/A vssd1 vssd1 vccd1 vccd1 _1597_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1520_ _1747_/Q _1386_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1747_/D sky130_fd_sc_hd__mux2_1
X_1451_ _1435_/A _0948_/B _1449_/X _1450_/X vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__o2bb2a_1
X_1382_ _1428_/B _1368_/Y _1410_/B1 _1730_/Q vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1649_ _1791_/Q _1648_/B _1645_/X _1648_/Y vssd1 vssd1 vccd1 vccd1 _1791_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1718_ _1788_/CLK _1718_/D vssd1 vssd1 vccd1 vccd1 _1718_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0951_ _1162_/A _1162_/C _1162_/B _0917_/A vssd1 vssd1 vccd1 vccd1 _1282_/B sky130_fd_sc_hd__or4bb_4
X_0882_ _0952_/A _1511_/A vssd1 vssd1 vccd1 vccd1 _0977_/A sky130_fd_sc_hd__nor2_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1503_ _1712_/Q _1472_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1712_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1365_ _0970_/A _0904_/B _1083_/B _0968_/A vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__a31o_1
X_1296_ _1344_/A _1655_/B _1636_/D _1626_/C vssd1 vssd1 vccd1 vccd1 _1296_/X sky130_fd_sc_hd__or4_1
X_1434_ _1740_/Q _0870_/X _1425_/Y _1723_/Q vssd1 vssd1 vccd1 vccd1 _1434_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _1150_/A _1150_/B vssd1 vssd1 vccd1 vccd1 _1721_/D sky130_fd_sc_hd__xnor2_1
X_1081_ _1754_/Q _1081_/B vssd1 vssd1 vccd1 vccd1 _1090_/A sky130_fd_sc_hd__nand2_1
X_0934_ _0926_/B _0926_/C _0933_/X _0926_/A _0850_/X vssd1 vssd1 vccd1 vccd1 _1515_/B
+ sky130_fd_sc_hd__a32o_1
X_0865_ _0932_/B _0925_/B vssd1 vssd1 vccd1 vccd1 _1518_/A sky130_fd_sc_hd__or2_4
X_1417_ _1742_/Q _1423_/A2 _1406_/X _1811_/Q _1416_/X vssd1 vssd1 vccd1 vccd1 _1417_/X
+ sky130_fd_sc_hd__a221o_1
X_1348_ _1696_/D _1348_/B _1348_/C _1318_/B vssd1 vssd1 vccd1 vccd1 _1349_/B sky130_fd_sc_hd__or4b_1
X_1279_ _1626_/B _1291_/A _1655_/C vssd1 vssd1 vccd1 vccd1 _1292_/B sky130_fd_sc_hd__and3_2
XFILLER_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1202_ _1203_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1212_/A sky130_fd_sc_hd__nor2_2
Xclkbuf_4_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1799_/CLK sky130_fd_sc_hd__clkbuf_8
X_1064_ _1730_/Q _0950_/B _0974_/X input1/X vssd1 vssd1 vccd1 vccd1 _1076_/S sky130_fd_sc_hd__a22oi_4
X_1133_ _0984_/A _1728_/D _1135_/S _1132_/Y vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__a31o_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0848_ _1701_/Q _0914_/A vssd1 vssd1 vccd1 vccd1 _0848_/Y sky130_fd_sc_hd__nand2b_1
X_0917_ _0917_/A _1162_/A _1162_/B _1162_/C vssd1 vssd1 vccd1 vccd1 _1373_/B sky130_fd_sc_hd__or4_4
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _1826_/CLK _1820_/D vssd1 vssd1 vccd1 vccd1 _1820_/Q sky130_fd_sc_hd__dfxtp_1
X_1751_ _1808_/CLK _1751_/D vssd1 vssd1 vccd1 vccd1 _1751_/Q sky130_fd_sc_hd__dfxtp_1
X_1682_ _1682_/A _1682_/B vssd1 vssd1 vccd1 vccd1 _1690_/S sky130_fd_sc_hd__and2_4
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1047_ _1010_/A _0992_/A _1047_/S vssd1 vssd1 vccd1 vccd1 _1048_/B sky130_fd_sc_hd__mux2_1
X_1116_ _1719_/Q _0957_/X _1114_/Y _1115_/X vssd1 vssd1 vccd1 vccd1 _1728_/D sky130_fd_sc_hd__a211o_4
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1803_ _1803_/CLK _1803_/D vssd1 vssd1 vccd1 vccd1 _1803_/Q sky130_fd_sc_hd__dfxtp_1
X_1596_ _1641_/C _1596_/B vssd1 vssd1 vccd1 vccd1 _1596_/Y sky130_fd_sc_hd__nor2_1
X_1665_ _1807_/Q _1408_/X _1666_/S vssd1 vssd1 vccd1 vccd1 _1807_/D sky130_fd_sc_hd__mux2_1
X_1734_ _1808_/CLK _1734_/D vssd1 vssd1 vccd1 vccd1 _1734_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1450_ _1744_/Q _1369_/B _1425_/Y _1727_/Q _1435_/A vssd1 vssd1 vccd1 vccd1 _1450_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ _1381_/A _1381_/B _1381_/C _1514_/B vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__or4_4
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1579_ _1579_/A _1648_/A _1579_/C vssd1 vssd1 vccd1 vccd1 _1602_/B sky130_fd_sc_hd__and3_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1648_ _1648_/A _1648_/B vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__nor2_1
X_1717_ _1830_/CLK _1717_/D vssd1 vssd1 vccd1 vccd1 _1717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0881_ _1698_/Q _1162_/C _0894_/A vssd1 vssd1 vccd1 vccd1 _1511_/A sky130_fd_sc_hd__or3_4
X_0950_ _1297_/A _0950_/B vssd1 vssd1 vccd1 vccd1 _0950_/X sky130_fd_sc_hd__or2_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1433_ _1732_/Q _1372_/A _1424_/X _1760_/Q vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__a22o_1
X_1502_ _1711_/Q _1466_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1711_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1364_ _1364_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1366_/C sky130_fd_sc_hd__nand2_1
X_1295_ _1359_/A _1295_/B vssd1 vssd1 vccd1 vccd1 _1297_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1080_ _0833_/Y _0834_/Y _1105_/B _1513_/C _1787_/Q vssd1 vssd1 vccd1 vccd1 _1081_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0933_ _0933_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__xor2_2
X_0864_ _0932_/B _0925_/B vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__nor2_8
X_1347_ _1347_/A _1352_/C _1360_/A _1347_/D vssd1 vssd1 vccd1 vccd1 _1348_/C sky130_fd_sc_hd__or4_1
X_1416_ input5/X _1375_/A _1377_/C _1725_/Q vssd1 vssd1 vccd1 vccd1 _1416_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1278_ _1650_/S _1655_/C vssd1 vssd1 vccd1 vccd1 _1278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1201_ _1737_/Q _1183_/Y _1200_/X vssd1 vssd1 vccd1 vccd1 _1203_/B sky130_fd_sc_hd__a21oi_2
X_1132_ _0982_/X _1135_/S _0903_/Y vssd1 vssd1 vccd1 vccd1 _1132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1063_ _1063_/A _1063_/B vssd1 vssd1 vccd1 vccd1 _1063_/X sky130_fd_sc_hd__or2_2
X_0916_ _1083_/A _0912_/B _1083_/B _1373_/A vssd1 vssd1 vccd1 vccd1 _0928_/A sky130_fd_sc_hd__o22ai_4
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0847_ _1624_/B vssd1 vssd1 vccd1 vccd1 _1803_/D sky130_fd_sc_hd__inv_2
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1750_ _1808_/CLK _1750_/D vssd1 vssd1 vccd1 vccd1 _1750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1681_ _1822_/Q _1498_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1822_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1115_ input8/X _0950_/X _1206_/A _1814_/Q vssd1 vssd1 vccd1 vccd1 _1115_/X sky130_fd_sc_hd__a22o_2
X_1046_ _1063_/A _1020_/X _1044_/Y _1045_/X vssd1 vssd1 vccd1 vccd1 _1048_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1797_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1802_ _1804_/CLK _1802_/D vssd1 vssd1 vccd1 vccd1 _1802_/Q sky130_fd_sc_hd__dfxtp_1
X_1733_ _1829_/CLK _1733_/D vssd1 vssd1 vccd1 vccd1 _1733_/Q sky130_fd_sc_hd__dfxtp_2
X_1595_ _1772_/Q _1577_/B _1695_/A vssd1 vssd1 vccd1 vccd1 _1772_/D sky130_fd_sc_hd__a21o_1
X_1664_ _0828_/Y _1559_/A _1663_/X vssd1 vssd1 vccd1 vccd1 _1806_/D sky130_fd_sc_hd__o21ai_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1029_ _1030_/B vssd1 vssd1 vccd1 vccd1 _1029_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1380_ _1381_/A _1381_/B _1381_/C _1514_/B vssd1 vssd1 vccd1 vccd1 _1380_/Y sky130_fd_sc_hd__nor4_4
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1716_ _1829_/CLK _1716_/D vssd1 vssd1 vccd1 vccd1 _1716_/Q sky130_fd_sc_hd__dfxtp_1
X_1578_ _1568_/B _1577_/Y _1695_/A vssd1 vssd1 vccd1 vccd1 _1770_/D sky130_fd_sc_hd__a21oi_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1647_ _1790_/Q _1643_/X _1650_/S vssd1 vssd1 vccd1 vccd1 _1790_/D sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0880_ _0952_/A _1084_/B vssd1 vssd1 vccd1 vccd1 _1513_/B sky130_fd_sc_hd__nor2_2
X_1363_ _1363_/A _1456_/B vssd1 vssd1 vccd1 vccd1 _1372_/C sky130_fd_sc_hd__nand2_1
X_1432_ _1445_/A _1052_/X _1430_/X _1431_/X vssd1 vssd1 vccd1 vccd1 _1432_/X sky130_fd_sc_hd__o22a_2
X_1501_ _1710_/Q _1458_/X _1508_/S vssd1 vssd1 vccd1 vccd1 _1710_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1294_ _1804_/D _1630_/B _1641_/C _1596_/B vssd1 vssd1 vccd1 vccd1 _1295_/B sky130_fd_sc_hd__or4_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0932_ _1298_/A _0932_/B vssd1 vssd1 vccd1 vccd1 _1282_/A sky130_fd_sc_hd__and2_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0863_ _1162_/A _1162_/B _1162_/C _0927_/A vssd1 vssd1 vccd1 vccd1 _0925_/B sky130_fd_sc_hd__or4b_4
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1346_ _1346_/A _1346_/B vssd1 vssd1 vccd1 vccd1 _1347_/D sky130_fd_sc_hd__nand2_1
X_1415_ _1741_/Q _1423_/A2 _1406_/X _1810_/Q _1414_/X vssd1 vssd1 vccd1 vccd1 _1415_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1277_ _1630_/B _1277_/B vssd1 vssd1 vccd1 vccd1 _1655_/C sky130_fd_sc_hd__nor2_4
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1200_ _1719_/Q _1173_/C _1206_/B _1753_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1200_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1062_ _1049_/Y _1060_/X _1061_/X vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__o21a_1
X_1131_ _1004_/A _1135_/S _1728_/D vssd1 vssd1 vccd1 vccd1 _1131_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0915_ _1298_/A _1083_/B vssd1 vssd1 vccd1 vccd1 _1374_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0846_ _1579_/A _1579_/C vssd1 vssd1 vccd1 vccd1 _1624_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ _1308_/A _1641_/D _1320_/X _1295_/B _1303_/B vssd1 vssd1 vccd1 vccd1 _1359_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _1821_/Q _1492_/X _1681_/S vssd1 vssd1 vccd1 vccd1 _1821_/D sky130_fd_sc_hd__mux2_1
X_1114_ _1114_/A _1114_/B vssd1 vssd1 vccd1 vccd1 _1114_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1045_ _1049_/B _1041_/Y _1091_/A vssd1 vssd1 vccd1 vccd1 _1045_/X sky130_fd_sc_hd__a21o_1
X_0829_ _1760_/Q vssd1 vssd1 vccd1 vccd1 _0829_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_6502_90 vssd1 vssd1 vccd1 vccd1 wrapped_6502_90/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1663_ _1806_/Q _1805_/Q _1805_/D vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__or3b_1
X_1801_ _1804_/CLK _1801_/D vssd1 vssd1 vccd1 vccd1 _1801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1732_ _1829_/CLK _1732_/D vssd1 vssd1 vccd1 vccd1 _1732_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _1771_/Q _1593_/X _1650_/S vssd1 vssd1 vccd1 vccd1 _1771_/D sky130_fd_sc_hd__mux2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1028_ _1010_/A _0992_/A _1028_/S vssd1 vssd1 vccd1 vccd1 _1030_/B sky130_fd_sc_hd__mux2_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1646_ _1643_/X _1644_/Y _1789_/Q _1650_/S vssd1 vssd1 vccd1 vccd1 _1789_/D sky130_fd_sc_hd__o2bb2a_1
X_1715_ _1829_/CLK _1715_/D vssd1 vssd1 vccd1 vccd1 _1715_/Q sky130_fd_sc_hd__dfxtp_1
X_1577_ _1770_/Q _1577_/B vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1500_ _1500_/A _1682_/B vssd1 vssd1 vccd1 vccd1 _1508_/S sky130_fd_sc_hd__and2_4
X_1293_ _1586_/A _1652_/B vssd1 vssd1 vccd1 vccd1 _1596_/B sky130_fd_sc_hd__or2_2
X_1362_ _0927_/A _1162_/A _0868_/A _0932_/B _1346_/A vssd1 vssd1 vccd1 vccd1 _1456_/B
+ sky130_fd_sc_hd__o41a_2
X_1431_ _1739_/Q _1369_/B _1425_/Y _1722_/Q _1435_/A vssd1 vssd1 vccd1 vccd1 _1431_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1629_ _1784_/Q _1624_/C _1628_/X _1759_/Q vssd1 vssd1 vccd1 vccd1 _1784_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0862_ _0914_/A _1701_/Q vssd1 vssd1 vccd1 vccd1 _0862_/Y sky130_fd_sc_hd__nand2b_2
X_0931_ _1166_/A _1083_/A vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__nor2_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1345_ _1345_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__nand2_1
X_1414_ input4/X _1375_/A _1377_/C _1724_/Q vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__a22o_1
X_1276_ _1586_/C _1630_/B vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1130_ _1737_/Q _0950_/B _0974_/X input8/X vssd1 vssd1 vccd1 vccd1 _1135_/S sky130_fd_sc_hd__a22o_2
X_1061_ _1010_/Y _0994_/A _1061_/S vssd1 vssd1 vccd1 vccd1 _1061_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0845_ input7/X _1768_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1579_/C sky130_fd_sc_hd__mux2_4
X_0914_ _0914_/A _0925_/B vssd1 vssd1 vccd1 vccd1 _1515_/A sky130_fd_sc_hd__nor2_1
X_1259_ _1628_/A _1652_/B _1586_/C _1626_/C vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__or4_1
X_1328_ _1327_/X _1328_/B _1328_/C vssd1 vssd1 vccd1 vccd1 _1333_/B sky130_fd_sc_hd__and3b_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1113_ _1830_/Q _1682_/A _1500_/A _1717_/Q _1112_/X vssd1 vssd1 vccd1 vccd1 _1114_/B
+ sky130_fd_sc_hd__a221oi_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1044_ _1047_/S _1043_/Y _1042_/X vssd1 vssd1 vccd1 vccd1 _1044_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0828_ _1806_/Q vssd1 vssd1 vccd1 vccd1 _0828_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_6502_91 vssd1 vssd1 vccd1 vccd1 wrapped_6502_91/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1800_ _1804_/CLK _1800_/D vssd1 vssd1 vccd1 vccd1 _1800_/Q sky130_fd_sc_hd__dfxtp_4
X_1662_ _1801_/Q _1359_/A _1297_/B _1624_/B vssd1 vssd1 vccd1 vccd1 _1801_/D sky130_fd_sc_hd__a22o_1
X_1731_ _1829_/CLK _1731_/D vssd1 vssd1 vccd1 vccd1 _1731_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1593_/A _1593_/B _1593_/C _1592_/X vssd1 vssd1 vccd1 vccd1 _1593_/X sky130_fd_sc_hd__or4b_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1027_ _1063_/A _1006_/B _1025_/X _1026_/X vssd1 vssd1 vccd1 vccd1 _1031_/S sky130_fd_sc_hd__o22a_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1576_ input8/X _1769_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1769_/D sky130_fd_sc_hd__mux2_1
X_1645_ _1628_/A _1624_/B _1626_/D _1643_/X vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__a31o_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1714_ _1829_/CLK _1714_/D vssd1 vssd1 vccd1 vccd1 _1714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1430_ _1731_/Q _1372_/A _1424_/X _1757_/Q vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__a22o_1
X_1292_ _1340_/A _1292_/B _1292_/C vssd1 vssd1 vccd1 vccd1 _1696_/D sky130_fd_sc_hd__or3_1
X_1361_ _1308_/X _1333_/B _1359_/A vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1559_ _1559_/A _1559_/B vssd1 vssd1 vccd1 vccd1 _1760_/D sky130_fd_sc_hd__or2_1
X_1628_ _1628_/A _1628_/B _1628_/C vssd1 vssd1 vccd1 vccd1 _1628_/X sky130_fd_sc_hd__and3_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0930_ _1373_/A _0954_/B _0953_/C vssd1 vssd1 vccd1 vccd1 _1346_/A sky130_fd_sc_hd__or3_4
X_0861_ _1373_/A _0970_/A vssd1 vssd1 vccd1 vccd1 _0861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1413_ _1740_/Q _1423_/A2 _1406_/X _1809_/Q _1412_/X vssd1 vssd1 vccd1 vccd1 _1413_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1344_ _1344_/A _1344_/B _1344_/C _1641_/B vssd1 vssd1 vccd1 vccd1 _1364_/B sky130_fd_sc_hd__or4_2
X_1275_ _1804_/D _1580_/A vssd1 vssd1 vccd1 vccd1 _1291_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ _0985_/Y _1058_/X _1059_/X _1063_/A vssd1 vssd1 vccd1 vccd1 _1060_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0913_ _0897_/A _0973_/B _0912_/X vssd1 vssd1 vccd1 vccd1 _1568_/B sky130_fd_sc_hd__o21a_2
X_0844_ _1655_/A vssd1 vssd1 vccd1 vccd1 _1802_/D sky130_fd_sc_hd__clkinv_4
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1327_ _1804_/D _1242_/X _1267_/B _1276_/Y vssd1 vssd1 vccd1 vccd1 _1327_/X sky130_fd_sc_hd__o31a_1
X_1258_ _1614_/B _1641_/B vssd1 vssd1 vccd1 vccd1 _1626_/C sky130_fd_sc_hd__nand2_2
X_1189_ _1734_/Q _1183_/Y _1188_/X vssd1 vssd1 vccd1 vccd1 _1191_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1112_ _1822_/Q _1050_/S _1052_/S _1111_/X vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__o211a_1
X_1043_ _1043_/A _1049_/B vssd1 vssd1 vccd1 vccd1 _1043_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ _1636_/D _1582_/Y _1588_/Y _1300_/A _1586_/X vssd1 vssd1 vccd1 vccd1 _1592_/X
+ sky130_fd_sc_hd__o221a_1
X_1661_ _1800_/Q _1549_/D _1292_/B _1624_/B vssd1 vssd1 vccd1 vccd1 _1800_/D sky130_fd_sc_hd__a22o_1
X_1730_ _1807_/CLK _1730_/D vssd1 vssd1 vccd1 vccd1 _1730_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1026_ _1020_/X _1022_/Y _1091_/A vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _1826_/CLK _1713_/D vssd1 vssd1 vccd1 vccd1 _1713_/Q sky130_fd_sc_hd__dfxtp_1
X_1575_ input7/X _1768_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1768_/D sky130_fd_sc_hd__mux2_1
X_1644_ _1648_/B _1644_/B vssd1 vssd1 vccd1 vccd1 _1644_/Y sky130_fd_sc_hd__nor2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1009_/A _1124_/A vssd1 vssd1 vccd1 vccd1 _1010_/A sky130_fd_sc_hd__or2_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1360_ _1360_/A _1360_/B _1360_/C _1360_/D vssd1 vssd1 vccd1 vccd1 _1700_/D sky130_fd_sc_hd__or4_1
X_1291_ _1291_/A _1655_/C vssd1 vssd1 vccd1 vccd1 _1328_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1558_ _1760_/Q _1557_/X _1558_/S vssd1 vssd1 vccd1 vccd1 _1559_/B sky130_fd_sc_hd__mux2_1
X_1627_ _1783_/Q _1653_/A _1626_/X vssd1 vssd1 vccd1 vccd1 _1783_/D sky130_fd_sc_hd__a21o_1
X_1489_ _1727_/Q _1489_/B vssd1 vssd1 vccd1 vccd1 _1489_/Y sky130_fd_sc_hd__nand2_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0860_ _0952_/A _0970_/A vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__or2_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1343_ _1359_/A _1320_/X _1557_/S vssd1 vssd1 vccd1 vccd1 _1352_/C sky130_fd_sc_hd__o21ai_1
X_1412_ input3/X _1375_/A _1377_/C _1723_/Q vssd1 vssd1 vccd1 vccd1 _1412_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1274_ _1628_/A _1630_/C vssd1 vssd1 vccd1 vccd1 _1274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0989_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0994_/A sky130_fd_sc_hd__inv_2
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ _1298_/A _0912_/B vssd1 vssd1 vccd1 vccd1 _0912_/X sky130_fd_sc_hd__or2_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0843_ _1256_/A _1583_/A vssd1 vssd1 vccd1 vccd1 _1586_/A sky130_fd_sc_hd__nand2_2
X_1326_ _1630_/B _1633_/B vssd1 vssd1 vccd1 vccd1 _1589_/A sky130_fd_sc_hd__or2_2
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1257_ _1614_/B _1257_/B vssd1 vssd1 vccd1 vccd1 _1630_/B sky130_fd_sc_hd__or2_4
X_1188_ _1725_/Q _1173_/C _1206_/B _1750_/Q _0957_/B vssd1 vssd1 vccd1 vccd1 _1188_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1111_ _1709_/Q _1673_/A vssd1 vssd1 vccd1 vccd1 _1111_/X sky130_fd_sc_hd__or2_1
X_1042_ _1049_/B _1041_/Y _0982_/X vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1309_ _1641_/D _1320_/C _1344_/A _1308_/A vssd1 vssd1 vccd1 vccd1 _1309_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_4_15_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1814_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ _1630_/C _1655_/C vssd1 vssd1 vccd1 vccd1 _1593_/C sky130_fd_sc_hd__and2_2
X_1660_ _1799_/Q _1648_/B _1644_/Y _1655_/X vssd1 vssd1 vccd1 vccd1 _1799_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1025_ _1020_/X _1024_/Y _1023_/Y vssd1 vssd1 vccd1 vccd1 _1025_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1789_ _1797_/CLK _1789_/D vssd1 vssd1 vccd1 vccd1 _1789_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _1643_/A _1643_/B _1643_/C _1643_/D vssd1 vssd1 vccd1 vccd1 _1643_/X sky130_fd_sc_hd__or4_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1712_ _1825_/CLK _1712_/D vssd1 vssd1 vccd1 vccd1 _1712_/Q sky130_fd_sc_hd__dfxtp_1
X_1574_ input6/X _1767_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1767_/D sky130_fd_sc_hd__mux2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1008_ _0966_/Y _1007_/X _1063_/A vssd1 vssd1 vccd1 vccd1 _1012_/A sky130_fd_sc_hd__mux2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1290_ _1356_/B _1290_/B _1290_/C _1288_/X vssd1 vssd1 vccd1 vccd1 _1292_/C sky130_fd_sc_hd__or4b_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1628_/A _1626_/B _1626_/C _1626_/D vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__and4_1
X_1557_ input3/X _1554_/X _1557_/S vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__mux2_1
X_1488_ _1727_/Q _1489_/B vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__or2_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1342_ _1359_/A _1342_/B vssd1 vssd1 vccd1 vccd1 _1348_/B sky130_fd_sc_hd__nor2_1
X_1273_ _1352_/A _1358_/B _1273_/C vssd1 vssd1 vccd1 vccd1 _1340_/A sky130_fd_sc_hd__or3_1
X_1411_ _1739_/Q _1381_/X _1410_/X vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0988_ _1790_/Q _1513_/C _1406_/C _1756_/Q _0878_/A vssd1 vssd1 vccd1 vccd1 _0992_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1609_ _1802_/D _1652_/B _1589_/Y _1608_/X vssd1 vssd1 vccd1 vccd1 _1609_/X sky130_fd_sc_hd__a31o_1
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0842_ input6/X _1767_/Q _1770_/Q vssd1 vssd1 vccd1 vccd1 _1583_/A sky130_fd_sc_hd__mux2_2
X_0911_ _1369_/A _1512_/A _1554_/S _1356_/B vssd1 vssd1 vccd1 vccd1 _0973_/D sky130_fd_sc_hd__nor4_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1256_ _1256_/A _1256_/B vssd1 vssd1 vccd1 vccd1 _1641_/B sky130_fd_sc_hd__nand2_8
X_1325_ _1641_/C _1320_/B _1321_/X _1324_/X vssd1 vssd1 vccd1 vccd1 _1342_/B sky130_fd_sc_hd__o31a_1
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1187_ _1187_/A _1187_/B vssd1 vssd1 vccd1 vccd1 _1733_/D sky130_fd_sc_hd__xor2_1
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1014_/A _1240_/A _1109_/Y _1128_/A vssd1 vssd1 vccd1 vccd1 _1144_/A sky130_fd_sc_hd__o211ai_4
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1041_ _1041_/A _1047_/S vssd1 vssd1 vccd1 vccd1 _1041_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1308_ _1308_/A _1320_/C vssd1 vssd1 vccd1 vccd1 _1308_/X sky130_fd_sc_hd__or2_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1239_ _1239_/A _1239_/B _1239_/C vssd1 vssd1 vccd1 vccd1 _1240_/B sky130_fd_sc_hd__and3_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1274_/Y _1588_/Y _1589_/A vssd1 vssd1 vccd1 vccd1 _1593_/B sky130_fd_sc_hd__a21oi_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1024_ _1024_/A _1028_/S vssd1 vssd1 vccd1 vccd1 _1024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1788_ _1788_/CLK _1788_/D vssd1 vssd1 vccd1 vccd1 _1788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 _1559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1642_ _1630_/C _1655_/C _1583_/Y _1633_/Y vssd1 vssd1 vccd1 vccd1 _1643_/D sky130_fd_sc_hd__a31o_1
Xclkbuf_4_14_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1808_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1711_ _1825_/CLK _1711_/D vssd1 vssd1 vccd1 vccd1 _1711_/Q sky130_fd_sc_hd__dfxtp_1
X_1573_ input5/X _1766_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1766_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ _1006_/B _1004_/Y _1005_/Y _1006_/X vssd1 vssd1 vccd1 vccd1 _1007_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1556_ _1554_/S _1510_/B _1542_/S _1555_/X vssd1 vssd1 vccd1 vccd1 _1558_/S sky130_fd_sc_hd__o31a_1
X_1625_ _1782_/Q _1624_/C _1628_/B _1628_/C vssd1 vssd1 vccd1 vccd1 _1782_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1707_/Q _1486_/X _1499_/S vssd1 vssd1 vccd1 vccd1 _1707_/D sky130_fd_sc_hd__mux2_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1410_ _1722_/Q _1377_/C _1410_/B1 _1409_/X vssd1 vssd1 vccd1 vccd1 _1410_/X sky130_fd_sc_hd__a211o_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1341_ _1341_/A _1349_/A _1341_/C vssd1 vssd1 vccd1 vccd1 _1698_/D sky130_fd_sc_hd__or3_1
X_1272_ _1359_/A _1328_/C vssd1 vssd1 vccd1 vccd1 _1273_/C sky130_fd_sc_hd__nor2_1
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0987_ _1063_/A _0979_/X _0986_/X _0960_/Y vssd1 vssd1 vccd1 vccd1 _0996_/B sky130_fd_sc_hd__a31o_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1608_ _1582_/Y _1606_/X _1607_/Y _1653_/A vssd1 vssd1 vccd1 vccd1 _1608_/X sky130_fd_sc_hd__a31o_1
X_1539_ _1725_/Q _1726_/Q _1727_/Q _1719_/Q vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__or4_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0910_ _0927_/A _1351_/A vssd1 vssd1 vccd1 vccd1 _1356_/B sky130_fd_sc_hd__and2b_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0841_ _1628_/A vssd1 vssd1 vccd1 vccd1 _1804_/D sky130_fd_sc_hd__clkinv_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1255_ _1256_/A _1256_/B vssd1 vssd1 vccd1 vccd1 _1257_/B sky130_fd_sc_hd__and2_1
X_1324_ _1636_/D _1633_/B _1320_/B _1655_/B vssd1 vssd1 vccd1 vccd1 _1324_/X sky130_fd_sc_hd__a211o_1
X_1186_ _1187_/A _1187_/B vssd1 vssd1 vccd1 vccd1 _1191_/A sky130_fd_sc_hd__or2_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ _1732_/Q _0950_/B _0974_/X input3/X vssd1 vssd1 vccd1 vccd1 _1047_/S sky130_fd_sc_hd__a22o_2
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1238_ _1238_/A _1238_/B vssd1 vssd1 vccd1 vccd1 _1745_/D sky130_fd_sc_hd__xnor2_1
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1307_ _1653_/B _1596_/B vssd1 vssd1 vccd1 vccd1 _1320_/C sky130_fd_sc_hd__or2_2
X_1169_ _1170_/A _1170_/B vssd1 vssd1 vccd1 vccd1 _1181_/B sky130_fd_sc_hd__or2_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1023_ _1020_/X _1022_/Y _0982_/X vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1787_ _1804_/CLK _1787_/D vssd1 vssd1 vccd1 vccd1 _1787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1572_ input4/X _1765_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1765_/D sky130_fd_sc_hd__mux2_1
X_1641_ _1655_/A _1641_/B _1641_/C _1641_/D vssd1 vssd1 vccd1 vccd1 _1643_/C sky130_fd_sc_hd__nor4_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1710_ _1830_/CLK _1710_/D vssd1 vssd1 vccd1 vccd1 _1710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ _1043_/A _1006_/B _1011_/S vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__or3b_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1555_ _1795_/Q _1794_/Q _1084_/B _0868_/A _1801_/Q vssd1 vssd1 vccd1 vccd1 _1555_/X
+ sky130_fd_sc_hd__o32a_1
X_1624_ _1655_/A _1624_/B _1624_/C vssd1 vssd1 vccd1 vccd1 _1628_/C sky130_fd_sc_hd__nor3_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1486_ input6/X _1479_/S _1485_/X vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__a21bo_2
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _1806_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ _1340_/A _1340_/B _1347_/A _1340_/D vssd1 vssd1 vccd1 vccd1 _1341_/C sky130_fd_sc_hd__or4_1
X_1271_ _1308_/A _1580_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _1328_/C sky130_fd_sc_hd__or3_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0986_ _0982_/X _0984_/Y _0986_/S vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__mux2_1
X_1607_ _1803_/D _1652_/B _1641_/C vssd1 vssd1 vccd1 vccd1 _1607_/Y sky130_fd_sc_hd__a21oi_1
X_1538_ _1560_/A _1542_/S _1510_/A vssd1 vssd1 vccd1 vccd1 _1543_/S sky130_fd_sc_hd__o21ba_1
X_1469_ _1723_/Q _1469_/B vssd1 vssd1 vccd1 vccd1 _1469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0840_ _1256_/A _1648_/A vssd1 vssd1 vccd1 vccd1 _1628_/A sky130_fd_sc_hd__nand2_8
X_1323_ _1586_/C _1323_/B vssd1 vssd1 vccd1 vccd1 _1633_/B sky130_fd_sc_hd__or2_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1254_ _1586_/C _1323_/B vssd1 vssd1 vccd1 vccd1 _1636_/D sky130_fd_sc_hd__nand2_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1185_ _1733_/Q _1183_/Y _1184_/X vssd1 vssd1 vccd1 vccd1 _1187_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0969_ _0914_/A _1282_/B _1345_/A vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1306_ _1596_/B _1644_/B vssd1 vssd1 vccd1 vccd1 _1641_/D sky130_fd_sc_hd__or2_4
X_1237_ input8/X _1156_/B _1205_/Y _1745_/Q _1236_/X vssd1 vssd1 vccd1 vccd1 _1238_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1168_ _0914_/A _1152_/A _1163_/Y _1167_/X vssd1 vssd1 vccd1 vccd1 _1170_/B sky130_fd_sc_hd__o211a_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1099_ _1102_/A _1102_/B _1098_/A vssd1 vssd1 vccd1 vccd1 _1100_/B sky130_fd_sc_hd__o21a_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1022_ _1041_/A _1028_/S vssd1 vssd1 vccd1 vccd1 _1022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1786_ _1797_/CLK _1786_/D vssd1 vssd1 vccd1 vccd1 _1786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1571_ input3/X _1764_/Q _1576_/S vssd1 vssd1 vccd1 vccd1 _1764_/D sky130_fd_sc_hd__mux2_1
X_1640_ _1628_/B _1580_/Y _1639_/X _1602_/B vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__o31a_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1005_ _1006_/B _1004_/Y _0982_/X vssd1 vssd1 vccd1 vccd1 _1005_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1769_ _1769_/CLK _1769_/D vssd1 vssd1 vccd1 vccd1 _1769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput30 _1423_/X vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_4
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1554_ _1723_/Q _0832_/Y _1554_/S vssd1 vssd1 vccd1 vccd1 _1554_/X sky130_fd_sc_hd__mux2_1
X_1623_ _1781_/Q _1648_/B _1602_/X _1622_/X vssd1 vssd1 vccd1 vccd1 _1781_/D sky130_fd_sc_hd__a22o_1
X_1485_ _1485_/A _1485_/B _1484_/X vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__or3b_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

