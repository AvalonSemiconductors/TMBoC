magic
tech sky130B
magscale 1 2
timestamp 1680210569
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 198 756 68816 67584
<< metal2 >>
rect 3514 0 3570 800
rect 10506 0 10562 800
rect 17498 0 17554 800
rect 24490 0 24546 800
rect 31482 0 31538 800
rect 38474 0 38530 800
rect 45466 0 45522 800
rect 52458 0 52514 800
rect 59450 0 59506 800
rect 66442 0 66498 800
<< obsm2 >>
rect 202 856 68152 67969
rect 202 750 3458 856
rect 3626 750 10450 856
rect 10618 750 17442 856
rect 17610 750 24434 856
rect 24602 750 31426 856
rect 31594 750 38418 856
rect 38586 750 45410 856
rect 45578 750 52402 856
rect 52570 750 59394 856
rect 59562 750 66386 856
rect 66554 750 68152 856
<< metal3 >>
rect 0 67872 800 67992
rect 0 65424 800 65544
rect 0 62976 800 63096
rect 0 60528 800 60648
rect 0 58080 800 58200
rect 0 55632 800 55752
rect 0 53184 800 53304
rect 0 50736 800 50856
rect 0 48288 800 48408
rect 0 45840 800 45960
rect 0 43392 800 43512
rect 0 40944 800 41064
rect 0 38496 800 38616
rect 0 36048 800 36168
rect 0 33600 800 33720
rect 0 31152 800 31272
rect 0 28704 800 28824
rect 0 26256 800 26376
rect 0 23808 800 23928
rect 0 21360 800 21480
rect 0 18912 800 19032
rect 0 16464 800 16584
rect 0 14016 800 14136
rect 0 11568 800 11688
rect 0 9120 800 9240
rect 0 6672 800 6792
rect 0 4224 800 4344
rect 0 1776 800 1896
<< obsm3 >>
rect 880 67792 67607 67965
rect 197 65624 67607 67792
rect 880 65344 67607 65624
rect 197 63176 67607 65344
rect 880 62896 67607 63176
rect 197 60728 67607 62896
rect 880 60448 67607 60728
rect 197 58280 67607 60448
rect 880 58000 67607 58280
rect 197 55832 67607 58000
rect 880 55552 67607 55832
rect 197 53384 67607 55552
rect 880 53104 67607 53384
rect 197 50936 67607 53104
rect 880 50656 67607 50936
rect 197 48488 67607 50656
rect 880 48208 67607 48488
rect 197 46040 67607 48208
rect 880 45760 67607 46040
rect 197 43592 67607 45760
rect 880 43312 67607 43592
rect 197 41144 67607 43312
rect 880 40864 67607 41144
rect 197 38696 67607 40864
rect 880 38416 67607 38696
rect 197 36248 67607 38416
rect 880 35968 67607 36248
rect 197 33800 67607 35968
rect 880 33520 67607 33800
rect 197 31352 67607 33520
rect 880 31072 67607 31352
rect 197 28904 67607 31072
rect 880 28624 67607 28904
rect 197 26456 67607 28624
rect 880 26176 67607 26456
rect 197 24008 67607 26176
rect 880 23728 67607 24008
rect 197 21560 67607 23728
rect 880 21280 67607 21560
rect 197 19112 67607 21280
rect 880 18832 67607 19112
rect 197 16664 67607 18832
rect 880 16384 67607 16664
rect 197 14216 67607 16384
rect 880 13936 67607 14216
rect 197 11768 67607 13936
rect 880 11488 67607 11768
rect 197 9320 67607 11488
rect 880 9040 67607 9320
rect 197 6872 67607 9040
rect 880 6592 67607 6872
rect 197 4424 67607 6592
rect 880 4144 67607 4424
rect 197 1976 67607 4144
rect 880 1696 67607 1976
rect 197 987 67607 1696
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 611 2048 4128 66333
rect 4608 2048 19488 66333
rect 19968 2048 34848 66333
rect 35328 2048 50208 66333
rect 50688 2048 59557 66333
rect 611 987 59557 2048
<< labels >>
rlabel metal2 s 59450 0 59506 800 6 clk
port 1 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 io_oeb
port 10 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 io_out[10]
port 12 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 io_out[11]
port 13 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 io_out[12]
port 14 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 io_out[13]
port 15 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[14]
port 16 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_out[15]
port 17 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_out[16]
port 18 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_out[17]
port 19 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_out[18]
port 20 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_out[19]
port 21 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[1]
port 22 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 io_out[20]
port 23 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 io_out[21]
port 24 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_out[22]
port 25 nsew signal output
rlabel metal3 s 0 58080 800 58200 6 io_out[23]
port 26 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 io_out[24]
port 27 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 io_out[25]
port 28 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 io_out[26]
port 29 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_out[2]
port 30 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_out[3]
port 31 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[4]
port 32 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_out[5]
port 33 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 io_out[6]
port 34 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 io_out[7]
port 35 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[8]
port 36 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_out[9]
port 37 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 rst
port 38 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16171546
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS2650/runs/23_03_30_22_54/results/signoff/wrapped_as2650.magic.gds
string GDS_START 1393958
<< end >>

