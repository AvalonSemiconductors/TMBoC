magic
tech sky130B
magscale 1 2
timestamp 1680007425
<< viali >>
rect 15117 17221 15151 17255
rect 10609 17153 10643 17187
rect 15301 17017 15335 17051
rect 10701 16949 10735 16983
rect 11437 16609 11471 16643
rect 11713 16541 11747 16575
rect 14565 16541 14599 16575
rect 15025 16541 15059 16575
rect 15853 16541 15887 16575
rect 9689 16473 9723 16507
rect 14473 16405 14507 16439
rect 15117 16405 15151 16439
rect 15761 16405 15795 16439
rect 9137 16201 9171 16235
rect 11069 16201 11103 16235
rect 13461 16133 13495 16167
rect 15209 16133 15243 16167
rect 8585 16065 8619 16099
rect 9045 16065 9079 16099
rect 9873 16065 9907 16099
rect 10517 16065 10551 16099
rect 11161 16065 11195 16099
rect 12173 16065 12207 16099
rect 13001 16065 13035 16099
rect 15485 16065 15519 16099
rect 16129 16065 16163 16099
rect 8493 15861 8527 15895
rect 9781 15861 9815 15895
rect 10425 15861 10459 15895
rect 12265 15861 12299 15895
rect 12909 15861 12943 15895
rect 16037 15861 16071 15895
rect 9137 15521 9171 15555
rect 11161 15521 11195 15555
rect 11713 15521 11747 15555
rect 13461 15521 13495 15555
rect 13737 15521 13771 15555
rect 14565 15521 14599 15555
rect 16313 15521 16347 15555
rect 7941 15453 7975 15487
rect 8401 15453 8435 15487
rect 14289 15453 14323 15487
rect 7849 15385 7883 15419
rect 9413 15385 9447 15419
rect 8493 15317 8527 15351
rect 12725 15113 12759 15147
rect 14105 15113 14139 15147
rect 15669 15113 15703 15147
rect 8585 14977 8619 15011
rect 12817 14977 12851 15011
rect 14197 14977 14231 15011
rect 14933 14977 14967 15011
rect 15577 14977 15611 15011
rect 8861 14909 8895 14943
rect 10609 14909 10643 14943
rect 15117 14909 15151 14943
rect 14749 14841 14783 14875
rect 9873 14365 9907 14399
rect 14473 14365 14507 14399
rect 15117 14365 15151 14399
rect 9965 14229 9999 14263
rect 14381 14229 14415 14263
rect 15025 14229 15059 14263
rect 9413 14025 9447 14059
rect 13921 13957 13955 13991
rect 15669 13957 15703 13991
rect 9505 13889 9539 13923
rect 10977 13889 11011 13923
rect 13645 13821 13679 13855
rect 10885 13685 10919 13719
rect 13645 13481 13679 13515
rect 9965 13345 9999 13379
rect 7389 13277 7423 13311
rect 13737 13277 13771 13311
rect 14657 13277 14691 13311
rect 10241 13209 10275 13243
rect 11989 13209 12023 13243
rect 7297 13141 7331 13175
rect 14565 13141 14599 13175
rect 11805 12937 11839 12971
rect 7358 12869 7392 12903
rect 7113 12801 7147 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 14473 12801 14507 12835
rect 14933 12801 14967 12835
rect 15577 12801 15611 12835
rect 8493 12597 8527 12631
rect 11069 12597 11103 12631
rect 14381 12597 14415 12631
rect 15025 12597 15059 12631
rect 15669 12597 15703 12631
rect 11897 12393 11931 12427
rect 14565 12257 14599 12291
rect 16313 12257 16347 12291
rect 4721 12189 4755 12223
rect 5917 12189 5951 12223
rect 6009 12189 6043 12223
rect 6561 12189 6595 12223
rect 9321 12189 9355 12223
rect 13553 12189 13587 12223
rect 13645 12189 13679 12223
rect 14289 12189 14323 12223
rect 6837 12121 6871 12155
rect 8585 12121 8619 12155
rect 10425 12121 10459 12155
rect 4629 12053 4663 12087
rect 9229 12053 9263 12087
rect 6009 11849 6043 11883
rect 9873 11849 9907 11883
rect 5641 11781 5675 11815
rect 5857 11781 5891 11815
rect 11161 11781 11195 11815
rect 15117 11781 15151 11815
rect 4270 11713 4304 11747
rect 4537 11713 4571 11747
rect 8677 11713 8711 11747
rect 8401 11645 8435 11679
rect 13369 11645 13403 11679
rect 15393 11645 15427 11679
rect 3157 11509 3191 11543
rect 5825 11509 5859 11543
rect 6929 11509 6963 11543
rect 6377 11305 6411 11339
rect 8033 11237 8067 11271
rect 10057 11237 10091 11271
rect 7297 11169 7331 11203
rect 10885 11169 10919 11203
rect 12633 11169 12667 11203
rect 3157 11101 3191 11135
rect 3341 11101 3375 11135
rect 5825 11101 5859 11135
rect 6285 11101 6319 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7849 11101 7883 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 9413 11101 9447 11135
rect 9965 11101 9999 11135
rect 3433 11033 3467 11067
rect 5549 11033 5583 11067
rect 11161 11033 11195 11067
rect 4077 10965 4111 10999
rect 9229 10965 9263 10999
rect 7021 10761 7055 10795
rect 7665 10761 7699 10795
rect 11897 10761 11931 10795
rect 2329 10625 2363 10659
rect 7113 10625 7147 10659
rect 10977 10625 11011 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 2237 10557 2271 10591
rect 2789 10557 2823 10591
rect 3065 10557 3099 10591
rect 9137 10557 9171 10591
rect 9413 10557 9447 10591
rect 4537 10421 4571 10455
rect 11069 10421 11103 10455
rect 2697 10217 2731 10251
rect 3341 10217 3375 10251
rect 13185 10217 13219 10251
rect 4077 10149 4111 10183
rect 2789 10013 2823 10047
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 7757 10013 7791 10047
rect 7941 10013 7975 10047
rect 10517 10013 10551 10047
rect 11161 10013 11195 10047
rect 11253 10013 11287 10047
rect 11805 10013 11839 10047
rect 12081 10013 12115 10047
rect 7573 9945 7607 9979
rect 7665 9945 7699 9979
rect 10609 9877 10643 9911
rect 11069 9605 11103 9639
rect 11989 9605 12023 9639
rect 7113 9537 7147 9571
rect 7665 9537 7699 9571
rect 8125 9537 8159 9571
rect 10977 9537 11011 9571
rect 11713 9537 11747 9571
rect 2605 9469 2639 9503
rect 2881 9469 2915 9503
rect 8401 9469 8435 9503
rect 8493 9401 8527 9435
rect 4353 9333 4387 9367
rect 13461 9333 13495 9367
rect 2697 9129 2731 9163
rect 3341 9129 3375 9163
rect 3985 9129 4019 9163
rect 5917 9129 5951 9163
rect 13001 9129 13035 9163
rect 13553 9061 13587 9095
rect 14565 9061 14599 9095
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 5825 8925 5859 8959
rect 6009 8925 6043 8959
rect 7389 8925 7423 8959
rect 9873 8925 9907 8959
rect 10793 8925 10827 8959
rect 13185 8925 13219 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 4537 8857 4571 8891
rect 6929 8857 6963 8891
rect 7021 8857 7055 8891
rect 7757 8857 7791 8891
rect 4353 8789 4387 8823
rect 6653 8789 6687 8823
rect 7941 8789 7975 8823
rect 9781 8789 9815 8823
rect 12081 8789 12115 8823
rect 13277 8789 13311 8823
rect 5089 8585 5123 8619
rect 6745 8585 6779 8619
rect 7849 8585 7883 8619
rect 11805 8585 11839 8619
rect 7481 8517 7515 8551
rect 9413 8517 9447 8551
rect 11161 8517 11195 8551
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 7021 8449 7055 8483
rect 7113 8449 7147 8483
rect 14013 8449 14047 8483
rect 2513 8381 2547 8415
rect 2789 8381 2823 8415
rect 4537 8381 4571 8415
rect 9137 8381 9171 8415
rect 13277 8381 13311 8415
rect 13553 8381 13587 8415
rect 14105 8381 14139 8415
rect 8033 8313 8067 8347
rect 2513 8041 2547 8075
rect 3157 8041 3191 8075
rect 9137 8041 9171 8075
rect 12725 7973 12759 8007
rect 3985 7905 4019 7939
rect 9689 7905 9723 7939
rect 16313 7905 16347 7939
rect 2605 7837 2639 7871
rect 3249 7837 3283 7871
rect 4169 7837 4203 7871
rect 4353 7837 4387 7871
rect 9321 7837 9355 7871
rect 10425 7837 10459 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 7021 7769 7055 7803
rect 12173 7769 12207 7803
rect 14289 7769 14323 7803
rect 16037 7769 16071 7803
rect 5733 7701 5767 7735
rect 9505 7701 9539 7735
rect 5089 7497 5123 7531
rect 7021 7497 7055 7531
rect 8309 7497 8343 7531
rect 10425 7497 10459 7531
rect 11989 7497 12023 7531
rect 15301 7497 15335 7531
rect 15945 7497 15979 7531
rect 9597 7429 9631 7463
rect 10425 7361 10459 7395
rect 10701 7361 10735 7395
rect 11897 7361 11931 7395
rect 14289 7361 14323 7395
rect 15393 7361 15427 7395
rect 15853 7361 15887 7395
rect 4905 7293 4939 7327
rect 4997 7293 5031 7327
rect 6653 7225 6687 7259
rect 7205 7225 7239 7259
rect 5457 7157 5491 7191
rect 7021 7157 7055 7191
rect 14197 7157 14231 7191
rect 11989 6817 12023 6851
rect 14289 6817 14323 6851
rect 4169 6749 4203 6783
rect 4813 6749 4847 6783
rect 7021 6749 7055 6783
rect 7849 6749 7883 6783
rect 8222 6749 8256 6783
rect 9505 6749 9539 6783
rect 9597 6749 9631 6783
rect 10425 6749 10459 6783
rect 4721 6681 4755 6715
rect 8033 6681 8067 6715
rect 8125 6681 8159 6715
rect 14565 6681 14599 6715
rect 4077 6613 4111 6647
rect 5733 6613 5767 6647
rect 8409 6613 8443 6647
rect 16037 6613 16071 6647
rect 4813 6409 4847 6443
rect 7573 6409 7607 6443
rect 14197 6409 14231 6443
rect 15577 6409 15611 6443
rect 3341 6341 3375 6375
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 10609 6273 10643 6307
rect 11897 6273 11931 6307
rect 14105 6273 14139 6307
rect 15485 6273 15519 6307
rect 3065 6205 3099 6239
rect 8217 6205 8251 6239
rect 9689 6205 9723 6239
rect 9965 6205 9999 6239
rect 10517 6205 10551 6239
rect 11805 6069 11839 6103
rect 5733 5865 5767 5899
rect 8493 5865 8527 5899
rect 9229 5865 9263 5899
rect 12633 5865 12667 5899
rect 3341 5797 3375 5831
rect 3985 5729 4019 5763
rect 11161 5729 11195 5763
rect 2605 5661 2639 5695
rect 3065 5661 3099 5695
rect 3341 5661 3375 5695
rect 7941 5661 7975 5695
rect 8401 5661 8435 5695
rect 9321 5661 9355 5695
rect 10885 5661 10919 5695
rect 13369 5661 13403 5695
rect 16037 5661 16071 5695
rect 2513 5593 2547 5627
rect 4261 5593 4295 5627
rect 7849 5525 7883 5559
rect 13277 5525 13311 5559
rect 15945 5525 15979 5559
rect 3433 5321 3467 5355
rect 4813 5321 4847 5355
rect 11069 5321 11103 5355
rect 12173 5321 12207 5355
rect 3525 5253 3559 5287
rect 2513 5185 2547 5219
rect 3341 5185 3375 5219
rect 4537 5185 4571 5219
rect 4813 5185 4847 5219
rect 8125 5185 8159 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 11161 5185 11195 5219
rect 12265 5185 12299 5219
rect 12909 5185 12943 5219
rect 13921 5185 13955 5219
rect 14749 5185 14783 5219
rect 14933 5185 14967 5219
rect 16957 5185 16991 5219
rect 17877 5185 17911 5219
rect 3157 5117 3191 5151
rect 8861 5117 8895 5151
rect 15853 5117 15887 5151
rect 18153 5117 18187 5151
rect 7941 5049 7975 5083
rect 16221 5049 16255 5083
rect 16313 5049 16347 5083
rect 2605 4981 2639 5015
rect 3709 4981 3743 5015
rect 12817 4981 12851 5015
rect 14013 4981 14047 5015
rect 14565 4981 14599 5015
rect 17049 4981 17083 5015
rect 2513 4777 2547 4811
rect 11437 4777 11471 4811
rect 9137 4709 9171 4743
rect 15209 4709 15243 4743
rect 17141 4709 17175 4743
rect 7297 4641 7331 4675
rect 13185 4641 13219 4675
rect 14841 4641 14875 4675
rect 15761 4641 15795 4675
rect 1961 4573 1995 4607
rect 2421 4573 2455 4607
rect 3065 4573 3099 4607
rect 3341 4573 3375 4607
rect 4169 4573 4203 4607
rect 4261 4573 4295 4607
rect 7389 4573 7423 4607
rect 8033 4573 8067 4607
rect 8309 4573 8343 4607
rect 9413 4573 9447 4607
rect 17601 4573 17635 4607
rect 9137 4505 9171 4539
rect 12909 4505 12943 4539
rect 16028 4505 16062 4539
rect 17877 4505 17911 4539
rect 1869 4437 1903 4471
rect 3341 4437 3375 4471
rect 4077 4437 4111 4471
rect 7849 4437 7883 4471
rect 8217 4437 8251 4471
rect 9321 4437 9355 4471
rect 15301 4437 15335 4471
rect 8769 4233 8803 4267
rect 13461 4233 13495 4267
rect 16313 4233 16347 4267
rect 9505 4165 9539 4199
rect 15853 4165 15887 4199
rect 17110 4165 17144 4199
rect 2421 4097 2455 4131
rect 4445 4097 4479 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 7849 4097 7883 4131
rect 8585 4097 8619 4131
rect 8861 4097 8895 4131
rect 9689 4097 9723 4131
rect 10149 4097 10183 4131
rect 10333 4097 10367 4131
rect 12633 4097 12667 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13369 4097 13403 4131
rect 14013 4097 14047 4131
rect 14280 4097 14314 4131
rect 16865 4097 16899 4131
rect 2697 4029 2731 4063
rect 7665 3961 7699 3995
rect 10149 3961 10183 3995
rect 16221 3961 16255 3995
rect 6837 3893 6871 3927
rect 7389 3893 7423 3927
rect 8401 3893 8435 3927
rect 9413 3893 9447 3927
rect 15393 3893 15427 3927
rect 18245 3893 18279 3927
rect 3065 3689 3099 3723
rect 4077 3689 4111 3723
rect 6377 3689 6411 3723
rect 7205 3689 7239 3723
rect 9229 3689 9263 3723
rect 12725 3689 12759 3723
rect 16773 3689 16807 3723
rect 7297 3553 7331 3587
rect 17417 3553 17451 3587
rect 3157 3485 3191 3519
rect 5190 3485 5224 3519
rect 5457 3485 5491 3519
rect 6193 3485 6227 3519
rect 6377 3485 6411 3519
rect 7021 3485 7055 3519
rect 8033 3485 8067 3519
rect 8125 3485 8159 3519
rect 8217 3485 8251 3519
rect 8401 3485 8435 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 10701 3485 10735 3519
rect 10793 3485 10827 3519
rect 11345 3485 11379 3519
rect 14289 3485 14323 3519
rect 14381 3485 14415 3519
rect 14933 3485 14967 3519
rect 15200 3485 15234 3519
rect 11590 3417 11624 3451
rect 17141 3417 17175 3451
rect 6837 3349 6871 3383
rect 7757 3349 7791 3383
rect 9597 3349 9631 3383
rect 16313 3349 16347 3383
rect 17233 3349 17267 3383
rect 4445 3145 4479 3179
rect 5549 3145 5583 3179
rect 15209 3145 15243 3179
rect 16865 3145 16899 3179
rect 17233 3145 17267 3179
rect 2973 3077 3007 3111
rect 15577 3077 15611 3111
rect 17325 3077 17359 3111
rect 2697 3009 2731 3043
rect 5641 3009 5675 3043
rect 6929 3009 6963 3043
rect 7757 3009 7791 3043
rect 8677 3009 8711 3043
rect 6653 2941 6687 2975
rect 6837 2941 6871 2975
rect 7849 2941 7883 2975
rect 8401 2941 8435 2975
rect 8493 2941 8527 2975
rect 15669 2941 15703 2975
rect 15761 2941 15795 2975
rect 17509 2941 17543 2975
rect 6745 2805 6779 2839
rect 7389 2805 7423 2839
rect 8861 2805 8895 2839
rect 16865 2601 16899 2635
rect 17325 2465 17359 2499
rect 17509 2465 17543 2499
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4721 2397 4755 2431
rect 7021 2397 7055 2431
rect 7573 2397 7607 2431
rect 9229 2397 9263 2431
rect 11713 2397 11747 2431
rect 13093 2397 13127 2431
rect 14749 2397 14783 2431
rect 16313 2397 16347 2431
rect 1777 2329 1811 2363
rect 2789 2329 2823 2363
rect 4445 2329 4479 2363
rect 6745 2329 6779 2363
rect 7849 2329 7883 2363
rect 9505 2329 9539 2363
rect 11989 2329 12023 2363
rect 12817 2329 12851 2363
rect 14473 2329 14507 2363
rect 16037 2329 16071 2363
rect 17233 2329 17267 2363
<< metal1 >>
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 14918 17212 14924 17264
rect 14976 17252 14982 17264
rect 15105 17255 15163 17261
rect 15105 17252 15117 17255
rect 14976 17224 15117 17252
rect 14976 17212 14982 17224
rect 15105 17221 15117 17224
rect 15151 17221 15163 17255
rect 15105 17215 15163 17221
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10560 17156 10609 17184
rect 10560 17144 10566 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 15286 17008 15292 17060
rect 15344 17008 15350 17060
rect 10686 16940 10692 16992
rect 10744 16940 10750 16992
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 10468 16612 11437 16640
rect 10468 16600 10474 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14148 16612 14596 16640
rect 14148 16600 14154 16612
rect 11698 16532 11704 16584
rect 11756 16532 11762 16584
rect 14568 16581 14596 16612
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16574 14611 16575
rect 14599 16546 14633 16574
rect 14599 16541 14611 16546
rect 14553 16535 14611 16541
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 16114 16572 16120 16584
rect 15887 16544 16120 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9677 16507 9735 16513
rect 9677 16504 9689 16507
rect 9088 16476 9689 16504
rect 9088 16464 9094 16476
rect 9677 16473 9689 16476
rect 9723 16473 9735 16507
rect 9677 16467 9735 16473
rect 10686 16464 10692 16516
rect 10744 16464 10750 16516
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 14642 16436 14648 16448
rect 14507 16408 14648 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 15102 16396 15108 16448
rect 15160 16396 15166 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15528 16408 15761 16436
rect 15528 16396 15534 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 15749 16399 15807 16405
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 9125 16235 9183 16241
rect 9125 16201 9137 16235
rect 9171 16232 9183 16235
rect 10410 16232 10416 16244
rect 9171 16204 10416 16232
rect 9171 16201 9183 16204
rect 9125 16195 9183 16201
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 11057 16235 11115 16241
rect 11057 16201 11069 16235
rect 11103 16232 11115 16235
rect 11698 16232 11704 16244
rect 11103 16204 11704 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 15010 16232 15016 16244
rect 13464 16204 15016 16232
rect 13464 16173 13492 16204
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 13449 16167 13507 16173
rect 13449 16133 13461 16167
rect 13495 16133 13507 16167
rect 13449 16127 13507 16133
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 9030 16096 9036 16108
rect 8619 16068 9036 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10502 16096 10508 16108
rect 9907 16068 10508 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10502 16056 10508 16068
rect 10560 16096 10566 16108
rect 11054 16096 11060 16108
rect 10560 16068 11060 16096
rect 10560 16056 10566 16068
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11698 16096 11704 16108
rect 11195 16068 11704 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11698 16056 11704 16068
rect 11756 16096 11762 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11756 16068 12173 16096
rect 11756 16056 11762 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13464 16096 13492 16127
rect 14642 16124 14648 16176
rect 14700 16124 14706 16176
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 15197 16167 15255 16173
rect 15197 16164 15209 16167
rect 15160 16136 15209 16164
rect 15160 16124 15166 16136
rect 15197 16133 15209 16136
rect 15243 16133 15255 16167
rect 15197 16127 15255 16133
rect 13035 16068 13492 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 15470 16056 15476 16108
rect 15528 16056 15534 16108
rect 16114 16056 16120 16108
rect 16172 16056 16178 16108
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 10778 15960 10784 15972
rect 5040 15932 10784 15960
rect 5040 15920 5046 15932
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10226 15892 10232 15904
rect 9815 15864 10232 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12802 15892 12808 15904
rect 12299 15864 12808 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13722 15892 13728 15904
rect 12943 15864 13728 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 14608 15864 16037 15892
rect 14608 15852 14614 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 8404 15592 9260 15620
rect 8404 15493 8432 15592
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8536 15524 9137 15552
rect 8536 15512 8542 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9232 15552 9260 15592
rect 11149 15555 11207 15561
rect 11149 15552 11161 15555
rect 9232 15524 11161 15552
rect 9125 15515 9183 15521
rect 11149 15521 11161 15524
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11698 15512 11704 15564
rect 11756 15512 11762 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 12860 15524 13461 15552
rect 12860 15512 12866 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 13722 15512 13728 15564
rect 13780 15512 13786 15564
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 16172 15524 16313 15552
rect 16172 15512 16178 15524
rect 16301 15521 16313 15524
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8389 15487 8447 15493
rect 8389 15484 8401 15487
rect 7975 15456 8401 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8389 15453 8401 15456
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 14240 15456 14289 15484
rect 14240 15444 14246 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 15654 15444 15660 15496
rect 15712 15444 15718 15496
rect 7837 15419 7895 15425
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 9401 15419 9459 15425
rect 9401 15416 9413 15419
rect 7883 15388 9413 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 9401 15385 9413 15388
rect 9447 15385 9459 15419
rect 9401 15379 9459 15385
rect 10410 15376 10416 15428
rect 10468 15376 10474 15428
rect 12710 15376 12716 15428
rect 12768 15376 12774 15428
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 12710 15104 12716 15156
rect 12768 15104 12774 15156
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14182 15144 14188 15156
rect 14139 15116 14188 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 15654 15104 15660 15156
rect 15712 15104 15718 15156
rect 10226 15076 10232 15088
rect 10074 15048 10232 15076
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 15102 15076 15108 15088
rect 14108 15048 15108 15076
rect 14108 15020 14136 15048
rect 15102 15036 15108 15048
rect 15160 15076 15166 15088
rect 15160 15048 15608 15076
rect 15160 15036 15166 15048
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8536 14980 8585 15008
rect 8536 14968 8542 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11882 15008 11888 15020
rect 11112 14980 11888 15008
rect 11112 14968 11118 14980
rect 11882 14968 11888 14980
rect 11940 15008 11946 15020
rect 12805 15011 12863 15017
rect 12805 15008 12817 15011
rect 11940 14980 12817 15008
rect 11940 14968 11946 14980
rect 12805 14977 12817 14980
rect 12851 15008 12863 15011
rect 14090 15008 14096 15020
rect 12851 14980 14096 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15378 15008 15384 15020
rect 14967 14980 15384 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15580 15017 15608 15048
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9398 14940 9404 14952
rect 8895 14912 9404 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 10597 14943 10655 14949
rect 10597 14940 10609 14943
rect 9916 14912 10609 14940
rect 9916 14900 9922 14912
rect 10597 14909 10609 14912
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14884 14912 15117 14940
rect 14884 14900 14890 14912
rect 15105 14909 15117 14912
rect 15151 14940 15163 14943
rect 15286 14940 15292 14952
rect 15151 14912 15292 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 14737 14875 14795 14881
rect 14737 14872 14749 14875
rect 13872 14844 14749 14872
rect 13872 14832 13878 14844
rect 14737 14841 14749 14844
rect 14783 14841 14795 14875
rect 14737 14835 14795 14841
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14240 14368 14473 14396
rect 14240 14356 14246 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14476 14328 14504 14359
rect 15102 14356 15108 14408
rect 15160 14356 15166 14408
rect 15654 14328 15660 14340
rect 14476 14300 15660 14328
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 10226 14260 10232 14272
rect 9999 14232 10232 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 13964 14232 14381 14260
rect 13964 14220 13970 14232
rect 14369 14229 14381 14232
rect 14415 14229 14427 14263
rect 14369 14223 14427 14229
rect 15010 14220 15016 14272
rect 15068 14220 15074 14272
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 9398 14016 9404 14068
rect 9456 14016 9462 14068
rect 13906 13948 13912 14000
rect 13964 13948 13970 14000
rect 15654 13948 15660 14000
rect 15712 13948 15718 14000
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9674 13920 9680 13932
rect 9539 13892 9680 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11146 13920 11152 13932
rect 11011 13892 11152 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10376 13688 10885 13716
rect 10376 13676 10382 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 13630 13472 13636 13524
rect 13688 13472 13694 13524
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10226 13376 10232 13388
rect 9999 13348 10232 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 14645 13311 14703 13317
rect 14645 13308 14657 13311
rect 13771 13280 14657 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 14645 13277 14657 13280
rect 14691 13308 14703 13311
rect 16298 13308 16304 13320
rect 14691 13280 16304 13308
rect 14691 13277 14703 13280
rect 14645 13271 14703 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 10229 13243 10287 13249
rect 10229 13209 10241 13243
rect 10275 13240 10287 13243
rect 10318 13240 10324 13252
rect 10275 13212 10324 13240
rect 10275 13209 10287 13212
rect 10229 13203 10287 13209
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 11790 13240 11796 13252
rect 11454 13212 11796 13240
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 11977 13243 12035 13249
rect 11977 13209 11989 13243
rect 12023 13209 12035 13243
rect 11977 13203 12035 13209
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 7156 13144 7297 13172
rect 7156 13132 7162 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11992 13172 12020 13203
rect 11204 13144 12020 13172
rect 14553 13175 14611 13181
rect 11204 13132 11210 13144
rect 14553 13141 14565 13175
rect 14599 13172 14611 13175
rect 14642 13172 14648 13184
rect 14599 13144 14648 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 7346 12903 7404 12909
rect 7346 12900 7358 12903
rect 7064 12872 7358 12900
rect 7064 12860 7070 12872
rect 7346 12869 7358 12872
rect 7392 12869 7404 12903
rect 15102 12900 15108 12912
rect 7346 12863 7404 12869
rect 14476 12872 15108 12900
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 14476 12841 14504 12872
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14608 12804 14933 12832
rect 14608 12792 14614 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 15120 12832 15148 12860
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15120 12804 15577 12832
rect 14921 12795 14979 12801
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 8478 12588 8484 12640
rect 8536 12588 8542 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 11146 12628 11152 12640
rect 11103 12600 11152 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14148 12600 14381 12628
rect 14148 12588 14154 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 15010 12588 15016 12640
rect 15068 12588 15074 12640
rect 15654 12588 15660 12640
rect 15712 12588 15718 12640
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 11882 12384 11888 12436
rect 11940 12384 11946 12436
rect 7374 12288 7380 12300
rect 4724 12260 7380 12288
rect 4724 12229 4752 12260
rect 7374 12248 7380 12260
rect 7432 12288 7438 12300
rect 8294 12288 8300 12300
rect 7432 12260 8300 12288
rect 7432 12248 7438 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 14642 12288 14648 12300
rect 14599 12260 14648 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6549 12223 6607 12229
rect 6549 12220 6561 12223
rect 6043 12192 6561 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6549 12189 6561 12192
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9582 12220 9588 12232
rect 9355 12192 9588 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 5920 12152 5948 12183
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12220 13691 12223
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13679 12192 14289 12220
rect 13679 12189 13691 12192
rect 13633 12183 13691 12189
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 6270 12152 6276 12164
rect 5920 12124 6276 12152
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 6914 12152 6920 12164
rect 6871 12124 6920 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 7282 12112 7288 12164
rect 7340 12112 7346 12164
rect 8573 12155 8631 12161
rect 8573 12121 8585 12155
rect 8619 12121 8631 12155
rect 8573 12115 8631 12121
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4580 12056 4629 12084
rect 4580 12044 4586 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4617 12047 4675 12053
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8588 12084 8616 12115
rect 10410 12112 10416 12164
rect 10468 12112 10474 12164
rect 13556 12152 13584 12183
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 13906 12152 13912 12164
rect 13556 12124 13912 12152
rect 13906 12112 13912 12124
rect 13964 12152 13970 12164
rect 14550 12152 14556 12164
rect 13964 12124 14556 12152
rect 13964 12112 13970 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 7156 12056 8616 12084
rect 7156 12044 7162 12056
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8720 12056 9229 12084
rect 8720 12044 8726 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 7006 11880 7012 11892
rect 6043 11852 7012 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 9122 11880 9128 11892
rect 7116 11852 9128 11880
rect 5629 11815 5687 11821
rect 5629 11781 5641 11815
rect 5675 11781 5687 11815
rect 5629 11775 5687 11781
rect 5845 11815 5903 11821
rect 5845 11781 5857 11815
rect 5891 11812 5903 11815
rect 7116 11812 7144 11852
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9861 11883 9919 11889
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 10410 11880 10416 11892
rect 9907 11852 10416 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 5891 11784 7144 11812
rect 5891 11781 5903 11784
rect 5845 11775 5903 11781
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4258 11747 4316 11753
rect 4258 11744 4270 11747
rect 3936 11716 4270 11744
rect 3936 11704 3942 11716
rect 4258 11713 4270 11716
rect 4304 11713 4316 11747
rect 4258 11707 4316 11713
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 5644 11744 5672 11775
rect 7926 11772 7932 11824
rect 7984 11772 7990 11824
rect 11149 11815 11207 11821
rect 11149 11781 11161 11815
rect 11195 11812 11207 11815
rect 13814 11812 13820 11824
rect 11195 11784 13820 11812
rect 11195 11781 11207 11784
rect 11149 11775 11207 11781
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 14090 11772 14096 11824
rect 14148 11772 14154 11824
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 15105 11815 15163 11821
rect 15105 11812 15117 11815
rect 15068 11784 15117 11812
rect 15068 11772 15074 11784
rect 15105 11781 15117 11784
rect 15151 11781 15163 11815
rect 15105 11775 15163 11781
rect 6270 11744 6276 11756
rect 5644 11716 6276 11744
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 6420 11648 8401 11676
rect 6420 11636 6426 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13906 11676 13912 11688
rect 13403 11648 13912 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 15378 11636 15384 11688
rect 15436 11636 15442 11688
rect 7098 11608 7104 11620
rect 6840 11580 7104 11608
rect 3145 11543 3203 11549
rect 3145 11509 3157 11543
rect 3191 11540 3203 11543
rect 4338 11540 4344 11552
rect 3191 11512 4344 11540
rect 3191 11509 3203 11512
rect 3145 11503 3203 11509
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 6840 11540 6868 11580
rect 7098 11568 7104 11580
rect 7156 11568 7162 11620
rect 5859 11512 6868 11540
rect 6917 11543 6975 11549
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 6917 11509 6929 11543
rect 6963 11540 6975 11543
rect 7190 11540 7196 11552
rect 6963 11512 7196 11540
rect 6963 11509 6975 11512
rect 6917 11503 6975 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 6362 11296 6368 11348
rect 6420 11296 6426 11348
rect 4338 11268 4344 11280
rect 3252 11240 4344 11268
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3252 11132 3280 11240
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 7190 11268 7196 11280
rect 6328 11240 7196 11268
rect 6328 11228 6334 11240
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8021 11271 8079 11277
rect 8021 11268 8033 11271
rect 7984 11240 8033 11268
rect 7984 11228 7990 11240
rect 8021 11237 8033 11240
rect 8067 11237 8079 11271
rect 8021 11231 8079 11237
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9180 11240 10057 11268
rect 9180 11228 9186 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 4154 11200 4160 11212
rect 3344 11172 4160 11200
rect 3344 11141 3372 11172
rect 4154 11160 4160 11172
rect 4212 11200 4218 11212
rect 4212 11172 7236 11200
rect 4212 11160 4218 11172
rect 3191 11104 3280 11132
rect 3329 11135 3387 11141
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 3421 11067 3479 11073
rect 3421 11033 3433 11067
rect 3467 11064 3479 11067
rect 3467 11036 4370 11064
rect 3467 11033 3479 11036
rect 3421 11027 3479 11033
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 5316 11036 5549 11064
rect 5316 11024 5322 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 5828 11064 5856 11095
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 7208 11141 7236 11172
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 8478 11200 8484 11212
rect 7852 11172 8484 11200
rect 7852 11141 7880 11172
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7193 11135 7251 11141
rect 7055 11104 7144 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7116 11064 7144 11104
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 5828 11036 7144 11064
rect 7208 11064 7236 11095
rect 7944 11064 7972 11095
rect 7208 11036 7972 11064
rect 5537 11027 5595 11033
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3568 10968 4077 10996
rect 3568 10956 3574 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 7116 10996 7144 11036
rect 8036 10996 8064 11172
rect 8478 11160 8484 11172
rect 8536 11200 8542 11212
rect 10873 11203 10931 11209
rect 8536 11172 9168 11200
rect 8536 11160 8542 11172
rect 9140 11141 9168 11172
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 11146 11200 11152 11212
rect 10919 11172 11152 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9416 11064 9444 11095
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9640 11104 9965 11132
rect 9640 11092 9646 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 9416 11036 11100 11064
rect 7116 10968 8064 10996
rect 4065 10959 4123 10965
rect 9214 10956 9220 11008
rect 9272 10956 9278 11008
rect 11072 10996 11100 11036
rect 11146 11024 11152 11076
rect 11204 11024 11210 11076
rect 11882 11024 11888 11076
rect 11940 11024 11946 11076
rect 11974 10996 11980 11008
rect 11072 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 6972 10764 7021 10792
rect 6972 10752 6978 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 7009 10755 7067 10761
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 8386 10792 8392 10804
rect 7699 10764 8392 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 8386 10752 8392 10764
rect 8444 10792 8450 10804
rect 9582 10792 9588 10804
rect 8444 10764 9588 10792
rect 8444 10752 8450 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 11882 10752 11888 10804
rect 11940 10752 11946 10804
rect 3326 10724 3332 10736
rect 2332 10696 3332 10724
rect 2332 10665 2360 10696
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 9214 10724 9220 10736
rect 8694 10696 9220 10724
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 12618 10724 12624 10736
rect 10980 10696 12624 10724
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4120 10628 4186 10656
rect 4120 10616 4126 10628
rect 7098 10616 7104 10668
rect 7156 10616 7162 10668
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10980 10665 11008 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10560 10628 10977 10656
rect 10560 10616 10566 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2777 10591 2835 10597
rect 2777 10588 2789 10591
rect 2271 10560 2789 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2777 10557 2789 10560
rect 2823 10557 2835 10591
rect 2777 10551 2835 10557
rect 3050 10548 3056 10600
rect 3108 10548 3114 10600
rect 9122 10548 9128 10600
rect 9180 10548 9186 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 11808 10588 11836 10619
rect 11974 10616 11980 10668
rect 12032 10616 12038 10668
rect 13170 10588 13176 10600
rect 9447 10560 13176 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 4488 10424 4537 10452
rect 4488 10412 4494 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 4525 10415 4583 10421
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11146 10452 11152 10464
rect 11103 10424 11152 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3050 10248 3056 10260
rect 2731 10220 3056 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 4246 10248 4252 10260
rect 3375 10220 4252 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 4246 10208 4252 10220
rect 4304 10248 4310 10260
rect 5258 10248 5264 10260
rect 4304 10220 5264 10248
rect 4304 10208 4310 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 13170 10208 13176 10260
rect 13228 10208 13234 10260
rect 4062 10140 4068 10192
rect 4120 10140 4126 10192
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8352 10084 11192 10112
rect 8352 10072 8358 10084
rect 2774 10004 2780 10056
rect 2832 10004 2838 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3510 10044 3516 10056
rect 3283 10016 3516 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7524 10016 7757 10044
rect 7524 10004 7530 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8386 10044 8392 10056
rect 7975 10016 8392 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 11164 10053 11192 10084
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11287 10016 11805 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12986 10044 12992 10056
rect 12115 10016 12992 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 7340 9948 7573 9976
rect 7340 9936 7346 9948
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 7561 9939 7619 9945
rect 7650 9936 7656 9988
rect 7708 9936 7714 9988
rect 10597 9911 10655 9917
rect 10597 9877 10609 9911
rect 10643 9908 10655 9911
rect 11698 9908 11704 9920
rect 10643 9880 11704 9908
rect 10643 9877 10655 9880
rect 10597 9871 10655 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11103 9608 11989 9636
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 3970 9528 3976 9580
rect 4028 9528 4034 9580
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 5960 9540 7113 9568
rect 5960 9528 5966 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8478 9568 8484 9580
rect 8159 9540 8484 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 14550 9568 14556 9580
rect 13110 9540 14556 9568
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 2590 9460 2596 9512
rect 2648 9460 2654 9512
rect 2866 9460 2872 9512
rect 2924 9460 2930 9512
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8570 9432 8576 9444
rect 8527 9404 8576 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 3108 9336 4353 9364
rect 3108 9324 3114 9336
rect 4341 9333 4353 9336
rect 4387 9364 4399 9367
rect 7374 9364 7380 9376
rect 4387 9336 7380 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 13446 9324 13452 9376
rect 13504 9324 13510 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2648 9132 2697 9160
rect 2648 9120 2654 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 2924 9132 3341 9160
rect 2924 9120 2930 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 2774 8916 2780 8968
rect 2832 8916 2838 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3108 8928 3249 8956
rect 3108 8916 3114 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3344 8956 3372 9123
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 3973 9163 4031 9169
rect 3973 9160 3985 9163
rect 3936 9132 3985 9160
rect 3936 9120 3942 9132
rect 3973 9129 3985 9132
rect 4019 9129 4031 9163
rect 3973 9123 4031 9129
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 12986 9120 12992 9172
rect 13044 9120 13050 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13228 9132 13676 9160
rect 13228 9120 13234 9132
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 10704 9064 13553 9092
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 3568 8996 5856 9024
rect 3568 8984 3574 8996
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3344 8928 4169 8956
rect 3237 8919 3295 8925
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 5828 8965 5856 8996
rect 7466 8984 7472 9036
rect 7524 8984 7530 9036
rect 10704 8968 10732 9064
rect 13541 9061 13553 9064
rect 13587 9061 13599 9095
rect 13541 9055 13599 9061
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 13446 9024 13452 9036
rect 11020 8996 13452 9024
rect 11020 8984 11026 8996
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6043 8928 7328 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 2792 8888 2820 8916
rect 2792 8860 4384 8888
rect 4356 8829 4384 8860
rect 4522 8848 4528 8900
rect 4580 8848 4586 8900
rect 6914 8848 6920 8900
rect 6972 8848 6978 8900
rect 7009 8891 7067 8897
rect 7009 8857 7021 8891
rect 7055 8888 7067 8891
rect 7300 8888 7328 8928
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9732 8928 9873 8956
rect 9732 8916 9738 8928
rect 9861 8925 9873 8928
rect 9907 8956 9919 8959
rect 10686 8956 10692 8968
rect 9907 8928 10692 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 11790 8956 11796 8968
rect 11072 8928 11796 8956
rect 7466 8888 7472 8900
rect 7055 8860 7236 8888
rect 7300 8860 7472 8888
rect 7055 8857 7067 8860
rect 7009 8851 7067 8857
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 4430 8820 4436 8832
rect 4387 8792 4436 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4430 8780 4436 8792
rect 4488 8820 4494 8832
rect 5166 8820 5172 8832
rect 4488 8792 5172 8820
rect 4488 8780 4494 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 6641 8823 6699 8829
rect 6641 8789 6653 8823
rect 6687 8820 6699 8823
rect 7098 8820 7104 8832
rect 6687 8792 7104 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7208 8820 7236 8860
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 9582 8888 9588 8900
rect 7791 8860 9588 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 9582 8848 9588 8860
rect 9640 8888 9646 8900
rect 11072 8888 11100 8928
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13262 8956 13268 8968
rect 13219 8928 13268 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13372 8965 13400 8996
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13648 8956 13676 9132
rect 14550 9052 14556 9104
rect 14608 9052 14614 9104
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13648 8928 14289 8956
rect 13357 8919 13415 8925
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 9640 8860 11100 8888
rect 9640 8848 9646 8860
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 11204 8860 13308 8888
rect 11204 8848 11210 8860
rect 7282 8820 7288 8832
rect 7208 8792 7288 8820
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7616 8792 7941 8820
rect 7616 8780 7622 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9456 8792 9781 8820
rect 9456 8780 9462 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 13280 8829 13308 8860
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 14476 8888 14504 8919
rect 14056 8860 14504 8888
rect 14056 8848 14062 8860
rect 12069 8823 12127 8829
rect 12069 8820 12081 8823
rect 11112 8792 12081 8820
rect 11112 8780 11118 8792
rect 12069 8789 12081 8792
rect 12115 8789 12127 8823
rect 12069 8783 12127 8789
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5092 8548 5120 8579
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 5224 8588 6745 8616
rect 5224 8576 5230 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7837 8619 7895 8625
rect 7340 8588 7788 8616
rect 7340 8576 7346 8588
rect 4002 8520 5120 8548
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 7469 8551 7527 8557
rect 7469 8548 7481 8551
rect 7248 8520 7481 8548
rect 7248 8508 7254 8520
rect 7469 8517 7481 8520
rect 7515 8517 7527 8551
rect 7469 8511 7527 8517
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4212 8452 4936 8480
rect 4212 8440 4218 8452
rect 2498 8372 2504 8424
rect 2556 8372 2562 8424
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 4908 8412 4936 8452
rect 4982 8440 4988 8492
rect 5040 8440 5046 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5184 8412 5212 8443
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7374 8480 7380 8492
rect 7147 8452 7380 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 5718 8412 5724 8424
rect 4908 8384 5724 8412
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7760 8412 7788 8588
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 10962 8616 10968 8628
rect 7883 8588 10968 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 13446 8576 13452 8628
rect 13504 8576 13510 8628
rect 9398 8508 9404 8560
rect 9456 8508 9462 8560
rect 10410 8508 10416 8560
rect 10468 8508 10474 8560
rect 10686 8508 10692 8560
rect 10744 8548 10750 8560
rect 11149 8551 11207 8557
rect 11149 8548 11161 8551
rect 10744 8520 11161 8548
rect 10744 8508 10750 8520
rect 11149 8517 11161 8520
rect 11195 8517 11207 8551
rect 11149 8511 11207 8517
rect 12710 8508 12716 8560
rect 12768 8508 12774 8560
rect 13464 8548 13492 8576
rect 13464 8520 14044 8548
rect 14016 8489 14044 8520
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 8110 8412 8116 8424
rect 7760 8398 8116 8412
rect 7774 8384 8116 8398
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9490 8412 9496 8424
rect 9171 8384 9496 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 13262 8372 13268 8424
rect 13320 8372 13326 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13587 8384 14105 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 8018 8304 8024 8356
rect 8076 8304 8082 8356
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 2498 8032 2504 8084
rect 2556 8032 2562 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2832 8044 3157 8072
rect 2832 8032 2838 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 7432 8044 9137 8072
rect 7432 8032 7438 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 12710 7964 12716 8016
rect 12768 7964 12774 8016
rect 3970 7896 3976 7948
rect 4028 7896 4034 7948
rect 4522 7936 4528 7948
rect 4080 7908 4528 7936
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 3050 7868 3056 7880
rect 2639 7840 3056 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 4080 7868 4108 7908
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 10502 7936 10508 7948
rect 9723 7908 10508 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 13998 7936 14004 7948
rect 12728 7908 14004 7936
rect 3283 7840 4108 7868
rect 4157 7871 4215 7877
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4172 7800 4200 7831
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4982 7868 4988 7880
rect 4396 7840 4988 7868
rect 4396 7828 4402 7840
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8168 7840 9321 7868
rect 8168 7828 8174 7840
rect 9309 7837 9321 7840
rect 9355 7868 9367 7871
rect 10226 7868 10232 7880
rect 9355 7840 10232 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 11054 7868 11060 7880
rect 10459 7840 11060 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12728 7877 12756 7908
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 15378 7936 15384 7948
rect 14200 7908 15384 7936
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 11940 7840 12725 7868
rect 11940 7828 11946 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13170 7868 13176 7880
rect 13035 7840 13176 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 4172 7772 4936 7800
rect 4908 7744 4936 7772
rect 7006 7760 7012 7812
rect 7064 7760 7070 7812
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 12161 7803 12219 7809
rect 8536 7772 9536 7800
rect 8536 7760 8542 7772
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5721 7735 5779 7741
rect 5721 7732 5733 7735
rect 4948 7704 5733 7732
rect 4948 7692 4954 7704
rect 5721 7701 5733 7704
rect 5767 7732 5779 7735
rect 9306 7732 9312 7744
rect 5767 7704 9312 7732
rect 5767 7701 5779 7704
rect 5721 7695 5779 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 9508 7741 9536 7772
rect 12161 7769 12173 7803
rect 12207 7800 12219 7803
rect 14200 7800 14228 7908
rect 15378 7896 15384 7908
rect 15436 7936 15442 7948
rect 16298 7936 16304 7948
rect 15436 7908 16304 7936
rect 15436 7896 15442 7908
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 12207 7772 14228 7800
rect 14277 7803 14335 7809
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 14277 7769 14289 7803
rect 14323 7769 14335 7803
rect 14277 7763 14335 7769
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14292 7732 14320 7763
rect 15286 7760 15292 7812
rect 15344 7760 15350 7812
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 15988 7772 16037 7800
rect 15988 7760 15994 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 14240 7704 14320 7732
rect 14240 7692 14246 7704
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4580 7500 5089 7528
rect 4580 7488 4586 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 8110 7528 8116 7540
rect 7055 7500 8116 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7024 7460 7052 7491
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7488 8300 7540
rect 8352 7488 8358 7540
rect 10410 7488 10416 7540
rect 10468 7488 10474 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 13262 7528 13268 7540
rect 12023 7500 13268 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 15286 7488 15292 7540
rect 15344 7488 15350 7540
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 4908 7432 7052 7460
rect 9585 7463 9643 7469
rect 4908 7333 4936 7432
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 11054 7460 11060 7472
rect 9631 7432 11060 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 13170 7460 13176 7472
rect 11440 7432 13176 7460
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10413 7395 10471 7401
rect 10413 7392 10425 7395
rect 9364 7364 10425 7392
rect 9364 7352 9370 7364
rect 10413 7361 10425 7364
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 11440 7392 11468 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 13998 7420 14004 7472
rect 14056 7460 14062 7472
rect 14056 7432 15424 7460
rect 14056 7420 14062 7432
rect 10735 7364 11468 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11848 7364 11897 7392
rect 11848 7352 11854 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 15396 7401 15424 7432
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 14240 7364 14289 7392
rect 14240 7352 14246 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 15470 7392 15476 7404
rect 15427 7364 15476 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 14292 7324 14320 7355
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 15856 7324 15884 7355
rect 14292 7296 15884 7324
rect 6638 7216 6644 7268
rect 6696 7216 6702 7268
rect 7193 7259 7251 7265
rect 7193 7225 7205 7259
rect 7239 7256 7251 7259
rect 8386 7256 8392 7268
rect 7239 7228 8392 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 6914 7188 6920 7200
rect 5491 7160 6920 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7374 7188 7380 7200
rect 7055 7160 7380 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 7300 6820 10364 6848
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4798 6780 4804 6792
rect 4203 6752 4804 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4798 6740 4804 6752
rect 4856 6780 4862 6792
rect 6638 6780 6644 6792
rect 4856 6752 6644 6780
rect 4856 6740 4862 6752
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7300 6780 7328 6820
rect 10336 6792 10364 6820
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11940 6820 11989 6848
rect 11940 6808 11946 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 14240 6820 14289 6848
rect 14240 6808 14246 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 7064 6752 7328 6780
rect 7064 6740 7070 6752
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7834 6780 7840 6792
rect 7432 6752 7840 6780
rect 7432 6740 7438 6752
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8210 6783 8268 6789
rect 8210 6780 8222 6783
rect 7984 6752 8222 6780
rect 7984 6740 7990 6752
rect 8210 6749 8222 6752
rect 8256 6749 8268 6783
rect 8210 6743 8268 6749
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10376 6752 10425 6780
rect 10376 6740 10382 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 3384 6684 4721 6712
rect 3384 6672 3390 6684
rect 4709 6681 4721 6684
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 6972 6684 8033 6712
rect 6972 6672 6978 6684
rect 8021 6681 8033 6684
rect 8067 6681 8079 6715
rect 8021 6675 8079 6681
rect 8113 6715 8171 6721
rect 8113 6681 8125 6715
rect 8159 6712 8171 6715
rect 9674 6712 9680 6724
rect 8159 6684 9680 6712
rect 8159 6681 8171 6684
rect 8113 6675 8171 6681
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 14553 6715 14611 6721
rect 14553 6712 14565 6715
rect 14240 6684 14565 6712
rect 14240 6672 14246 6684
rect 14553 6681 14565 6684
rect 14599 6681 14611 6715
rect 14553 6675 14611 6681
rect 15562 6672 15568 6724
rect 15620 6672 15626 6724
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 4028 6616 4077 6644
rect 4028 6604 4034 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 5718 6604 5724 6656
rect 5776 6604 5782 6656
rect 8386 6604 8392 6656
rect 8444 6653 8450 6656
rect 8444 6607 8455 6653
rect 8444 6604 8450 6607
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 16025 6647 16083 6653
rect 16025 6644 16037 6647
rect 14148 6616 16037 6644
rect 14148 6604 14154 6616
rect 16025 6613 16037 6616
rect 16071 6613 16083 6647
rect 16025 6607 16083 6613
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 7561 6443 7619 6449
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 7926 6440 7932 6452
rect 7607 6412 7932 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 14182 6400 14188 6452
rect 14240 6400 14246 6452
rect 15562 6400 15568 6452
rect 15620 6400 15626 6452
rect 3326 6332 3332 6384
rect 3384 6332 3390 6384
rect 3786 6332 3792 6384
rect 3844 6332 3850 6384
rect 8110 6372 8116 6384
rect 7484 6344 8116 6372
rect 7484 6313 7512 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 9214 6332 9220 6384
rect 9272 6332 9278 6384
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7699 6276 7880 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 7852 6248 7880 6276
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 10284 6276 10609 6304
rect 10284 6264 10290 6276
rect 10597 6273 10609 6276
rect 10643 6304 10655 6307
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 10643 6276 11897 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 11885 6273 11897 6276
rect 11931 6304 11943 6307
rect 12618 6304 12624 6316
rect 11931 6276 12624 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 4338 6236 4344 6248
rect 3099 6208 4344 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8202 6236 8208 6248
rect 7892 6208 8208 6236
rect 7892 6196 7898 6208
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 8536 6208 9689 6236
rect 8536 6196 8542 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9999 6208 10517 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11204 6072 11805 6100
rect 11204 6060 11210 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 7098 5896 7104 5908
rect 5776 5868 7104 5896
rect 5776 5856 5782 5868
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 3786 5828 3792 5840
rect 3375 5800 3792 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 3970 5720 3976 5772
rect 4028 5720 4034 5772
rect 8570 5760 8576 5772
rect 7944 5732 8576 5760
rect 2590 5652 2596 5704
rect 2648 5652 2654 5704
rect 3050 5652 3056 5704
rect 3108 5652 3114 5704
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 3510 5692 3516 5704
rect 3375 5664 3516 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 7944 5701 7972 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 11146 5720 11152 5772
rect 11204 5720 11210 5772
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 8260 5664 8401 5692
rect 8260 5652 8266 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 14090 5692 14096 5704
rect 13403 5664 14096 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 2547 5596 4261 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 4249 5593 4261 5596
rect 4295 5593 4307 5627
rect 4249 5587 4307 5593
rect 4798 5584 4804 5636
rect 4856 5584 4862 5636
rect 10888 5624 10916 5655
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 16022 5652 16028 5704
rect 16080 5692 16086 5704
rect 16298 5692 16304 5704
rect 16080 5664 16304 5692
rect 16080 5652 16086 5664
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 11054 5624 11060 5636
rect 10888 5596 11060 5624
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 12158 5584 12164 5636
rect 12216 5584 12222 5636
rect 7837 5559 7895 5565
rect 7837 5525 7849 5559
rect 7883 5556 7895 5559
rect 8202 5556 8208 5568
rect 7883 5528 8208 5556
rect 7883 5525 7895 5528
rect 7837 5519 7895 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 13262 5516 13268 5568
rect 13320 5516 13326 5568
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 15933 5559 15991 5565
rect 15933 5556 15945 5559
rect 15804 5528 15945 5556
rect 15804 5516 15810 5528
rect 15933 5525 15945 5528
rect 15979 5525 15991 5559
rect 15933 5519 15991 5525
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 3418 5312 3424 5364
rect 3476 5312 3482 5364
rect 4798 5312 4804 5364
rect 4856 5312 4862 5364
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 12158 5312 12164 5364
rect 12216 5312 12222 5364
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 3513 5287 3571 5293
rect 3513 5284 3525 5287
rect 3016 5256 3525 5284
rect 3016 5244 3022 5256
rect 3513 5253 3525 5256
rect 3559 5253 3571 5287
rect 5718 5284 5724 5296
rect 3513 5247 3571 5253
rect 3896 5256 5724 5284
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2590 5216 2596 5228
rect 2547 5188 2596 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2590 5176 2596 5188
rect 2648 5216 2654 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 2648 5188 3341 5216
rect 2648 5176 2654 5188
rect 3329 5185 3341 5188
rect 3375 5216 3387 5219
rect 3896 5216 3924 5256
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 16022 5284 16028 5296
rect 8076 5256 8984 5284
rect 8076 5244 8082 5256
rect 3375 5188 3924 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4028 5188 4537 5216
rect 4028 5176 4034 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 4890 5216 4896 5228
rect 4847 5188 4896 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 7340 5188 8125 5216
rect 7340 5176 7346 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 4062 5148 4068 5160
rect 3191 5120 4068 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 8128 5148 8156 5179
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8956 5225 8984 5256
rect 13924 5256 16028 5284
rect 13924 5228 13952 5256
rect 16022 5244 16028 5256
rect 16080 5284 16086 5296
rect 16080 5256 16574 5284
rect 16080 5244 16086 5256
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8628 5188 8769 5216
rect 8628 5176 8634 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 11146 5176 11152 5228
rect 11204 5176 11210 5228
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 11940 5188 12265 5216
rect 11940 5176 11946 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12299 5188 12909 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13906 5176 13912 5228
rect 13964 5176 13970 5228
rect 14737 5219 14795 5225
rect 14737 5185 14749 5219
rect 14783 5216 14795 5219
rect 14826 5216 14832 5228
rect 14783 5188 14832 5216
rect 14783 5185 14795 5188
rect 14737 5179 14795 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15654 5216 15660 5228
rect 14967 5188 15660 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16546 5216 16574 5256
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16546 5188 16957 5216
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17862 5176 17868 5228
rect 17920 5176 17926 5228
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8128 5120 8861 5148
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 14844 5148 14872 5176
rect 15838 5148 15844 5160
rect 14844 5120 15844 5148
rect 8849 5111 8907 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5148 18199 5151
rect 19058 5148 19064 5160
rect 18187 5120 19064 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 7926 5040 7932 5092
rect 7984 5040 7990 5092
rect 16206 5040 16212 5092
rect 16264 5040 16270 5092
rect 16301 5083 16359 5089
rect 16301 5049 16313 5083
rect 16347 5080 16359 5083
rect 16942 5080 16948 5092
rect 16347 5052 16948 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 5166 5012 5172 5024
rect 3743 4984 5172 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 12802 4972 12808 5024
rect 12860 4972 12866 5024
rect 13998 4972 14004 5024
rect 14056 4972 14062 5024
rect 14553 5015 14611 5021
rect 14553 4981 14565 5015
rect 14599 5012 14611 5015
rect 14642 5012 14648 5024
rect 14599 4984 14648 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16908 4984 17049 5012
rect 16908 4972 16914 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17037 4975 17095 4981
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4808 2559 4811
rect 2958 4808 2964 4820
rect 2547 4780 2964 4808
rect 2547 4777 2559 4780
rect 2501 4771 2559 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 9674 4808 9680 4820
rect 7524 4780 9680 4808
rect 7524 4768 7530 4780
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 11425 4811 11483 4817
rect 11425 4808 11437 4811
rect 11204 4780 11437 4808
rect 11204 4768 11210 4780
rect 11425 4777 11437 4780
rect 11471 4777 11483 4811
rect 11425 4771 11483 4777
rect 4430 4740 4436 4752
rect 2746 4712 4436 4740
rect 2746 4672 2774 4712
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 9122 4700 9128 4752
rect 9180 4700 9186 4752
rect 15197 4743 15255 4749
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 15286 4740 15292 4752
rect 15243 4712 15292 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 15286 4700 15292 4712
rect 15344 4700 15350 4752
rect 17129 4743 17187 4749
rect 17129 4709 17141 4743
rect 17175 4709 17187 4743
rect 17129 4703 17187 4709
rect 4890 4672 4896 4684
rect 2424 4644 2774 4672
rect 4172 4644 4896 4672
rect 2424 4613 2452 4644
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 1995 4576 2421 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 3050 4564 3056 4616
rect 3108 4564 3114 4616
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 3510 4604 3516 4616
rect 3375 4576 3516 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3510 4564 3516 4576
rect 3568 4604 3574 4616
rect 4172 4613 4200 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 13173 4675 13231 4681
rect 7331 4644 8064 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3568 4576 4169 4604
rect 3568 4564 3574 4576
rect 4157 4573 4169 4576
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7466 4604 7472 4616
rect 7423 4576 7472 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 3068 4536 3096 4564
rect 3970 4536 3976 4548
rect 3068 4508 3976 4536
rect 3970 4496 3976 4508
rect 4028 4536 4034 4548
rect 4264 4536 4292 4567
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8036 4613 8064 4644
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13262 4672 13268 4684
rect 13219 4644 13268 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14826 4632 14832 4684
rect 14884 4632 14890 4684
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8110 4604 8116 4616
rect 8067 4576 8116 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8570 4604 8576 4616
rect 8343 4576 8576 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8570 4564 8576 4576
rect 8628 4604 8634 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8628 4576 9413 4604
rect 8628 4564 8634 4576
rect 9401 4573 9413 4576
rect 9447 4604 9459 4607
rect 9582 4604 9588 4616
rect 9447 4576 9588 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 17144 4604 17172 4703
rect 17218 4604 17224 4616
rect 17144 4576 17224 4604
rect 17218 4564 17224 4576
rect 17276 4604 17282 4616
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17276 4576 17601 4604
rect 17276 4564 17282 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 4028 4508 4292 4536
rect 8128 4536 8156 4564
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8128 4508 9137 4536
rect 4028 4496 4034 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 12802 4536 12808 4548
rect 12466 4508 12808 4536
rect 9125 4499 9183 4505
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 12894 4496 12900 4548
rect 12952 4496 12958 4548
rect 16016 4539 16074 4545
rect 16016 4505 16028 4539
rect 16062 4536 16074 4539
rect 16298 4536 16304 4548
rect 16062 4508 16304 4536
rect 16062 4505 16074 4508
rect 16016 4499 16074 4505
rect 16298 4496 16304 4508
rect 16356 4496 16362 4548
rect 17402 4496 17408 4548
rect 17460 4536 17466 4548
rect 17865 4539 17923 4545
rect 17865 4536 17877 4539
rect 17460 4508 17877 4536
rect 17460 4496 17466 4508
rect 17865 4505 17877 4508
rect 17911 4505 17923 4539
rect 17865 4499 17923 4505
rect 1854 4428 1860 4480
rect 1912 4428 1918 4480
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4062 4428 4068 4480
rect 4120 4428 4126 4480
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 7837 4471 7895 4477
rect 7837 4468 7849 4471
rect 7432 4440 7849 4468
rect 7432 4428 7438 4440
rect 7837 4437 7849 4440
rect 7883 4437 7895 4471
rect 7837 4431 7895 4437
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 8076 4440 8217 4468
rect 8076 4428 8082 4440
rect 8205 4437 8217 4440
rect 8251 4468 8263 4471
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 8251 4440 9321 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 9309 4431 9367 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15289 4471 15347 4477
rect 15289 4468 15301 4471
rect 15252 4440 15301 4468
rect 15252 4428 15258 4440
rect 15289 4437 15301 4440
rect 15335 4437 15347 4471
rect 15289 4431 15347 4437
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 7190 4264 7196 4276
rect 4488 4236 7196 4264
rect 4488 4224 4494 4236
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8757 4267 8815 4273
rect 8757 4264 8769 4267
rect 8076 4236 8769 4264
rect 8076 4224 8082 4236
rect 8757 4233 8769 4236
rect 8803 4264 8815 4267
rect 8803 4236 9536 4264
rect 8803 4233 8815 4236
rect 8757 4227 8815 4233
rect 3326 4156 3332 4208
rect 3384 4156 3390 4208
rect 9508 4205 9536 4236
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12952 4236 13461 4264
rect 12952 4224 12958 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 16298 4224 16304 4276
rect 16356 4224 16362 4276
rect 9493 4199 9551 4205
rect 6840 4168 7972 4196
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1912 4100 2421 4128
rect 1912 4088 1918 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4212 4100 4445 4128
rect 4212 4088 4218 4100
rect 4433 4097 4445 4100
rect 4479 4128 4491 4131
rect 4982 4128 4988 4140
rect 4479 4100 4988 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6840 4137 6868 4168
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6788 4100 6837 4128
rect 6788 4088 6794 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 6972 4100 7573 4128
rect 6972 4088 6978 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7944 4128 7972 4168
rect 9493 4165 9505 4199
rect 9539 4165 9551 4199
rect 9493 4159 9551 4165
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 12912 4196 12940 4224
rect 15010 4196 15016 4208
rect 9640 4168 10180 4196
rect 9640 4156 9646 4168
rect 8386 4128 8392 4140
rect 7944 4100 8392 4128
rect 7837 4091 7895 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3050 4060 3056 4072
rect 2731 4032 3056 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 7852 4060 7880 4091
rect 8386 4088 8392 4100
rect 8444 4128 8450 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8444 4100 8585 4128
rect 8444 4088 8450 4100
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 6840 4032 7880 4060
rect 6840 3936 6868 4032
rect 8110 4020 8116 4072
rect 8168 4060 8174 4072
rect 8864 4060 8892 4091
rect 9674 4088 9680 4140
rect 9732 4088 9738 4140
rect 10152 4137 10180 4168
rect 12636 4168 12940 4196
rect 13004 4168 15016 4196
rect 12636 4137 12664 4168
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 8168 4032 8892 4060
rect 9692 4060 9720 4088
rect 10336 4060 10364 4091
rect 12710 4088 12716 4140
rect 12768 4088 12774 4140
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13004 4128 13032 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 15838 4156 15844 4208
rect 15896 4156 15902 4208
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 17098 4199 17156 4205
rect 17098 4196 17110 4199
rect 17000 4168 17110 4196
rect 17000 4156 17006 4168
rect 17098 4165 17110 4168
rect 17144 4165 17156 4199
rect 17098 4159 17156 4165
rect 12943 4100 13032 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13354 4088 13360 4140
rect 13412 4088 13418 4140
rect 13998 4088 14004 4140
rect 14056 4088 14062 4140
rect 14268 4131 14326 4137
rect 14268 4097 14280 4131
rect 14314 4128 14326 4131
rect 14642 4128 14648 4140
rect 14314 4100 14648 4128
rect 14314 4097 14326 4100
rect 14268 4091 14326 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 16850 4088 16856 4140
rect 16908 4088 16914 4140
rect 9692 4032 10364 4060
rect 8168 4020 8174 4032
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 7653 3995 7711 4001
rect 7653 3992 7665 3995
rect 7156 3964 7665 3992
rect 7156 3952 7162 3964
rect 7653 3961 7665 3964
rect 7699 3992 7711 3995
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 7699 3964 10149 3992
rect 7699 3961 7711 3964
rect 7653 3955 7711 3961
rect 10137 3961 10149 3964
rect 10183 3961 10195 3995
rect 10137 3955 10195 3961
rect 16209 3995 16267 4001
rect 16209 3961 16221 3995
rect 16255 3992 16267 3995
rect 16850 3992 16856 4004
rect 16255 3964 16856 3992
rect 16255 3961 16267 3964
rect 16209 3955 16267 3961
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 6822 3884 6828 3936
rect 6880 3884 6886 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 7064 3896 7389 3924
rect 7064 3884 7070 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 8386 3924 8392 3936
rect 7800 3896 8392 3924
rect 7800 3884 7806 3896
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 8628 3896 9413 3924
rect 8628 3884 8634 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 15381 3927 15439 3933
rect 15381 3893 15393 3927
rect 15427 3924 15439 3927
rect 15562 3924 15568 3936
rect 15427 3896 15568 3924
rect 15427 3893 15439 3896
rect 15381 3887 15439 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17920 3896 18245 3924
rect 17920 3884 17926 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 3050 3680 3056 3732
rect 3108 3680 3114 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 4028 3692 4077 3720
rect 4028 3680 4034 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 6914 3720 6920 3732
rect 6411 3692 6920 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7374 3720 7380 3732
rect 7239 3692 7380 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7208 3584 7236 3683
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 8444 3692 9229 3720
rect 8444 3680 8450 3692
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 9217 3683 9275 3689
rect 12710 3680 12716 3732
rect 12768 3680 12774 3732
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 15712 3692 16773 3720
rect 15712 3680 15718 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 16761 3683 16819 3689
rect 6380 3556 7236 3584
rect 7285 3587 7343 3593
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 4154 3516 4160 3528
rect 3191 3488 4160 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 5166 3476 5172 3528
rect 5224 3525 5230 3528
rect 5224 3516 5236 3525
rect 5445 3519 5503 3525
rect 5224 3488 5269 3516
rect 5224 3479 5236 3488
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5718 3516 5724 3528
rect 5491 3488 5724 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5224 3476 5230 3479
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6380 3525 6408 3556
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7926 3584 7932 3596
rect 7331 3556 7932 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 17405 3587 17463 3593
rect 8352 3556 10732 3584
rect 8352 3544 8358 3556
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 6196 3448 6224 3479
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6880 3488 7021 3516
rect 6880 3476 6886 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7024 3448 7052 3479
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8202 3476 8208 3528
rect 8260 3476 8266 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8404 3448 8432 3479
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 10704 3525 10732 3556
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 17494 3584 17500 3596
rect 17451 3556 17500 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 10827 3488 11345 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 13354 3516 13360 3528
rect 11333 3479 11391 3485
rect 12406 3488 13360 3516
rect 8662 3448 8668 3460
rect 6196 3420 6960 3448
rect 7024 3420 8668 3448
rect 6822 3340 6828 3392
rect 6880 3340 6886 3392
rect 6932 3380 6960 3420
rect 8662 3408 8668 3420
rect 8720 3448 8726 3460
rect 9416 3448 9444 3479
rect 8720 3420 9444 3448
rect 8720 3408 8726 3420
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11578 3451 11636 3457
rect 11578 3448 11590 3451
rect 11204 3420 11590 3448
rect 11204 3408 11210 3420
rect 11578 3417 11590 3420
rect 11624 3448 11636 3451
rect 12406 3448 12434 3488
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 15194 3525 15200 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13964 3488 14289 3516
rect 13964 3476 13970 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14415 3488 14933 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 15188 3516 15200 3525
rect 15155 3488 15200 3516
rect 14921 3479 14979 3485
rect 15188 3479 15200 3488
rect 15194 3476 15200 3479
rect 15252 3476 15258 3528
rect 11624 3420 12434 3448
rect 11624 3417 11636 3420
rect 11578 3411 11636 3417
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 17129 3451 17187 3457
rect 17129 3448 17141 3451
rect 15620 3420 17141 3448
rect 15620 3408 15626 3420
rect 17129 3417 17141 3420
rect 17175 3417 17187 3451
rect 17129 3411 17187 3417
rect 7282 3380 7288 3392
rect 6932 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7524 3352 7757 3380
rect 7524 3340 7530 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7745 3343 7803 3349
rect 9585 3383 9643 3389
rect 9585 3349 9597 3383
rect 9631 3380 9643 3383
rect 11698 3380 11704 3392
rect 9631 3352 11704 3380
rect 9631 3349 9643 3352
rect 9585 3343 9643 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 16298 3340 16304 3392
rect 16356 3340 16362 3392
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 17310 3380 17316 3392
rect 17267 3352 17316 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 17310 3340 17316 3352
rect 17368 3380 17374 3392
rect 17862 3380 17868 3392
rect 17368 3352 17868 3380
rect 17368 3340 17374 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 4430 3136 4436 3188
rect 4488 3136 4494 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5718 3176 5724 3188
rect 5583 3148 5724 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15286 3176 15292 3188
rect 15243 3148 15292 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 16850 3136 16856 3188
rect 16908 3136 16914 3188
rect 17218 3136 17224 3188
rect 17276 3136 17282 3188
rect 2958 3068 2964 3120
rect 3016 3068 3022 3120
rect 8294 3108 8300 3120
rect 5644 3080 8300 3108
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2648 3012 2697 3040
rect 2648 3000 2654 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 5644 3049 5672 3080
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 16298 3108 16304 3120
rect 15611 3080 16304 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 16298 3068 16304 3080
rect 16356 3108 16362 3120
rect 17313 3111 17371 3117
rect 17313 3108 17325 3111
rect 16356 3080 17325 3108
rect 16356 3068 16362 3080
rect 17313 3077 17325 3080
rect 17359 3077 17371 3111
rect 17313 3071 17371 3077
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6788 3012 6929 3040
rect 6788 3000 6794 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 8570 3040 8576 3052
rect 7791 3012 8576 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 6638 2932 6644 2984
rect 6696 2932 6702 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 7098 2972 7104 2984
rect 6871 2944 7104 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 6656 2904 6684 2932
rect 7760 2904 7788 3003
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 8662 3000 8668 3052
rect 8720 3000 8726 3052
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15068 3012 15792 3040
rect 15068 3000 15074 3012
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2972 7895 2975
rect 7926 2972 7932 2984
rect 7883 2944 7932 2972
rect 7883 2941 7895 2944
rect 7837 2935 7895 2941
rect 7926 2932 7932 2944
rect 7984 2972 7990 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7984 2944 8401 2972
rect 7984 2932 7990 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 9122 2972 9128 2984
rect 8527 2944 9128 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 15654 2932 15660 2984
rect 15712 2932 15718 2984
rect 15764 2981 15792 3012
rect 15749 2975 15807 2981
rect 15749 2941 15761 2975
rect 15795 2972 15807 2975
rect 17494 2972 17500 2984
rect 15795 2944 17500 2972
rect 15795 2941 15807 2944
rect 15749 2935 15807 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 6656 2876 7788 2904
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 6733 2839 6791 2845
rect 6733 2836 6745 2839
rect 5592 2808 6745 2836
rect 5592 2796 5598 2808
rect 6733 2805 6745 2808
rect 6779 2805 6791 2839
rect 6733 2799 6791 2805
rect 7374 2796 7380 2848
rect 7432 2796 7438 2848
rect 8849 2839 8907 2845
rect 8849 2805 8861 2839
rect 8895 2836 8907 2839
rect 9214 2836 9220 2848
rect 8895 2808 9220 2836
rect 8895 2805 8907 2808
rect 8849 2799 8907 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16264 2604 16865 2632
rect 16264 2592 16270 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 16853 2595 16911 2601
rect 7374 2496 7380 2508
rect 2056 2468 7380 2496
rect 2056 2437 2084 2468
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7524 2468 7604 2496
rect 7524 2456 7530 2468
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 4709 2431 4767 2437
rect 3099 2400 4660 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 842 2320 848 2372
rect 900 2360 906 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 900 2332 1777 2360
rect 900 2320 906 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2556 2332 2789 2360
rect 2556 2320 2562 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4433 2363 4491 2369
rect 4433 2360 4445 2363
rect 4212 2332 4445 2360
rect 4212 2320 4218 2332
rect 4433 2329 4445 2332
rect 4479 2329 4491 2363
rect 4632 2360 4660 2400
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5534 2428 5540 2440
rect 4755 2400 5540 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6822 2428 6828 2440
rect 5644 2400 6828 2428
rect 5644 2360 5672 2400
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 7006 2388 7012 2440
rect 7064 2388 7070 2440
rect 7576 2437 7604 2468
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 17276 2468 17325 2496
rect 17276 2456 17282 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17494 2456 17500 2508
rect 17552 2456 17558 2508
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 9214 2388 9220 2440
rect 9272 2388 9278 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 13354 2428 13360 2440
rect 13127 2400 13360 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2428 14795 2431
rect 15654 2428 15660 2440
rect 14783 2400 15660 2428
rect 14783 2397 14795 2400
rect 14737 2391 14795 2397
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 16298 2388 16304 2440
rect 16356 2388 16362 2440
rect 4632 2332 5672 2360
rect 4433 2323 4491 2329
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 5868 2332 6745 2360
rect 5868 2320 5874 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 6733 2323 6791 2329
rect 7466 2320 7472 2372
rect 7524 2360 7530 2372
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 7524 2332 7849 2360
rect 7524 2320 7530 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 7837 2323 7895 2329
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 9180 2332 9505 2360
rect 9180 2320 9186 2332
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 9493 2323 9551 2329
rect 11054 2320 11060 2372
rect 11112 2360 11118 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11112 2332 11989 2360
rect 11112 2320 11118 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12805 2363 12863 2369
rect 12805 2360 12817 2363
rect 12492 2332 12817 2360
rect 12492 2320 12498 2332
rect 12805 2329 12817 2332
rect 12851 2329 12863 2363
rect 12805 2323 12863 2329
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 14148 2332 14473 2360
rect 14148 2320 14154 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 15746 2320 15752 2372
rect 15804 2360 15810 2372
rect 16025 2363 16083 2369
rect 16025 2360 16037 2363
rect 15804 2332 16037 2360
rect 15804 2320 15810 2332
rect 16025 2329 16037 2332
rect 16071 2329 16083 2363
rect 16025 2323 16083 2329
rect 17221 2363 17279 2369
rect 17221 2329 17233 2363
rect 17267 2360 17279 2363
rect 17310 2360 17316 2372
rect 17267 2332 17316 2360
rect 17267 2329 17279 2332
rect 17221 2323 17279 2329
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 14924 17212 14976 17264
rect 10508 17144 10560 17196
rect 15292 17051 15344 17060
rect 15292 17017 15301 17051
rect 15301 17017 15335 17051
rect 15335 17017 15344 17051
rect 15292 17008 15344 17017
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 10416 16600 10468 16652
rect 14096 16600 14148 16652
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 16120 16532 16172 16584
rect 9036 16464 9088 16516
rect 10692 16464 10744 16516
rect 14648 16396 14700 16448
rect 15108 16439 15160 16448
rect 15108 16405 15117 16439
rect 15117 16405 15151 16439
rect 15151 16405 15160 16439
rect 15108 16396 15160 16405
rect 15476 16396 15528 16448
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 10416 16192 10468 16244
rect 11704 16192 11756 16244
rect 15016 16192 15068 16244
rect 9036 16099 9088 16108
rect 9036 16065 9045 16099
rect 9045 16065 9079 16099
rect 9079 16065 9088 16099
rect 9036 16056 9088 16065
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 11060 16056 11112 16108
rect 11704 16056 11756 16108
rect 14648 16124 14700 16176
rect 15108 16124 15160 16176
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 4988 15920 5040 15972
rect 10784 15920 10836 15972
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 10232 15852 10284 15904
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 12808 15852 12860 15904
rect 13728 15852 13780 15904
rect 14556 15852 14608 15904
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 8484 15512 8536 15564
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 12808 15512 12860 15564
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 16120 15512 16172 15564
rect 14188 15444 14240 15496
rect 15660 15444 15712 15496
rect 10416 15376 10468 15428
rect 12716 15376 12768 15428
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 12716 15147 12768 15156
rect 12716 15113 12725 15147
rect 12725 15113 12759 15147
rect 12759 15113 12768 15147
rect 12716 15104 12768 15113
rect 14188 15104 14240 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 10232 15036 10284 15088
rect 15108 15036 15160 15088
rect 8484 14968 8536 15020
rect 11060 14968 11112 15020
rect 11888 14968 11940 15020
rect 14096 14968 14148 15020
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 15384 14968 15436 15020
rect 9404 14900 9456 14952
rect 9864 14900 9916 14952
rect 14832 14900 14884 14952
rect 15292 14900 15344 14952
rect 13820 14832 13872 14884
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 14188 14356 14240 14408
rect 15108 14399 15160 14408
rect 15108 14365 15117 14399
rect 15117 14365 15151 14399
rect 15151 14365 15160 14399
rect 15108 14356 15160 14365
rect 15660 14288 15712 14340
rect 10232 14220 10284 14272
rect 13912 14220 13964 14272
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 13912 13991 13964 14000
rect 13912 13957 13921 13991
rect 13921 13957 13955 13991
rect 13955 13957 13964 13991
rect 13912 13948 13964 13957
rect 15660 13991 15712 14000
rect 15660 13957 15669 13991
rect 15669 13957 15703 13991
rect 15703 13957 15712 13991
rect 15660 13948 15712 13957
rect 9680 13880 9732 13932
rect 11152 13880 11204 13932
rect 15016 13880 15068 13932
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 10324 13676 10376 13728
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 10232 13336 10284 13388
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 16304 13268 16356 13320
rect 10324 13200 10376 13252
rect 11796 13200 11848 13252
rect 7104 13132 7156 13184
rect 11152 13132 11204 13184
rect 14648 13132 14700 13184
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 7012 12860 7064 12912
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 15108 12860 15160 12912
rect 14556 12792 14608 12844
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 11152 12588 11204 12640
rect 14096 12588 14148 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 7380 12248 7432 12300
rect 8300 12248 8352 12300
rect 14648 12248 14700 12300
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 9588 12180 9640 12232
rect 6276 12112 6328 12164
rect 6920 12112 6972 12164
rect 7288 12112 7340 12164
rect 4528 12044 4580 12096
rect 7104 12044 7156 12096
rect 10416 12155 10468 12164
rect 10416 12121 10425 12155
rect 10425 12121 10459 12155
rect 10459 12121 10468 12155
rect 10416 12112 10468 12121
rect 15660 12180 15712 12232
rect 13912 12112 13964 12164
rect 14556 12112 14608 12164
rect 8668 12044 8720 12096
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 7012 11840 7064 11892
rect 9128 11840 9180 11892
rect 10416 11840 10468 11892
rect 3884 11704 3936 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 7932 11772 7984 11824
rect 13820 11772 13872 11824
rect 14096 11772 14148 11824
rect 15016 11772 15068 11824
rect 6276 11704 6328 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 6368 11636 6420 11688
rect 13912 11636 13964 11688
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 4344 11500 4396 11552
rect 7104 11568 7156 11620
rect 7196 11500 7248 11552
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 4344 11228 4396 11280
rect 6276 11228 6328 11280
rect 7196 11228 7248 11280
rect 7932 11228 7984 11280
rect 9128 11228 9180 11280
rect 4160 11160 4212 11212
rect 5264 11024 5316 11076
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 3516 10956 3568 11008
rect 8484 11160 8536 11212
rect 11152 11160 11204 11212
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 9588 11092 9640 11144
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 11152 11067 11204 11076
rect 11152 11033 11161 11067
rect 11161 11033 11195 11067
rect 11195 11033 11204 11067
rect 11152 11024 11204 11033
rect 11888 11024 11940 11076
rect 11980 10956 12032 11008
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 6920 10752 6972 10804
rect 8392 10752 8444 10804
rect 9588 10752 9640 10804
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 3332 10684 3384 10736
rect 9220 10684 9272 10736
rect 4068 10616 4120 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 10508 10616 10560 10668
rect 12624 10684 12676 10736
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 13176 10548 13228 10600
rect 4436 10412 4488 10464
rect 11152 10412 11204 10464
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 3056 10208 3108 10260
rect 4252 10208 4304 10260
rect 5264 10208 5316 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 4068 10183 4120 10192
rect 4068 10149 4077 10183
rect 4077 10149 4111 10183
rect 4111 10149 4120 10183
rect 4068 10140 4120 10149
rect 8300 10072 8352 10124
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 3516 10004 3568 10056
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 7472 10004 7524 10056
rect 8392 10004 8444 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 12992 10004 13044 10056
rect 7288 9936 7340 9988
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 7656 9936 7708 9945
rect 11704 9868 11756 9920
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 3976 9528 4028 9580
rect 5908 9528 5960 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 8484 9528 8536 9580
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 14556 9528 14608 9580
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 8576 9392 8628 9444
rect 3056 9324 3108 9376
rect 7380 9324 7432 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 2596 9120 2648 9172
rect 2872 9120 2924 9172
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 3056 8916 3108 8968
rect 3884 9120 3936 9172
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 12992 9163 13044 9172
rect 12992 9129 13001 9163
rect 13001 9129 13035 9163
rect 13035 9129 13044 9163
rect 12992 9120 13044 9129
rect 13176 9120 13228 9172
rect 3516 8984 3568 9036
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 7472 8984 7524 9036
rect 10968 8984 11020 9036
rect 4528 8891 4580 8900
rect 4528 8857 4537 8891
rect 4537 8857 4571 8891
rect 4571 8857 4580 8891
rect 4528 8848 4580 8857
rect 6920 8891 6972 8900
rect 6920 8857 6929 8891
rect 6929 8857 6963 8891
rect 6963 8857 6972 8891
rect 6920 8848 6972 8857
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 9680 8916 9732 8968
rect 10692 8916 10744 8968
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 4436 8780 4488 8832
rect 5172 8780 5224 8832
rect 7104 8780 7156 8832
rect 7472 8848 7524 8900
rect 9588 8848 9640 8900
rect 11796 8916 11848 8968
rect 13268 8916 13320 8968
rect 13452 8984 13504 9036
rect 14556 9095 14608 9104
rect 14556 9061 14565 9095
rect 14565 9061 14599 9095
rect 14599 9061 14608 9095
rect 14556 9052 14608 9061
rect 11152 8848 11204 8900
rect 7288 8780 7340 8832
rect 7564 8780 7616 8832
rect 9404 8780 9456 8832
rect 11060 8780 11112 8832
rect 14004 8848 14056 8900
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 5172 8576 5224 8628
rect 7288 8576 7340 8628
rect 7196 8508 7248 8560
rect 4160 8440 4212 8492
rect 2504 8415 2556 8424
rect 2504 8381 2513 8415
rect 2513 8381 2547 8415
rect 2547 8381 2556 8415
rect 2504 8372 2556 8381
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7380 8440 7432 8492
rect 5724 8372 5776 8424
rect 10968 8576 11020 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 13452 8576 13504 8628
rect 9404 8551 9456 8560
rect 9404 8517 9413 8551
rect 9413 8517 9447 8551
rect 9447 8517 9456 8551
rect 9404 8508 9456 8517
rect 10416 8508 10468 8560
rect 10692 8508 10744 8560
rect 12716 8508 12768 8560
rect 8116 8372 8168 8424
rect 9496 8372 9548 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 2504 8032 2556 8041
rect 2780 8032 2832 8084
rect 7380 8032 7432 8084
rect 12716 8007 12768 8016
rect 12716 7973 12725 8007
rect 12725 7973 12759 8007
rect 12759 7973 12768 8007
rect 12716 7964 12768 7973
rect 3976 7939 4028 7948
rect 3976 7905 3985 7939
rect 3985 7905 4019 7939
rect 4019 7905 4028 7939
rect 3976 7896 4028 7905
rect 3056 7828 3108 7880
rect 4528 7896 4580 7948
rect 10508 7896 10560 7948
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4988 7828 5040 7880
rect 8116 7828 8168 7880
rect 10232 7828 10284 7880
rect 11060 7828 11112 7880
rect 11888 7828 11940 7880
rect 14004 7896 14056 7948
rect 13176 7828 13228 7880
rect 7012 7803 7064 7812
rect 7012 7769 7021 7803
rect 7021 7769 7055 7803
rect 7055 7769 7064 7803
rect 7012 7760 7064 7769
rect 8484 7760 8536 7812
rect 4896 7692 4948 7744
rect 9312 7692 9364 7744
rect 15384 7896 15436 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 14188 7692 14240 7744
rect 15292 7760 15344 7812
rect 15936 7760 15988 7812
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 4528 7488 4580 7540
rect 8116 7488 8168 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 10416 7531 10468 7540
rect 10416 7497 10425 7531
rect 10425 7497 10459 7531
rect 10459 7497 10468 7531
rect 10416 7488 10468 7497
rect 13268 7488 13320 7540
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 11060 7420 11112 7472
rect 9312 7352 9364 7404
rect 13176 7420 13228 7472
rect 14004 7420 14056 7472
rect 11796 7352 11848 7404
rect 14188 7352 14240 7404
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 15476 7352 15528 7404
rect 6644 7259 6696 7268
rect 6644 7225 6653 7259
rect 6653 7225 6687 7259
rect 6687 7225 6696 7259
rect 6644 7216 6696 7225
rect 8392 7216 8444 7268
rect 6920 7148 6972 7200
rect 7380 7148 7432 7200
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 6644 6740 6696 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 11888 6808 11940 6860
rect 14188 6808 14240 6860
rect 7012 6740 7064 6749
rect 7380 6740 7432 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 7932 6740 7984 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10324 6740 10376 6792
rect 3332 6672 3384 6724
rect 6920 6672 6972 6724
rect 9680 6672 9732 6724
rect 14188 6672 14240 6724
rect 15568 6672 15620 6724
rect 3976 6604 4028 6656
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 8392 6647 8444 6656
rect 8392 6613 8409 6647
rect 8409 6613 8443 6647
rect 8443 6613 8444 6647
rect 8392 6604 8444 6613
rect 14096 6604 14148 6656
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 7932 6400 7984 6452
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 15568 6443 15620 6452
rect 15568 6409 15577 6443
rect 15577 6409 15611 6443
rect 15611 6409 15620 6443
rect 15568 6400 15620 6409
rect 3332 6375 3384 6384
rect 3332 6341 3341 6375
rect 3341 6341 3375 6375
rect 3375 6341 3384 6375
rect 3332 6332 3384 6341
rect 3792 6332 3844 6384
rect 8116 6332 8168 6384
rect 9220 6332 9272 6384
rect 10232 6264 10284 6316
rect 12624 6264 12676 6316
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 4344 6196 4396 6248
rect 7840 6196 7892 6248
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 8484 6196 8536 6248
rect 11152 6060 11204 6112
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 7104 5856 7156 5908
rect 8484 5899 8536 5908
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 3792 5788 3844 5840
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3516 5652 3568 5704
rect 8576 5720 8628 5772
rect 11152 5763 11204 5772
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11152 5720 11204 5729
rect 8208 5652 8260 5704
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 4804 5584 4856 5636
rect 14096 5652 14148 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16304 5652 16356 5704
rect 11060 5584 11112 5636
rect 12164 5584 12216 5636
rect 8208 5516 8260 5568
rect 13268 5559 13320 5568
rect 13268 5525 13277 5559
rect 13277 5525 13311 5559
rect 13311 5525 13320 5559
rect 13268 5516 13320 5525
rect 15752 5516 15804 5568
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 3424 5355 3476 5364
rect 3424 5321 3433 5355
rect 3433 5321 3467 5355
rect 3467 5321 3476 5355
rect 3424 5312 3476 5321
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 2964 5244 3016 5296
rect 2596 5176 2648 5228
rect 5724 5244 5776 5296
rect 8024 5244 8076 5296
rect 3976 5176 4028 5228
rect 4896 5176 4948 5228
rect 7288 5176 7340 5228
rect 4068 5108 4120 5160
rect 8392 5176 8444 5228
rect 8576 5176 8628 5228
rect 16028 5244 16080 5296
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 11888 5176 11940 5228
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 14832 5176 14884 5228
rect 15660 5176 15712 5228
rect 17868 5219 17920 5228
rect 17868 5185 17877 5219
rect 17877 5185 17911 5219
rect 17911 5185 17920 5219
rect 17868 5176 17920 5185
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 19064 5108 19116 5160
rect 7932 5083 7984 5092
rect 7932 5049 7941 5083
rect 7941 5049 7975 5083
rect 7975 5049 7984 5083
rect 7932 5040 7984 5049
rect 16212 5083 16264 5092
rect 16212 5049 16221 5083
rect 16221 5049 16255 5083
rect 16255 5049 16264 5083
rect 16212 5040 16264 5049
rect 16948 5040 17000 5092
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 5172 4972 5224 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 14648 4972 14700 5024
rect 16856 4972 16908 5024
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 2964 4768 3016 4820
rect 7472 4768 7524 4820
rect 9680 4768 9732 4820
rect 11152 4768 11204 4820
rect 4436 4700 4488 4752
rect 9128 4743 9180 4752
rect 9128 4709 9137 4743
rect 9137 4709 9171 4743
rect 9171 4709 9180 4743
rect 9128 4700 9180 4709
rect 15292 4700 15344 4752
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3516 4564 3568 4616
rect 4896 4632 4948 4684
rect 3976 4496 4028 4548
rect 7472 4564 7524 4616
rect 13268 4632 13320 4684
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 8116 4564 8168 4616
rect 8576 4564 8628 4616
rect 9588 4564 9640 4616
rect 17224 4564 17276 4616
rect 12808 4496 12860 4548
rect 12900 4539 12952 4548
rect 12900 4505 12909 4539
rect 12909 4505 12943 4539
rect 12943 4505 12952 4539
rect 12900 4496 12952 4505
rect 16304 4496 16356 4548
rect 17408 4496 17460 4548
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 7380 4428 7432 4480
rect 8024 4428 8076 4480
rect 15200 4428 15252 4480
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 4436 4224 4488 4276
rect 7196 4224 7248 4276
rect 8024 4224 8076 4276
rect 3332 4156 3384 4208
rect 12900 4224 12952 4276
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 1860 4088 1912 4140
rect 4160 4088 4212 4140
rect 4988 4088 5040 4140
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6736 4088 6788 4140
rect 6920 4088 6972 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 9588 4156 9640 4208
rect 3056 4020 3108 4072
rect 8392 4088 8444 4140
rect 8116 4020 8168 4072
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 15016 4156 15068 4208
rect 15844 4199 15896 4208
rect 15844 4165 15853 4199
rect 15853 4165 15887 4199
rect 15887 4165 15896 4199
rect 15844 4156 15896 4165
rect 16948 4156 17000 4208
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 14648 4088 14700 4140
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 7104 3952 7156 4004
rect 16856 3952 16908 4004
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7012 3884 7064 3936
rect 7748 3884 7800 3936
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 8576 3884 8628 3936
rect 15568 3884 15620 3936
rect 17868 3884 17920 3936
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 3056 3723 3108 3732
rect 3056 3689 3065 3723
rect 3065 3689 3099 3723
rect 3099 3689 3108 3723
rect 3056 3680 3108 3689
rect 3976 3680 4028 3732
rect 6920 3680 6972 3732
rect 7380 3680 7432 3732
rect 8392 3680 8444 3732
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 15660 3680 15712 3732
rect 4160 3476 4212 3528
rect 5172 3519 5224 3528
rect 5172 3485 5190 3519
rect 5190 3485 5224 3519
rect 5172 3476 5224 3485
rect 5724 3476 5776 3528
rect 7932 3544 7984 3596
rect 8300 3544 8352 3596
rect 6828 3476 6880 3528
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 17500 3544 17552 3596
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 8668 3408 8720 3460
rect 11152 3408 11204 3460
rect 13360 3476 13412 3528
rect 13912 3476 13964 3528
rect 15200 3519 15252 3528
rect 15200 3485 15234 3519
rect 15234 3485 15252 3519
rect 15200 3476 15252 3485
rect 15568 3408 15620 3460
rect 7288 3340 7340 3392
rect 7472 3340 7524 3392
rect 11704 3340 11756 3392
rect 16304 3383 16356 3392
rect 16304 3349 16313 3383
rect 16313 3349 16347 3383
rect 16347 3349 16356 3383
rect 16304 3340 16356 3349
rect 17316 3340 17368 3392
rect 17868 3340 17920 3392
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 4436 3179 4488 3188
rect 4436 3145 4445 3179
rect 4445 3145 4479 3179
rect 4479 3145 4488 3179
rect 4436 3136 4488 3145
rect 5724 3136 5776 3188
rect 15292 3136 15344 3188
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17224 3179 17276 3188
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 2964 3111 3016 3120
rect 2964 3077 2973 3111
rect 2973 3077 3007 3111
rect 3007 3077 3016 3111
rect 2964 3068 3016 3077
rect 2596 3000 2648 3052
rect 4068 3000 4120 3052
rect 8300 3068 8352 3120
rect 16304 3068 16356 3120
rect 6736 3000 6788 3052
rect 6644 2975 6696 2984
rect 6644 2941 6653 2975
rect 6653 2941 6687 2975
rect 6687 2941 6696 2975
rect 6644 2932 6696 2941
rect 7104 2932 7156 2984
rect 8576 3000 8628 3052
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 15016 3000 15068 3052
rect 7932 2932 7984 2984
rect 9128 2932 9180 2984
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 5540 2796 5592 2848
rect 7380 2839 7432 2848
rect 7380 2805 7389 2839
rect 7389 2805 7423 2839
rect 7423 2805 7432 2839
rect 7380 2796 7432 2805
rect 9220 2796 9272 2848
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 16212 2592 16264 2644
rect 7380 2456 7432 2508
rect 7472 2456 7524 2508
rect 848 2320 900 2372
rect 2504 2320 2556 2372
rect 4160 2320 4212 2372
rect 5540 2388 5592 2440
rect 6828 2388 6880 2440
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 17224 2456 17276 2508
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 13360 2388 13412 2440
rect 15660 2388 15712 2440
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 5816 2320 5868 2372
rect 7472 2320 7524 2372
rect 9128 2320 9180 2372
rect 11060 2320 11112 2372
rect 12440 2320 12492 2372
rect 14096 2320 14148 2372
rect 15752 2320 15804 2372
rect 17316 2320 17368 2372
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 4986 19200 5042 20000
rect 14922 19200 14978 20000
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 5000 15978 5028 19200
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 14936 17270 14964 19200
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 14924 17264 14976 17270
rect 14924 17206 14976 17212
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 9048 16114 9076 16458
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 10428 16250 10456 16594
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10520 16114 10548 17138
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16522 10732 16934
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 11716 16250 11744 16526
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 8496 15570 8524 15846
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 8496 15026 8524 15302
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 10244 15094 10272 15846
rect 10428 15434 10456 15846
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 9416 14074 9444 14894
rect 9876 14414 9904 14894
rect 9864 14408 9916 14414
rect 9692 14356 9864 14362
rect 9692 14350 9916 14356
rect 9692 14334 9904 14350
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9692 13938 9720 14334
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 10244 13394 10272 14214
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 5388 13019 5696 13028
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11762 4568 12038
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 6288 11762 6316 12106
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3332 10736 3384 10742
rect 3528 10724 3556 10950
rect 3384 10696 3556 10724
rect 3332 10678 3384 10684
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3528 10062 3556 10696
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 9178 2636 9454
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2792 8974 2820 9998
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9178 2912 9454
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3068 8974 3096 9318
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 3528 9042 3556 9998
rect 3896 9178 3924 11698
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11286 4384 11494
rect 6288 11286 6316 11698
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6380 11354 6408 11630
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4080 10198 4108 10610
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4172 10062 4200 11154
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2516 8090 2544 8366
rect 2792 8090 2820 8366
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3068 7886 3096 8910
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 3988 7954 4016 9522
rect 4172 8498 4200 9998
rect 4264 8974 4292 10202
rect 4356 10062 4384 11222
rect 6288 11150 6316 11222
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 4356 7886 4384 9998
rect 4448 8838 4476 10406
rect 5276 10266 5304 11018
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 6932 10810 6960 12106
rect 7024 11898 7052 12854
rect 7116 12850 7144 13126
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7392 12306 7420 13262
rect 10336 13258 10364 13670
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11626 7144 12038
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7116 10674 7144 11562
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11286 7236 11494
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5920 9178 5948 9522
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4540 8430 4568 8842
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 6932 8650 6960 8842
rect 7116 8838 7144 10610
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 5172 8628 5224 8634
rect 6932 8622 7144 8650
rect 5172 8570 5224 8576
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 7954 4568 8366
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 6390 3372 6666
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3344 6202 3372 6326
rect 3344 6174 3556 6202
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 3528 5896 3556 6174
rect 3436 5868 3556 5896
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2608 5234 2636 5646
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1872 4146 1900 4422
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2608 3058 2636 4966
rect 2976 4826 3004 5238
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2976 3126 3004 4762
rect 3068 4622 3096 5646
rect 3436 5370 3464 5868
rect 3804 5846 3832 6326
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3988 5778 4016 6598
rect 4356 6254 4384 7822
rect 4540 7546 4568 7890
rect 5000 7886 5028 8434
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 6458 4844 6734
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3528 4622 3556 5646
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4816 5370 4844 5578
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4908 5234 4936 7686
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3988 4554 4016 5170
rect 4068 5160 4120 5166
rect 4120 5108 4200 5114
rect 4068 5102 4200 5108
rect 4080 5086 4200 5102
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4214 3372 4422
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3068 3738 3096 4014
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 3988 3738 4016 4490
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 4080 3058 4108 4422
rect 4172 4146 4200 5086
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4448 4282 4476 4694
rect 4908 4690 4936 5170
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 3534 4200 4082
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4448 3194 4476 4218
rect 5000 4146 5028 7278
rect 5736 6662 5764 8366
rect 7024 7970 7052 8434
rect 7116 8072 7144 8622
rect 7208 8566 7236 11222
rect 7300 11218 7328 12106
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7944 11286 7972 11766
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 8312 10130 8340 12242
rect 8496 11218 8524 12582
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11762 8708 12038
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9140 11286 9168 11834
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7300 8838 7328 9930
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8974 7420 9318
rect 7484 9042 7512 9998
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9586 7696 9930
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7484 8906 7512 8978
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8634 7328 8774
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7196 8560 7248 8566
rect 7484 8514 7512 8842
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7196 8502 7248 8508
rect 7392 8498 7512 8514
rect 7380 8492 7512 8498
rect 7432 8486 7512 8492
rect 7380 8434 7432 8440
rect 7392 8090 7420 8434
rect 7576 8378 7604 8774
rect 7484 8350 7604 8378
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8356 8076 8362
rect 7380 8084 7432 8090
rect 7116 8044 7236 8072
rect 7024 7942 7144 7970
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6656 6798 6684 7210
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6932 6730 6960 7142
rect 7024 6798 7052 7754
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 7116 5914 7144 7942
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 5736 5302 5764 5850
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5184 3534 5212 4966
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 7208 4282 7236 8044
rect 7380 8026 7432 8032
rect 7392 7206 7420 8026
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 6798 7420 7142
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 5736 3194 5764 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 6656 2990 6684 4082
rect 6748 3058 6776 4082
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3534 6868 3878
rect 6932 3738 6960 4082
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 5552 2446 5580 2790
rect 6840 2446 6868 3334
rect 7024 2446 7052 3878
rect 7116 2990 7144 3946
rect 7300 3398 7328 5170
rect 7484 4826 7512 8350
rect 8024 8298 8076 8304
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7852 6254 7880 6734
rect 7944 6458 7972 6734
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 8036 5302 8064 8298
rect 8128 7886 8156 8366
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8312 7546 8340 10066
rect 8404 10062 8432 10746
rect 9140 10606 9168 11222
rect 9600 11150 9628 12174
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 10428 11898 10456 12106
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10742 9260 10950
rect 9600 10810 9628 11086
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8128 6390 8156 7482
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 5710 8248 6190
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4622 7512 4762
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 3738 7420 4422
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7760 3942 7788 4082
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7944 3602 7972 5034
rect 8036 4486 8064 5238
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4282 8064 4422
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7392 2514 7420 2790
rect 7484 2514 7512 3334
rect 7944 2990 7972 3538
rect 8036 3534 8064 4218
rect 8128 4078 8156 4558
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8128 3534 8156 4014
rect 8220 3534 8248 5510
rect 8312 3602 8340 7482
rect 8404 7274 8432 9454
rect 8496 7818 8524 9522
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 5234 8432 6598
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 5914 8524 6190
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8588 5778 8616 9386
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8566 9444 8774
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7410 9352 7686
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9232 5914 9260 6326
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5234 8616 5714
rect 9324 5710 9352 7346
rect 9508 6798 9536 8366
rect 9600 6798 9628 8842
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9692 6730 9720 8910
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 10428 8650 10456 11834
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10062 10548 10610
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10336 8622 10456 8650
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 10244 6322 10272 7822
rect 10336 6798 10364 8622
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10428 7546 10456 8502
rect 10520 7954 10548 9998
rect 10796 8974 10824 15914
rect 11072 15026 11100 16050
rect 11716 15570 11744 16050
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 12820 15570 12848 15846
rect 13740 15570 13768 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12728 15162 12756 15370
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 14108 15026 14136 16594
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 14660 16182 14688 16390
rect 15028 16250 15056 16526
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15120 16182 15148 16390
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 15570 14596 15846
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14200 15162 14228 15438
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11164 13190 11192 13874
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11808 12986 11836 13194
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12850 11928 14962
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 13648 13530 13676 13806
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 11218 11192 12582
rect 11900 12442 11928 12786
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 13832 11830 13860 14826
rect 14200 14414 14228 14962
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13924 14006 13952 14214
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13924 11694 13952 12106
rect 14108 11830 14136 12582
rect 14568 12170 14596 12786
rect 14660 12306 14688 13126
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11164 10470 11192 11018
rect 11900 10810 11928 11018
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11992 10674 12020 10950
rect 12636 10742 12664 11154
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11152 10464 11204 10470
rect 11992 10418 12020 10610
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 11152 10406 11204 10412
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9042 11008 9522
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10704 8566 10732 8910
rect 10980 8634 11008 8978
rect 11164 8906 11192 10406
rect 11900 10390 12020 10418
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9586 11744 9862
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 11072 7886 11100 8774
rect 11808 8634 11836 8910
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 11072 7478 11100 7822
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11808 7410 11836 8570
rect 11900 7886 11928 10390
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 13188 10266 13216 10542
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 13004 9178 13032 9998
rect 13188 9178 13216 10202
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 12728 8022 12756 8502
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 13188 7886 13216 9114
rect 13464 9042 13492 9318
rect 14568 9110 14596 9522
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8430 13308 8910
rect 13464 8634 13492 8978
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11900 6866 11928 7822
rect 13188 7478 13216 7822
rect 13280 7546 13308 8366
rect 14016 7954 14044 8842
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 14016 7478 14044 7890
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14200 7410 14228 7686
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 14200 6866 14228 7142
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5778 11192 6054
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 11072 5370 11100 5578
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11900 5234 11928 6802
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6322 14136 6598
rect 14200 6458 14228 6666
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 12636 5914 12664 6258
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 14108 5710 14136 6258
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 5370 12204 5578
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 8404 4146 8432 5170
rect 8588 4622 8616 5170
rect 11164 4826 11192 5170
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8404 3738 8432 3878
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8312 3126 8340 3538
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8588 3058 8616 3878
rect 9140 3534 9168 4694
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4214 9628 4558
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9692 4146 9720 4762
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8680 3058 8708 3402
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 9140 2990 9168 3470
rect 11164 3466 11192 4762
rect 12820 4554 12848 4966
rect 13280 4690 13308 5510
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 14844 5234 14872 14894
rect 15120 14414 15148 15030
rect 15304 14958 15332 17002
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16114 15516 16390
rect 16132 16114 16160 16526
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15570 16160 16050
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 15162 15700 15438
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 13938 15056 14214
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15120 12918 15148 14350
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 11830 15056 12582
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15396 11694 15424 14962
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 14006 15700 14282
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12238 15700 12582
rect 16316 12306 16344 13262
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 7954 15424 11630
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 18705 8732 19013 8741
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15304 7546 15332 7754
rect 15948 7546 15976 7754
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15488 6322 15516 7346
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6458 15608 6666
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 16316 5710 16344 7890
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12912 4282 12940 4490
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 12728 3738 12756 4082
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 13372 3534 13400 4082
rect 13924 3534 13952 5170
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14016 4146 14044 4966
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 14660 4146 14688 4966
rect 14844 4690 14872 5170
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 9232 2446 9260 2790
rect 11716 2446 11744 3334
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 13372 2446 13400 3470
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 15028 3058 15056 4150
rect 15212 3534 15240 4422
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15304 3194 15332 4694
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3466 15608 3878
rect 15672 3738 15700 5170
rect 15764 4690 15792 5510
rect 16040 5302 16068 5646
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15856 4214 15884 5102
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15580 2972 15608 3402
rect 15660 2984 15712 2990
rect 15580 2944 15660 2972
rect 15660 2926 15712 2932
rect 15672 2446 15700 2926
rect 16224 2650 16252 5034
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16304 4548 16356 4554
rect 16304 4490 16356 4496
rect 16316 4282 16344 4490
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16868 4146 16896 4966
rect 16960 4214 16988 5034
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3126 16344 3334
rect 16868 3194 16896 3946
rect 17236 3194 17264 4558
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16316 2446 16344 3062
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 17236 2514 17264 3130
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 17328 2378 17356 3334
rect 848 2372 900 2378
rect 848 2314 900 2320
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 860 800 888 2314
rect 2516 800 2544 2314
rect 4172 800 4200 2314
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 5828 800 5856 2314
rect 7484 800 7512 2314
rect 9140 800 9168 2314
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 11072 898 11100 2314
rect 10796 870 11100 898
rect 10796 800 10824 870
rect 12452 800 12480 2314
rect 14108 800 14136 2314
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 15764 800 15792 2314
rect 17420 800 17448 4490
rect 17880 3942 17908 5170
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17512 2990 17540 3538
rect 17880 3398 17908 3878
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17512 2514 17540 2926
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 19076 800 19104 5102
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9126 0 9182 800
rect 10782 0 10838 800
rect 12438 0 12494 800
rect 14094 0 14150 800
rect 15750 0 15806 800
rect 17406 0 17462 800
rect 19062 0 19118 800
<< via2 >>
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 5384 16352 5700 16353
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 18701 15199 19017 15200
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 5384 13088 5700 13089
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 5384 9824 5700 9825
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 18701 8671 19017 8672
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 16896 3483 17456
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 17440 5702 17456
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 16896 7922 17456
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 17440 10141 17456
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9821 15264 10141 16288
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9821 12000 10141 13024
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 16896 12361 17456
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 14720 12361 15744
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11456 12361 12480
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 17440 14580 17456
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 14260 15264 14580 16288
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 14260 10912 14580 11936
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 16896 16800 17456
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11456 16800 12480
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 17440 19019 17456
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1676037725
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_157
timestamp 1676037725
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_180
timestamp 1676037725
transform 1 0 17664 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_64
timestamp 1676037725
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_85
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1676037725
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp 1676037725
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1676037725
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1676037725
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_101
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_127
timestamp 1676037725
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1676037725
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_37
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1676037725
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1676037725
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1676037725
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1676037725
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1676037725
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_121
timestamp 1676037725
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1676037725
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1676037725
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_36
timestamp 1676037725
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_48
timestamp 1676037725
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_60
timestamp 1676037725
transform 1 0 6624 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1676037725
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1676037725
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_91
timestamp 1676037725
transform 1 0 9476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_103
timestamp 1676037725
transform 1 0 10580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1676037725
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1676037725
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1676037725
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_29
timestamp 1676037725
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1676037725
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1676037725
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_86
timestamp 1676037725
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_98
timestamp 1676037725
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1676037725
transform 1 0 10856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1676037725
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_129
timestamp 1676037725
transform 1 0 12972 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1676037725
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_151
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_159
timestamp 1676037725
transform 1 0 15732 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_175
timestamp 1676037725
transform 1 0 17204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_52
timestamp 1676037725
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_64
timestamp 1676037725
transform 1 0 6992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1676037725
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_90
timestamp 1676037725
transform 1 0 9384 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1676037725
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1676037725
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1676037725
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_163
timestamp 1676037725
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_175
timestamp 1676037725
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_187
timestamp 1676037725
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_42
timestamp 1676037725
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_72
timestamp 1676037725
transform 1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_97
timestamp 1676037725
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1676037725
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_118
timestamp 1676037725
transform 1 0 11960 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_138
timestamp 1676037725
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1676037725
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1676037725
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1676037725
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1676037725
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1676037725
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_176
timestamp 1676037725
transform 1 0 17296 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1676037725
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1676037725
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_67
timestamp 1676037725
transform 1 0 7268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1676037725
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1676037725
transform 1 0 13248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_140
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_144
timestamp 1676037725
transform 1 0 14352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_152
timestamp 1676037725
transform 1 0 15088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1676037725
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1676037725
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1676037725
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_94
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_100
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1676037725
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1676037725
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_143
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1676037725
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_38
timestamp 1676037725
transform 1 0 4600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1676037725
transform 1 0 5704 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1676037725
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1676037725
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1676037725
transform 1 0 9936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_104
timestamp 1676037725
transform 1 0 10672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1676037725
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_148
timestamp 1676037725
transform 1 0 14720 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_172
timestamp 1676037725
transform 1 0 16928 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_184
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_37
timestamp 1676037725
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_94
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1676037725
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1676037725
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_19
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_48
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_60
timestamp 1676037725
transform 1 0 6624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1676037725
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1676037725
transform 1 0 10396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1676037725
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1676037725
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1676037725
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_91
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1676037725
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1676037725
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1676037725
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1676037725
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1676037725
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_99
timestamp 1676037725
transform 1 0 10212 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1676037725
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_46
timestamp 1676037725
transform 1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1676037725
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_83
timestamp 1676037725
transform 1 0 8740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_156
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1676037725
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_40
timestamp 1676037725
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1676037725
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_90
timestamp 1676037725
transform 1 0 9384 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_166
timestamp 1676037725
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_178
timestamp 1676037725
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_94
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_106
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_118
timestamp 1676037725
transform 1 0 11960 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_130
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_142
timestamp 1676037725
transform 1 0 14168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_69
timestamp 1676037725
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_119
timestamp 1676037725
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_148
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_160
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_92
timestamp 1676037725
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_98
timestamp 1676037725
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1676037725
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1676037725
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_128
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_143
timestamp 1676037725
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1676037725
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_71
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1676037725
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1676037725
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_178
timestamp 1676037725
transform 1 0 17480 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1676037725
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1676037725
transform 1 0 8648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1676037725
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1676037725
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1676037725
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1676037725
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_157
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1676037725
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_116
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_128
timestamp 1676037725
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_161
timestamp 1676037725
transform 1 0 15916 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1676037725
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1676037725
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1676037725
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1676037725
transform -1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1676037725
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1676037725
transform -1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1676037725
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1676037725
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1676037725
transform -1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1676037725
transform -1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1676037725
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1676037725
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1676037725
transform -1 0 14720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1676037725
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1676037725
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1676037725
transform -1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1676037725
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1676037725
transform -1 0 8004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1676037725
transform -1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1676037725
transform 1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1676037725
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125__1
timestamp 1676037725
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15180 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _127__10
timestamp 1676037725
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _129_
timestamp 1676037725
transform -1 0 4416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _130_
timestamp 1676037725
transform -1 0 10764 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _131_
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _132_
timestamp 1676037725
transform 1 0 12512 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _136_
timestamp 1676037725
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 1676037725
transform 1 0 15180 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _138_
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14996 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4600 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _142_
timestamp 1676037725
transform 1 0 3128 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _144_
timestamp 1676037725
transform -1 0 13616 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  _146_
timestamp 1676037725
transform 1 0 6440 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1676037725
transform -1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9752 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9752 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_4  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1676037725
transform -1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _156_
timestamp 1676037725
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1676037725
transform -1 0 5520 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _159_
timestamp 1676037725
transform -1 0 8372 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8004 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1676037725
transform -1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _168_
timestamp 1676037725
transform 1 0 8372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _171_
timestamp 1676037725
transform -1 0 8924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _172_
timestamp 1676037725
transform -1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _173__11
timestamp 1676037725
transform -1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__12
timestamp 1676037725
transform -1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175__13
timestamp 1676037725
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _176_
timestamp 1676037725
transform -1 0 4416 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _177_
timestamp 1676037725
transform 1 0 3036 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _178_
timestamp 1676037725
transform -1 0 4416 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _179_
timestamp 1676037725
transform 1 0 4968 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _180_
timestamp 1676037725
transform -1 0 13064 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _181_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _182_
timestamp 1676037725
transform 1 0 11776 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _183_
timestamp 1676037725
transform 1 0 7728 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _184__14
timestamp 1676037725
transform -1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185__15
timestamp 1676037725
transform -1 0 12880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186__16
timestamp 1676037725
transform -1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187__17
timestamp 1676037725
transform 1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188__18
timestamp 1676037725
transform -1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189__19
timestamp 1676037725
transform -1 0 14628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190__20
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191__21
timestamp 1676037725
transform -1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192__22
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193__2
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194__3
timestamp 1676037725
transform -1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195__4
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196__5
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197__23
timestamp 1676037725
transform -1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1676037725
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1676037725
transform -1 0 14260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1676037725
transform -1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform -1 0 11224 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1676037725
transform -1 0 8648 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1676037725
transform -1 0 13064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207__6
timestamp 1676037725
transform -1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208__7
timestamp 1676037725
transform -1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _209_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1676037725
transform -1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1676037725
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1676037725
transform -1 0 11224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1676037725
transform 1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1676037725
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1676037725
transform -1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216__8
timestamp 1676037725
transform -1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217__9
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1676037725
transform -1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1676037725
transform -1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1676037725
transform -1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _221_
timestamp 1676037725
transform 1 0 3036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1676037725
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1676037725
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _225_
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1676037725
transform -1 0 10672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1676037725
transform -1 0 11224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1676037725
transform -1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1676037725
transform -1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230__24
timestamp 1676037725
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13984 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1676037725
transform 1 0 14904 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1676037725
transform 1 0 15732 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1676037725
transform 1 0 11316 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _237_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _238_
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _239_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _240_
timestamp 1676037725
transform -1 0 15548 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _241_
timestamp 1676037725
transform 1 0 9936 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _242_
timestamp 1676037725
transform -1 0 11776 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _243_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _244_
timestamp 1676037725
transform -1 0 13800 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _245_
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_2  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4600 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _247_
timestamp 1676037725
transform -1 0 5520 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9476 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _249_
timestamp 1676037725
transform -1 0 8740 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _250_
timestamp 1676037725
transform 1 0 6532 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _251_
timestamp 1676037725
transform 1 0 10856 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _252_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _253_
timestamp 1676037725
transform -1 0 13616 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _254_
timestamp 1676037725
transform 1 0 9108 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_2  _255_
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfrtp_4  _257_
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _258_
timestamp 1676037725
transform 1 0 2576 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _259_
timestamp 1676037725
transform 1 0 2760 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _260_
timestamp 1676037725
transform -1 0 5888 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _261_
timestamp 1676037725
transform 1 0 2392 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _262_
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _263_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _264_
timestamp 1676037725
transform 1 0 3036 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _265_
timestamp 1676037725
transform -1 0 10028 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _266_
timestamp 1676037725
transform 1 0 10856 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _267_
timestamp 1676037725
transform -1 0 13248 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _268_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _269_
timestamp 1676037725
transform -1 0 16376 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1676037725
transform 1 0 10764 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f__068_
timestamp 1676037725
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f__068_
timestamp 1676037725
transform -1 0 7084 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f__068_
timestamp 1676037725
transform 1 0 10396 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f__068_
timestamp 1676037725
transform 1 0 10396 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output3
timestamp 1676037725
transform 1 0 17572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1676037725
transform 1 0 17848 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform -1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform -1 0 4784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 9200 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 13156 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform -1 0 16376 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 4986 19200 5042 20000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 io_out[0]
port 1 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 io_out[10]
port 2 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 io_out[11]
port 3 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 io_out[1]
port 4 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 io_out[2]
port 5 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 io_out[3]
port 6 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 io_out[4]
port 7 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 io_out[5]
port 8 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 io_out[6]
port 9 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 io_out[7]
port 10 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[8]
port 11 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 io_out[9]
port 12 nsew signal tristate
flabel metal2 s 14922 19200 14978 20000 0 FreeSans 224 90 0 0 rst
port 13 nsew signal input
flabel metal4 s 3163 2128 3483 17456 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 7602 2128 7922 17456 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 12041 2128 12361 17456 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 16480 2128 16800 17456 0 FreeSans 1920 90 0 0 vccd1
port 14 nsew power bidirectional
flabel metal4 s 5382 2128 5702 17456 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 17456 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 17456 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 17456 0 FreeSans 1920 90 0 0 vssd1
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
