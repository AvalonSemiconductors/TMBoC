VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as1802
  CLASS BLOCK ;
  FOREIGN wrapped_as1802 ;
  ORIGIN 0.000 0.000 ;
  SIZE 325.000 BY 325.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.060 4.000 289.260 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.020 4.000 15.220 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.820 4.000 226.020 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.900 4.000 247.100 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.980 4.000 268.180 ;
    END
  END io_in[12]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.180 4.000 57.380 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.260 4.000 78.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.340 4.000 99.540 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.420 4.000 120.620 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.500 4.000 141.700 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.580 4.000 162.780 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.660 4.000 183.860 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.350 0.000 317.910 4.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 0.000 7.410 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.850 0.000 122.410 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 0.000 133.910 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 0.000 145.410 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 0.000 156.910 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 0.000 168.410 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.350 0.000 179.910 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.850 0.000 191.410 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 0.000 202.910 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.850 0.000 214.410 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 0.000 225.910 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.850 0.000 237.410 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.350 0.000 248.910 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.850 0.000 260.410 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 0.000 271.910 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.850 0.000 283.410 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 0.000 294.910 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 0.000 306.410 4.000 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.850 0.000 30.410 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 0.000 41.910 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.850 0.000 53.410 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.850 0.000 76.410 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 0.000 87.910 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 0.000 99.410 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.350 0.000 110.910 4.000 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.140 4.000 310.340 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 313.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 313.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 313.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 313.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 319.240 312.885 ;
      LAYER met1 ;
        RECT 5.520 8.540 319.240 313.040 ;
      LAYER met2 ;
        RECT 6.990 4.280 317.760 312.985 ;
        RECT 7.690 4.000 18.070 4.280 ;
        RECT 19.190 4.000 29.570 4.280 ;
        RECT 30.690 4.000 41.070 4.280 ;
        RECT 42.190 4.000 52.570 4.280 ;
        RECT 53.690 4.000 64.070 4.280 ;
        RECT 65.190 4.000 75.570 4.280 ;
        RECT 76.690 4.000 87.070 4.280 ;
        RECT 88.190 4.000 98.570 4.280 ;
        RECT 99.690 4.000 110.070 4.280 ;
        RECT 111.190 4.000 121.570 4.280 ;
        RECT 122.690 4.000 133.070 4.280 ;
        RECT 134.190 4.000 144.570 4.280 ;
        RECT 145.690 4.000 156.070 4.280 ;
        RECT 157.190 4.000 167.570 4.280 ;
        RECT 168.690 4.000 179.070 4.280 ;
        RECT 180.190 4.000 190.570 4.280 ;
        RECT 191.690 4.000 202.070 4.280 ;
        RECT 203.190 4.000 213.570 4.280 ;
        RECT 214.690 4.000 225.070 4.280 ;
        RECT 226.190 4.000 236.570 4.280 ;
        RECT 237.690 4.000 248.070 4.280 ;
        RECT 249.190 4.000 259.570 4.280 ;
        RECT 260.690 4.000 271.070 4.280 ;
        RECT 272.190 4.000 282.570 4.280 ;
        RECT 283.690 4.000 294.070 4.280 ;
        RECT 295.190 4.000 305.570 4.280 ;
        RECT 306.690 4.000 317.070 4.280 ;
      LAYER met3 ;
        RECT 3.070 310.740 303.995 312.965 ;
        RECT 4.400 308.740 303.995 310.740 ;
        RECT 3.070 289.660 303.995 308.740 ;
        RECT 4.400 287.660 303.995 289.660 ;
        RECT 3.070 268.580 303.995 287.660 ;
        RECT 4.400 266.580 303.995 268.580 ;
        RECT 3.070 247.500 303.995 266.580 ;
        RECT 4.400 245.500 303.995 247.500 ;
        RECT 3.070 226.420 303.995 245.500 ;
        RECT 4.400 224.420 303.995 226.420 ;
        RECT 3.070 205.340 303.995 224.420 ;
        RECT 4.400 203.340 303.995 205.340 ;
        RECT 3.070 184.260 303.995 203.340 ;
        RECT 4.400 182.260 303.995 184.260 ;
        RECT 3.070 163.180 303.995 182.260 ;
        RECT 4.400 161.180 303.995 163.180 ;
        RECT 3.070 142.100 303.995 161.180 ;
        RECT 4.400 140.100 303.995 142.100 ;
        RECT 3.070 121.020 303.995 140.100 ;
        RECT 4.400 119.020 303.995 121.020 ;
        RECT 3.070 99.940 303.995 119.020 ;
        RECT 4.400 97.940 303.995 99.940 ;
        RECT 3.070 78.860 303.995 97.940 ;
        RECT 4.400 76.860 303.995 78.860 ;
        RECT 3.070 57.780 303.995 76.860 ;
        RECT 4.400 55.780 303.995 57.780 ;
        RECT 3.070 36.700 303.995 55.780 ;
        RECT 4.400 34.700 303.995 36.700 ;
        RECT 3.070 15.620 303.995 34.700 ;
        RECT 4.400 13.620 303.995 15.620 ;
        RECT 3.070 9.695 303.995 13.620 ;
      LAYER met4 ;
        RECT 9.495 10.240 20.640 288.825 ;
        RECT 23.040 10.240 97.440 288.825 ;
        RECT 99.840 10.240 174.240 288.825 ;
        RECT 176.640 10.240 251.040 288.825 ;
        RECT 253.440 10.240 291.345 288.825 ;
        RECT 9.495 9.695 291.345 10.240 ;
  END
END wrapped_as1802
END LIBRARY

